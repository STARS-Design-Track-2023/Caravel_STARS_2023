// This is the unpowered netlist.
module silly_synthesizer (clk,
    cs,
    nrst,
    pwm,
    gpio);
 input clk;
 input cs;
 input nrst;
 output pwm;
 input [16:0] gpio;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \inputs.down.det_edge ;
 wire \inputs.down.ff_in ;
 wire \inputs.down.ff_out ;
 wire \inputs.down.in ;
 wire \inputs.frequency_lut.rng[0] ;
 wire \inputs.frequency_lut.rng[1] ;
 wire \inputs.frequency_lut.rng[2] ;
 wire \inputs.frequency_lut.rng[3] ;
 wire \inputs.frequency_lut.rng[4] ;
 wire \inputs.frequency_lut.rng[5] ;
 wire \inputs.key_encoder.mode_key ;
 wire \inputs.key_encoder.octave_key_up ;
 wire \inputs.key_encoder.sync_keys[0] ;
 wire \inputs.key_encoder.sync_keys[10] ;
 wire \inputs.key_encoder.sync_keys[11] ;
 wire \inputs.key_encoder.sync_keys[12] ;
 wire \inputs.key_encoder.sync_keys[13] ;
 wire \inputs.key_encoder.sync_keys[14] ;
 wire \inputs.key_encoder.sync_keys[15] ;
 wire \inputs.key_encoder.sync_keys[1] ;
 wire \inputs.key_encoder.sync_keys[2] ;
 wire \inputs.key_encoder.sync_keys[3] ;
 wire \inputs.key_encoder.sync_keys[4] ;
 wire \inputs.key_encoder.sync_keys[5] ;
 wire \inputs.key_encoder.sync_keys[6] ;
 wire \inputs.key_encoder.sync_keys[7] ;
 wire \inputs.key_encoder.sync_keys[8] ;
 wire \inputs.key_encoder.sync_keys[9] ;
 wire \inputs.keypad[0] ;
 wire \inputs.keypad[10] ;
 wire \inputs.keypad[11] ;
 wire \inputs.keypad[12] ;
 wire \inputs.keypad[13] ;
 wire \inputs.keypad[14] ;
 wire \inputs.keypad[15] ;
 wire \inputs.keypad[16] ;
 wire \inputs.keypad[1] ;
 wire \inputs.keypad[2] ;
 wire \inputs.keypad[3] ;
 wire \inputs.keypad[4] ;
 wire \inputs.keypad[5] ;
 wire \inputs.keypad[6] ;
 wire \inputs.keypad[7] ;
 wire \inputs.keypad[8] ;
 wire \inputs.keypad[9] ;
 wire \inputs.keypad_synchronizer.half_sync[0] ;
 wire \inputs.keypad_synchronizer.half_sync[10] ;
 wire \inputs.keypad_synchronizer.half_sync[11] ;
 wire \inputs.keypad_synchronizer.half_sync[12] ;
 wire \inputs.keypad_synchronizer.half_sync[13] ;
 wire \inputs.keypad_synchronizer.half_sync[14] ;
 wire \inputs.keypad_synchronizer.half_sync[15] ;
 wire \inputs.keypad_synchronizer.half_sync[16] ;
 wire \inputs.keypad_synchronizer.half_sync[1] ;
 wire \inputs.keypad_synchronizer.half_sync[2] ;
 wire \inputs.keypad_synchronizer.half_sync[3] ;
 wire \inputs.keypad_synchronizer.half_sync[4] ;
 wire \inputs.keypad_synchronizer.half_sync[5] ;
 wire \inputs.keypad_synchronizer.half_sync[6] ;
 wire \inputs.keypad_synchronizer.half_sync[7] ;
 wire \inputs.keypad_synchronizer.half_sync[8] ;
 wire \inputs.keypad_synchronizer.half_sync[9] ;
 wire \inputs.mode_edge.det_edge ;
 wire \inputs.mode_edge.ff_in ;
 wire \inputs.mode_edge.ff_out ;
 wire \inputs.octave_fsm.octave_key_up ;
 wire \inputs.octave_fsm.state[0] ;
 wire \inputs.octave_fsm.state[1] ;
 wire \inputs.octave_fsm.state[2] ;
 wire \inputs.random_note_generator.feedback ;
 wire \inputs.random_note_generator.out[0] ;
 wire \inputs.random_note_generator.out[10] ;
 wire \inputs.random_note_generator.out[11] ;
 wire \inputs.random_note_generator.out[12] ;
 wire \inputs.random_note_generator.out[13] ;
 wire \inputs.random_note_generator.out[14] ;
 wire \inputs.random_note_generator.out[15] ;
 wire \inputs.random_note_generator.out[1] ;
 wire \inputs.random_note_generator.out[2] ;
 wire \inputs.random_note_generator.out[3] ;
 wire \inputs.random_note_generator.out[4] ;
 wire \inputs.random_note_generator.out[5] ;
 wire \inputs.random_note_generator.out[6] ;
 wire \inputs.random_note_generator.out[7] ;
 wire \inputs.random_note_generator.out[8] ;
 wire \inputs.random_note_generator.out[9] ;
 wire \inputs.random_update_clock.count[0] ;
 wire \inputs.random_update_clock.count[10] ;
 wire \inputs.random_update_clock.count[11] ;
 wire \inputs.random_update_clock.count[12] ;
 wire \inputs.random_update_clock.count[13] ;
 wire \inputs.random_update_clock.count[14] ;
 wire \inputs.random_update_clock.count[15] ;
 wire \inputs.random_update_clock.count[16] ;
 wire \inputs.random_update_clock.count[17] ;
 wire \inputs.random_update_clock.count[18] ;
 wire \inputs.random_update_clock.count[19] ;
 wire \inputs.random_update_clock.count[1] ;
 wire \inputs.random_update_clock.count[20] ;
 wire \inputs.random_update_clock.count[21] ;
 wire \inputs.random_update_clock.count[22] ;
 wire \inputs.random_update_clock.count[2] ;
 wire \inputs.random_update_clock.count[3] ;
 wire \inputs.random_update_clock.count[4] ;
 wire \inputs.random_update_clock.count[5] ;
 wire \inputs.random_update_clock.count[6] ;
 wire \inputs.random_update_clock.count[7] ;
 wire \inputs.random_update_clock.count[8] ;
 wire \inputs.random_update_clock.count[9] ;
 wire \inputs.random_update_clock.next_count[0] ;
 wire \inputs.random_update_clock.next_count[10] ;
 wire \inputs.random_update_clock.next_count[11] ;
 wire \inputs.random_update_clock.next_count[12] ;
 wire \inputs.random_update_clock.next_count[13] ;
 wire \inputs.random_update_clock.next_count[14] ;
 wire \inputs.random_update_clock.next_count[15] ;
 wire \inputs.random_update_clock.next_count[16] ;
 wire \inputs.random_update_clock.next_count[17] ;
 wire \inputs.random_update_clock.next_count[18] ;
 wire \inputs.random_update_clock.next_count[19] ;
 wire \inputs.random_update_clock.next_count[1] ;
 wire \inputs.random_update_clock.next_count[20] ;
 wire \inputs.random_update_clock.next_count[21] ;
 wire \inputs.random_update_clock.next_count[22] ;
 wire \inputs.random_update_clock.next_count[2] ;
 wire \inputs.random_update_clock.next_count[3] ;
 wire \inputs.random_update_clock.next_count[4] ;
 wire \inputs.random_update_clock.next_count[5] ;
 wire \inputs.random_update_clock.next_count[6] ;
 wire \inputs.random_update_clock.next_count[7] ;
 wire \inputs.random_update_clock.next_count[8] ;
 wire \inputs.random_update_clock.next_count[9] ;
 wire \inputs.up.ff_in ;
 wire \inputs.up.ff_out ;
 wire \inputs.wavetype_fsm.next_state[0] ;
 wire \inputs.wavetype_fsm.next_state[1] ;
 wire \inputs.wavetype_fsm.state[0] ;
 wire \inputs.wavetype_fsm.state[1] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \outputs.div.a[0] ;
 wire \outputs.div.a[10] ;
 wire \outputs.div.a[11] ;
 wire \outputs.div.a[12] ;
 wire \outputs.div.a[13] ;
 wire \outputs.div.a[14] ;
 wire \outputs.div.a[15] ;
 wire \outputs.div.a[16] ;
 wire \outputs.div.a[17] ;
 wire \outputs.div.a[18] ;
 wire \outputs.div.a[19] ;
 wire \outputs.div.a[1] ;
 wire \outputs.div.a[20] ;
 wire \outputs.div.a[21] ;
 wire \outputs.div.a[22] ;
 wire \outputs.div.a[23] ;
 wire \outputs.div.a[24] ;
 wire \outputs.div.a[25] ;
 wire \outputs.div.a[2] ;
 wire \outputs.div.a[3] ;
 wire \outputs.div.a[4] ;
 wire \outputs.div.a[5] ;
 wire \outputs.div.a[6] ;
 wire \outputs.div.a[7] ;
 wire \outputs.div.a[8] ;
 wire \outputs.div.a[9] ;
 wire \outputs.div.count[0] ;
 wire \outputs.div.count[1] ;
 wire \outputs.div.count[2] ;
 wire \outputs.div.count[3] ;
 wire \outputs.div.count[4] ;
 wire \outputs.div.div ;
 wire \outputs.div.divisor[0] ;
 wire \outputs.div.divisor[10] ;
 wire \outputs.div.divisor[11] ;
 wire \outputs.div.divisor[12] ;
 wire \outputs.div.divisor[13] ;
 wire \outputs.div.divisor[14] ;
 wire \outputs.div.divisor[15] ;
 wire \outputs.div.divisor[16] ;
 wire \outputs.div.divisor[17] ;
 wire \outputs.div.divisor[1] ;
 wire \outputs.div.divisor[2] ;
 wire \outputs.div.divisor[3] ;
 wire \outputs.div.divisor[4] ;
 wire \outputs.div.divisor[5] ;
 wire \outputs.div.divisor[6] ;
 wire \outputs.div.divisor[7] ;
 wire \outputs.div.divisor[8] ;
 wire \outputs.div.divisor[9] ;
 wire \outputs.div.m[0] ;
 wire \outputs.div.m[10] ;
 wire \outputs.div.m[11] ;
 wire \outputs.div.m[12] ;
 wire \outputs.div.m[13] ;
 wire \outputs.div.m[14] ;
 wire \outputs.div.m[15] ;
 wire \outputs.div.m[16] ;
 wire \outputs.div.m[17] ;
 wire \outputs.div.m[1] ;
 wire \outputs.div.m[2] ;
 wire \outputs.div.m[3] ;
 wire \outputs.div.m[4] ;
 wire \outputs.div.m[5] ;
 wire \outputs.div.m[6] ;
 wire \outputs.div.m[7] ;
 wire \outputs.div.m[8] ;
 wire \outputs.div.m[9] ;
 wire \outputs.div.next_div ;
 wire \outputs.div.next_start ;
 wire \outputs.div.oscillator_out[0] ;
 wire \outputs.div.oscillator_out[10] ;
 wire \outputs.div.oscillator_out[11] ;
 wire \outputs.div.oscillator_out[12] ;
 wire \outputs.div.oscillator_out[13] ;
 wire \outputs.div.oscillator_out[14] ;
 wire \outputs.div.oscillator_out[15] ;
 wire \outputs.div.oscillator_out[16] ;
 wire \outputs.div.oscillator_out[17] ;
 wire \outputs.div.oscillator_out[1] ;
 wire \outputs.div.oscillator_out[2] ;
 wire \outputs.div.oscillator_out[3] ;
 wire \outputs.div.oscillator_out[4] ;
 wire \outputs.div.oscillator_out[5] ;
 wire \outputs.div.oscillator_out[6] ;
 wire \outputs.div.oscillator_out[7] ;
 wire \outputs.div.oscillator_out[8] ;
 wire \outputs.div.oscillator_out[9] ;
 wire \outputs.div.q[0] ;
 wire \outputs.div.q[10] ;
 wire \outputs.div.q[11] ;
 wire \outputs.div.q[12] ;
 wire \outputs.div.q[13] ;
 wire \outputs.div.q[14] ;
 wire \outputs.div.q[15] ;
 wire \outputs.div.q[16] ;
 wire \outputs.div.q[17] ;
 wire \outputs.div.q[18] ;
 wire \outputs.div.q[19] ;
 wire \outputs.div.q[1] ;
 wire \outputs.div.q[20] ;
 wire \outputs.div.q[21] ;
 wire \outputs.div.q[22] ;
 wire \outputs.div.q[23] ;
 wire \outputs.div.q[24] ;
 wire \outputs.div.q[25] ;
 wire \outputs.div.q[26] ;
 wire \outputs.div.q[2] ;
 wire \outputs.div.q[3] ;
 wire \outputs.div.q[4] ;
 wire \outputs.div.q[5] ;
 wire \outputs.div.q[6] ;
 wire \outputs.div.q[7] ;
 wire \outputs.div.q[8] ;
 wire \outputs.div.q[9] ;
 wire \outputs.div.q_out[0] ;
 wire \outputs.div.q_out[1] ;
 wire \outputs.div.q_out[2] ;
 wire \outputs.div.q_out[3] ;
 wire \outputs.div.q_out[4] ;
 wire \outputs.div.q_out[5] ;
 wire \outputs.div.q_out[6] ;
 wire \outputs.div.q_out[7] ;
 wire \outputs.div.start ;
 wire \outputs.divider_buffer2[0] ;
 wire \outputs.divider_buffer2[10] ;
 wire \outputs.divider_buffer2[11] ;
 wire \outputs.divider_buffer2[12] ;
 wire \outputs.divider_buffer2[13] ;
 wire \outputs.divider_buffer2[14] ;
 wire \outputs.divider_buffer2[15] ;
 wire \outputs.divider_buffer2[16] ;
 wire \outputs.divider_buffer2[17] ;
 wire \outputs.divider_buffer2[1] ;
 wire \outputs.divider_buffer2[2] ;
 wire \outputs.divider_buffer2[3] ;
 wire \outputs.divider_buffer2[4] ;
 wire \outputs.divider_buffer2[5] ;
 wire \outputs.divider_buffer2[6] ;
 wire \outputs.divider_buffer2[7] ;
 wire \outputs.divider_buffer2[8] ;
 wire \outputs.divider_buffer2[9] ;
 wire \outputs.divider_buffer[0] ;
 wire \outputs.divider_buffer[10] ;
 wire \outputs.divider_buffer[11] ;
 wire \outputs.divider_buffer[12] ;
 wire \outputs.divider_buffer[13] ;
 wire \outputs.divider_buffer[14] ;
 wire \outputs.divider_buffer[15] ;
 wire \outputs.divider_buffer[16] ;
 wire \outputs.divider_buffer[17] ;
 wire \outputs.divider_buffer[1] ;
 wire \outputs.divider_buffer[2] ;
 wire \outputs.divider_buffer[3] ;
 wire \outputs.divider_buffer[4] ;
 wire \outputs.divider_buffer[5] ;
 wire \outputs.divider_buffer[6] ;
 wire \outputs.divider_buffer[7] ;
 wire \outputs.divider_buffer[8] ;
 wire \outputs.divider_buffer[9] ;
 wire \outputs.output_gen.count[0] ;
 wire \outputs.output_gen.count[1] ;
 wire \outputs.output_gen.count[2] ;
 wire \outputs.output_gen.count[3] ;
 wire \outputs.output_gen.count[4] ;
 wire \outputs.output_gen.count[5] ;
 wire \outputs.output_gen.count[6] ;
 wire \outputs.output_gen.count[7] ;
 wire \outputs.output_gen.next_count[0] ;
 wire \outputs.output_gen.next_count[1] ;
 wire \outputs.output_gen.next_count[2] ;
 wire \outputs.output_gen.next_count[3] ;
 wire \outputs.output_gen.next_count[4] ;
 wire \outputs.output_gen.next_count[5] ;
 wire \outputs.output_gen.next_count[6] ;
 wire \outputs.output_gen.next_count[7] ;
 wire \outputs.output_gen.pwm_ff ;
 wire \outputs.output_gen.pwm_unff ;
 wire \outputs.pwm_output ;
 wire \outputs.sample_rate.count[0] ;
 wire \outputs.sample_rate.count[1] ;
 wire \outputs.sample_rate.count[2] ;
 wire \outputs.sample_rate.count[3] ;
 wire \outputs.sample_rate.count[4] ;
 wire \outputs.sample_rate.count[5] ;
 wire \outputs.sample_rate.count[6] ;
 wire \outputs.sample_rate.count[7] ;
 wire \outputs.sample_rate.next_count[0] ;
 wire \outputs.sample_rate.next_count[1] ;
 wire \outputs.sample_rate.next_count[2] ;
 wire \outputs.sample_rate.next_count[3] ;
 wire \outputs.sample_rate.next_count[4] ;
 wire \outputs.sample_rate.next_count[5] ;
 wire \outputs.sample_rate.next_count[6] ;
 wire \outputs.sample_rate.next_count[7] ;
 wire \outputs.scaled_buffer[0] ;
 wire \outputs.scaled_buffer[1] ;
 wire \outputs.scaled_buffer[2] ;
 wire \outputs.scaled_buffer[3] ;
 wire \outputs.scaled_buffer[4] ;
 wire \outputs.scaled_buffer[5] ;
 wire \outputs.scaled_buffer[6] ;
 wire \outputs.scaled_buffer[7] ;
 wire \outputs.shaper.count[0] ;
 wire \outputs.shaper.count[10] ;
 wire \outputs.shaper.count[11] ;
 wire \outputs.shaper.count[12] ;
 wire \outputs.shaper.count[13] ;
 wire \outputs.shaper.count[14] ;
 wire \outputs.shaper.count[15] ;
 wire \outputs.shaper.count[16] ;
 wire \outputs.shaper.count[17] ;
 wire \outputs.shaper.count[1] ;
 wire \outputs.shaper.count[2] ;
 wire \outputs.shaper.count[3] ;
 wire \outputs.shaper.count[4] ;
 wire \outputs.shaper.count[5] ;
 wire \outputs.shaper.count[6] ;
 wire \outputs.shaper.count[7] ;
 wire \outputs.shaper.count[8] ;
 wire \outputs.shaper.count[9] ;
 wire \outputs.sig_gen.count[0] ;
 wire \outputs.sig_gen.count[10] ;
 wire \outputs.sig_gen.count[11] ;
 wire \outputs.sig_gen.count[12] ;
 wire \outputs.sig_gen.count[13] ;
 wire \outputs.sig_gen.count[14] ;
 wire \outputs.sig_gen.count[15] ;
 wire \outputs.sig_gen.count[16] ;
 wire \outputs.sig_gen.count[17] ;
 wire \outputs.sig_gen.count[1] ;
 wire \outputs.sig_gen.count[2] ;
 wire \outputs.sig_gen.count[3] ;
 wire \outputs.sig_gen.count[4] ;
 wire \outputs.sig_gen.count[5] ;
 wire \outputs.sig_gen.count[6] ;
 wire \outputs.sig_gen.count[7] ;
 wire \outputs.sig_gen.count[8] ;
 wire \outputs.sig_gen.count[9] ;
 wire \outputs.sig_gen.next_count[0] ;
 wire \outputs.sig_gen.next_count[10] ;
 wire \outputs.sig_gen.next_count[11] ;
 wire \outputs.sig_gen.next_count[12] ;
 wire \outputs.sig_gen.next_count[13] ;
 wire \outputs.sig_gen.next_count[14] ;
 wire \outputs.sig_gen.next_count[15] ;
 wire \outputs.sig_gen.next_count[16] ;
 wire \outputs.sig_gen.next_count[17] ;
 wire \outputs.sig_gen.next_count[1] ;
 wire \outputs.sig_gen.next_count[2] ;
 wire \outputs.sig_gen.next_count[3] ;
 wire \outputs.sig_gen.next_count[4] ;
 wire \outputs.sig_gen.next_count[5] ;
 wire \outputs.sig_gen.next_count[6] ;
 wire \outputs.sig_gen.next_count[7] ;
 wire \outputs.sig_gen.next_count[8] ;
 wire \outputs.sig_gen.next_count[9] ;
 wire \outputs.signal_buffer2[0] ;
 wire \outputs.signal_buffer2[10] ;
 wire \outputs.signal_buffer2[11] ;
 wire \outputs.signal_buffer2[12] ;
 wire \outputs.signal_buffer2[13] ;
 wire \outputs.signal_buffer2[14] ;
 wire \outputs.signal_buffer2[15] ;
 wire \outputs.signal_buffer2[16] ;
 wire \outputs.signal_buffer2[17] ;
 wire \outputs.signal_buffer2[1] ;
 wire \outputs.signal_buffer2[2] ;
 wire \outputs.signal_buffer2[3] ;
 wire \outputs.signal_buffer2[4] ;
 wire \outputs.signal_buffer2[5] ;
 wire \outputs.signal_buffer2[6] ;
 wire \outputs.signal_buffer2[7] ;
 wire \outputs.signal_buffer2[8] ;
 wire \outputs.signal_buffer2[9] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__and3_1 _1295_ (.A(\outputs.sample_rate.count[2] ),
    .B(\outputs.sample_rate.count[1] ),
    .C(\outputs.sample_rate.count[0] ),
    .X(_0994_));
 sky130_fd_sc_hd__and2_1 _1296_ (.A(\outputs.sample_rate.count[3] ),
    .B(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__and3_1 _1297_ (.A(\outputs.sample_rate.count[4] ),
    .B(\outputs.sample_rate.count[5] ),
    .C(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__and2_1 _1298_ (.A(\outputs.sample_rate.count[6] ),
    .B(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__nand2_1 _1299_ (.A(\outputs.sample_rate.count[7] ),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__a21o_1 _1300_ (.A1(\outputs.div.count[1] ),
    .A2(\outputs.div.count[0] ),
    .B1(\outputs.div.count[2] ),
    .X(_0999_));
 sky130_fd_sc_hd__inv_2 _1301_ (.A(\outputs.div.start ),
    .Y(_1000_));
 sky130_fd_sc_hd__a31o_1 _1302_ (.A1(\outputs.div.count[3] ),
    .A2(\outputs.div.count[4] ),
    .A3(_0999_),
    .B1(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__and2_1 _1303_ (.A(_0998_),
    .B(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__clkbuf_4 _1304_ (.A(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_4 _1305_ (.A(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__inv_2 _1306_ (.A(_1004_),
    .Y(\outputs.div.next_start ));
 sky130_fd_sc_hd__clkbuf_4 _1307_ (.A(net1),
    .X(_1005_));
 sky130_fd_sc_hd__and2b_1 _1308_ (.A_N(_1005_),
    .B(net2),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_1 _1309_ (.A(_1006_),
    .X(\inputs.keypad[0] ));
 sky130_fd_sc_hd__and2b_1 _1310_ (.A_N(_1005_),
    .B(net10),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_1 _1311_ (.A(_1007_),
    .X(\inputs.keypad[1] ));
 sky130_fd_sc_hd__and2b_1 _1312_ (.A_N(_1005_),
    .B(net11),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_1 _1313_ (.A(_1008_),
    .X(\inputs.keypad[2] ));
 sky130_fd_sc_hd__and2b_1 _1314_ (.A_N(_1005_),
    .B(net12),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _1315_ (.A(_1009_),
    .X(\inputs.keypad[3] ));
 sky130_fd_sc_hd__and2b_1 _1316_ (.A_N(_1005_),
    .B(net13),
    .X(_1010_));
 sky130_fd_sc_hd__buf_1 _1317_ (.A(_1010_),
    .X(\inputs.keypad[4] ));
 sky130_fd_sc_hd__and2b_1 _1318_ (.A_N(_1005_),
    .B(net14),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_1 _1319_ (.A(_1011_),
    .X(\inputs.keypad[5] ));
 sky130_fd_sc_hd__and2b_1 _1320_ (.A_N(_1005_),
    .B(net15),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _1321_ (.A(_1012_),
    .X(\inputs.keypad[6] ));
 sky130_fd_sc_hd__and2b_1 _1322_ (.A_N(_1005_),
    .B(net16),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _1323_ (.A(_1013_),
    .X(\inputs.keypad[7] ));
 sky130_fd_sc_hd__and2b_1 _1324_ (.A_N(_1005_),
    .B(net17),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _1325_ (.A(_1014_),
    .X(\inputs.keypad[8] ));
 sky130_fd_sc_hd__and2b_1 _1326_ (.A_N(_1005_),
    .B(net18),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _1327_ (.A(_1015_),
    .X(\inputs.keypad[9] ));
 sky130_fd_sc_hd__and2b_1 _1328_ (.A_N(net1),
    .B(net3),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _1329_ (.A(_1016_),
    .X(\inputs.keypad[10] ));
 sky130_fd_sc_hd__and2b_1 _1330_ (.A_N(net1),
    .B(net4),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _1331_ (.A(_1017_),
    .X(\inputs.keypad[11] ));
 sky130_fd_sc_hd__and2b_1 _1332_ (.A_N(net1),
    .B(net5),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_1 _1333_ (.A(_1018_),
    .X(\inputs.keypad[12] ));
 sky130_fd_sc_hd__and2b_1 _1334_ (.A_N(net1),
    .B(net9),
    .X(_1019_));
 sky130_fd_sc_hd__clkbuf_1 _1335_ (.A(_1019_),
    .X(\inputs.keypad[13] ));
 sky130_fd_sc_hd__and2b_1 _1336_ (.A_N(net1),
    .B(net6),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_1 _1337_ (.A(_1020_),
    .X(\inputs.keypad[14] ));
 sky130_fd_sc_hd__and2b_1 _1338_ (.A_N(net1),
    .B(net7),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _1339_ (.A(_1021_),
    .X(\inputs.keypad[15] ));
 sky130_fd_sc_hd__and2b_1 _1340_ (.A_N(net1),
    .B(net8),
    .X(_1022_));
 sky130_fd_sc_hd__buf_1 _1341_ (.A(_1022_),
    .X(\inputs.keypad[16] ));
 sky130_fd_sc_hd__and2b_1 _1342_ (.A_N(net1),
    .B(\outputs.pwm_output ),
    .X(_1023_));
 sky130_fd_sc_hd__clkbuf_1 _1343_ (.A(_1023_),
    .X(net20));
 sky130_fd_sc_hd__inv_2 _1344_ (.A(net157),
    .Y(\inputs.random_update_clock.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _1345_ (.A(net174),
    .B(net157),
    .X(\inputs.random_update_clock.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1346_ (.A(\inputs.random_update_clock.count[1] ),
    .B(\inputs.random_update_clock.count[0] ),
    .C(\inputs.random_update_clock.count[2] ),
    .X(_1024_));
 sky130_fd_sc_hd__a21oi_1 _1347_ (.A1(net174),
    .A2(\inputs.random_update_clock.count[0] ),
    .B1(net194),
    .Y(_1025_));
 sky130_fd_sc_hd__nor2_1 _1348_ (.A(_1024_),
    .B(_1025_),
    .Y(\inputs.random_update_clock.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1349_ (.A(\inputs.random_update_clock.count[3] ),
    .B(_1024_),
    .X(_1026_));
 sky130_fd_sc_hd__nor2_1 _1350_ (.A(net198),
    .B(_1024_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_1 _1351_ (.A(_1026_),
    .B(_1027_),
    .Y(\inputs.random_update_clock.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _1352_ (.A(net176),
    .B(_1026_),
    .X(\inputs.random_update_clock.next_count[4] ));
 sky130_fd_sc_hd__a21oi_1 _1353_ (.A1(\inputs.random_update_clock.count[4] ),
    .A2(_1026_),
    .B1(net293),
    .Y(_1028_));
 sky130_fd_sc_hd__and3_1 _1354_ (.A(\inputs.random_update_clock.count[4] ),
    .B(\inputs.random_update_clock.count[5] ),
    .C(_1026_),
    .X(_1029_));
 sky130_fd_sc_hd__or4bb_1 _1355_ (.A(\inputs.random_update_clock.count[4] ),
    .B(\inputs.random_update_clock.count[6] ),
    .C_N(\inputs.random_update_clock.count[7] ),
    .D_N(\inputs.random_update_clock.count[5] ),
    .X(_1030_));
 sky130_fd_sc_hd__or4_1 _1356_ (.A(\inputs.random_update_clock.count[1] ),
    .B(\inputs.random_update_clock.count[0] ),
    .C(\inputs.random_update_clock.count[3] ),
    .D(\inputs.random_update_clock.count[2] ),
    .X(_1031_));
 sky130_fd_sc_hd__nor2_1 _1357_ (.A(_1030_),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__or4b_1 _1358_ (.A(\inputs.random_update_clock.count[12] ),
    .B(\inputs.random_update_clock.count[15] ),
    .C(\inputs.random_update_clock.count[14] ),
    .D_N(\inputs.random_update_clock.count[13] ),
    .X(_1033_));
 sky130_fd_sc_hd__or4bb_1 _1359_ (.A(\inputs.random_update_clock.count[9] ),
    .B(\inputs.random_update_clock.count[11] ),
    .C_N(\inputs.random_update_clock.count[10] ),
    .D_N(\inputs.random_update_clock.count[8] ),
    .X(_1034_));
 sky130_fd_sc_hd__nor2_1 _1360_ (.A(_1033_),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__and4bb_1 _1361_ (.A_N(\inputs.random_update_clock.count[16] ),
    .B_N(\inputs.random_update_clock.count[19] ),
    .C(\inputs.random_update_clock.count[18] ),
    .D(\inputs.random_update_clock.count[17] ),
    .X(_1036_));
 sky130_fd_sc_hd__nor3b_1 _1362_ (.A(\inputs.random_update_clock.count[20] ),
    .B(\inputs.random_update_clock.count[22] ),
    .C_N(\inputs.random_update_clock.count[21] ),
    .Y(_1037_));
 sky130_fd_sc_hd__and4_1 _1363_ (.A(_1032_),
    .B(_1035_),
    .C(_1036_),
    .D(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__buf_2 _1364_ (.A(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__nor3_1 _1365_ (.A(_1028_),
    .B(_1029_),
    .C(_1039_),
    .Y(\inputs.random_update_clock.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _1366_ (.A(\inputs.random_update_clock.count[6] ),
    .B(_1029_),
    .X(_1040_));
 sky130_fd_sc_hd__nor2_1 _1367_ (.A(net216),
    .B(_1029_),
    .Y(_1041_));
 sky130_fd_sc_hd__nor2_1 _1368_ (.A(_1040_),
    .B(_1041_),
    .Y(\inputs.random_update_clock.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _1369_ (.A(\inputs.random_update_clock.count[6] ),
    .B(\inputs.random_update_clock.count[7] ),
    .C(_1029_),
    .X(_1042_));
 sky130_fd_sc_hd__nand4_2 _1370_ (.A(_1032_),
    .B(_1035_),
    .C(_1036_),
    .D(_1037_),
    .Y(_1043_));
 sky130_fd_sc_hd__o21ai_1 _1371_ (.A1(net212),
    .A2(_1040_),
    .B1(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_1 _1372_ (.A(_1042_),
    .B(_1044_),
    .Y(\inputs.random_update_clock.next_count[7] ));
 sky130_fd_sc_hd__nor2_1 _1373_ (.A(\inputs.random_update_clock.count[8] ),
    .B(_1042_),
    .Y(_1045_));
 sky130_fd_sc_hd__and2_1 _1374_ (.A(\inputs.random_update_clock.count[8] ),
    .B(_1042_),
    .X(_1046_));
 sky130_fd_sc_hd__nor3_1 _1375_ (.A(_1039_),
    .B(_1045_),
    .C(_1046_),
    .Y(\inputs.random_update_clock.next_count[8] ));
 sky130_fd_sc_hd__and3_1 _1376_ (.A(\inputs.random_update_clock.count[9] ),
    .B(\inputs.random_update_clock.count[8] ),
    .C(_1042_),
    .X(_1047_));
 sky130_fd_sc_hd__nor2_1 _1377_ (.A(net196),
    .B(_1046_),
    .Y(_1048_));
 sky130_fd_sc_hd__nor2_1 _1378_ (.A(_1047_),
    .B(_1048_),
    .Y(\inputs.random_update_clock.next_count[9] ));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(\inputs.random_update_clock.count[10] ),
    .B(_1047_),
    .Y(_1049_));
 sky130_fd_sc_hd__or2_1 _1380_ (.A(\inputs.random_update_clock.count[10] ),
    .B(_1047_),
    .X(_1050_));
 sky130_fd_sc_hd__and3_1 _1381_ (.A(_1043_),
    .B(_1049_),
    .C(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_1 _1382_ (.A(_1051_),
    .X(\inputs.random_update_clock.next_count[10] ));
 sky130_fd_sc_hd__xnor2_1 _1383_ (.A(net191),
    .B(_1049_),
    .Y(\inputs.random_update_clock.next_count[11] ));
 sky130_fd_sc_hd__and4_1 _1384_ (.A(\inputs.random_update_clock.count[11] ),
    .B(\inputs.random_update_clock.count[10] ),
    .C(\inputs.random_update_clock.count[12] ),
    .D(_1047_),
    .X(_1052_));
 sky130_fd_sc_hd__a31o_1 _1385_ (.A1(\inputs.random_update_clock.count[11] ),
    .A2(\inputs.random_update_clock.count[10] ),
    .A3(_1047_),
    .B1(\inputs.random_update_clock.count[12] ),
    .X(_1053_));
 sky130_fd_sc_hd__and2b_1 _1386_ (.A_N(_1052_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_1 _1387_ (.A(_1054_),
    .X(\inputs.random_update_clock.next_count[12] ));
 sky130_fd_sc_hd__or2_1 _1388_ (.A(\inputs.random_update_clock.count[13] ),
    .B(_1052_),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_1 _1389_ (.A(\inputs.random_update_clock.count[13] ),
    .B(_1052_),
    .Y(_1056_));
 sky130_fd_sc_hd__and3_1 _1390_ (.A(_1043_),
    .B(_1055_),
    .C(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _1391_ (.A(_1057_),
    .X(\inputs.random_update_clock.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _1392_ (.A(\inputs.random_update_clock.count[13] ),
    .B(\inputs.random_update_clock.count[14] ),
    .C(_1052_),
    .X(_1058_));
 sky130_fd_sc_hd__a21oi_1 _1393_ (.A1(\inputs.random_update_clock.count[13] ),
    .A2(_1052_),
    .B1(net166),
    .Y(_1059_));
 sky130_fd_sc_hd__nor2_1 _1394_ (.A(_1058_),
    .B(net167),
    .Y(\inputs.random_update_clock.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _1395_ (.A(\inputs.random_update_clock.count[15] ),
    .B(_1058_),
    .X(_1060_));
 sky130_fd_sc_hd__nor2_1 _1396_ (.A(net187),
    .B(_1058_),
    .Y(_1061_));
 sky130_fd_sc_hd__nor2_1 _1397_ (.A(_1060_),
    .B(_1061_),
    .Y(\inputs.random_update_clock.next_count[15] ));
 sky130_fd_sc_hd__xor2_1 _1398_ (.A(net168),
    .B(_1060_),
    .X(\inputs.random_update_clock.next_count[16] ));
 sky130_fd_sc_hd__a21oi_1 _1399_ (.A1(\inputs.random_update_clock.count[16] ),
    .A2(_1060_),
    .B1(net284),
    .Y(_1062_));
 sky130_fd_sc_hd__and3_1 _1400_ (.A(\inputs.random_update_clock.count[16] ),
    .B(\inputs.random_update_clock.count[17] ),
    .C(_1060_),
    .X(_1063_));
 sky130_fd_sc_hd__nor3_1 _1401_ (.A(_1039_),
    .B(net285),
    .C(_1063_),
    .Y(\inputs.random_update_clock.next_count[17] ));
 sky130_fd_sc_hd__nor2_1 _1402_ (.A(net307),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__and2_1 _1403_ (.A(\inputs.random_update_clock.count[18] ),
    .B(_1063_),
    .X(_1065_));
 sky130_fd_sc_hd__nor3_1 _1404_ (.A(_1039_),
    .B(_1064_),
    .C(_1065_),
    .Y(\inputs.random_update_clock.next_count[18] ));
 sky130_fd_sc_hd__xor2_1 _1405_ (.A(net190),
    .B(_1065_),
    .X(\inputs.random_update_clock.next_count[19] ));
 sky130_fd_sc_hd__and3_1 _1406_ (.A(\inputs.random_update_clock.count[19] ),
    .B(\inputs.random_update_clock.count[20] ),
    .C(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__a21oi_1 _1407_ (.A1(\inputs.random_update_clock.count[19] ),
    .A2(_1065_),
    .B1(net177),
    .Y(_1067_));
 sky130_fd_sc_hd__nor2_1 _1408_ (.A(_1066_),
    .B(net178),
    .Y(\inputs.random_update_clock.next_count[20] ));
 sky130_fd_sc_hd__or2_1 _1409_ (.A(\inputs.random_update_clock.count[21] ),
    .B(_1066_),
    .X(_1068_));
 sky130_fd_sc_hd__nand2_1 _1410_ (.A(\inputs.random_update_clock.count[21] ),
    .B(_1066_),
    .Y(_1069_));
 sky130_fd_sc_hd__and3_1 _1411_ (.A(_1043_),
    .B(_1068_),
    .C(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__clkbuf_1 _1412_ (.A(_1070_),
    .X(\inputs.random_update_clock.next_count[21] ));
 sky130_fd_sc_hd__xnor2_1 _1413_ (.A(net96),
    .B(_1069_),
    .Y(\inputs.random_update_clock.next_count[22] ));
 sky130_fd_sc_hd__nor3b_1 _1414_ (.A(net94),
    .B(net88),
    .C_N(\inputs.key_encoder.sync_keys[14] ),
    .Y(\inputs.key_encoder.mode_key ));
 sky130_fd_sc_hd__and2b_1 _1415_ (.A_N(\inputs.key_encoder.octave_key_up ),
    .B(\inputs.key_encoder.sync_keys[15] ),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _1416_ (.A(_1071_),
    .X(\inputs.down.in ));
 sky130_fd_sc_hd__inv_2 _1417_ (.A(net90),
    .Y(\outputs.output_gen.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _1418_ (.A(\outputs.output_gen.count[1] ),
    .B(net90),
    .X(\outputs.output_gen.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1419_ (.A(\outputs.output_gen.count[2] ),
    .B(\outputs.output_gen.count[1] ),
    .C(\outputs.output_gen.count[0] ),
    .X(_1072_));
 sky130_fd_sc_hd__a21oi_1 _1420_ (.A1(\outputs.output_gen.count[1] ),
    .A2(net90),
    .B1(net218),
    .Y(_1073_));
 sky130_fd_sc_hd__nor2_1 _1421_ (.A(_1072_),
    .B(net219),
    .Y(\outputs.output_gen.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1422_ (.A(\outputs.output_gen.count[3] ),
    .B(_1072_),
    .X(_1074_));
 sky130_fd_sc_hd__nor2_1 _1423_ (.A(net268),
    .B(_1072_),
    .Y(_1075_));
 sky130_fd_sc_hd__nor2_1 _1424_ (.A(_1074_),
    .B(_1075_),
    .Y(\outputs.output_gen.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _1425_ (.A(net236),
    .B(_1074_),
    .X(\outputs.output_gen.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1426_ (.A(\outputs.output_gen.count[5] ),
    .B(\outputs.output_gen.count[4] ),
    .C(_1074_),
    .X(_1076_));
 sky130_fd_sc_hd__a21oi_1 _1427_ (.A1(net314),
    .A2(_1074_),
    .B1(net227),
    .Y(_1077_));
 sky130_fd_sc_hd__nor2_1 _1428_ (.A(_1076_),
    .B(_1077_),
    .Y(\outputs.output_gen.next_count[5] ));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(\outputs.output_gen.count[6] ),
    .B(_1076_),
    .Y(_1078_));
 sky130_fd_sc_hd__or2_1 _1430_ (.A(\outputs.output_gen.count[6] ),
    .B(_1076_),
    .X(_1079_));
 sky130_fd_sc_hd__and2_1 _1431_ (.A(_1078_),
    .B(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _1432_ (.A(_1080_),
    .X(\outputs.output_gen.next_count[6] ));
 sky130_fd_sc_hd__xnor2_1 _1433_ (.A(net148),
    .B(_1078_),
    .Y(\outputs.output_gen.next_count[7] ));
 sky130_fd_sc_hd__and3_1 _1434_ (.A(\outputs.sample_rate.count[6] ),
    .B(\outputs.sample_rate.count[7] ),
    .C(_0996_),
    .X(_1081_));
 sky130_fd_sc_hd__nor2_1 _1435_ (.A(_1081_),
    .B(_1001_),
    .Y(_1082_));
 sky130_fd_sc_hd__buf_2 _1436_ (.A(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__clkbuf_4 _1437_ (.A(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_4 _1438_ (.A(_1084_),
    .X(\outputs.div.next_div ));
 sky130_fd_sc_hd__inv_2 _1439_ (.A(net100),
    .Y(\outputs.sample_rate.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _1440_ (.A(net114),
    .B(net100),
    .X(\outputs.sample_rate.next_count[1] ));
 sky130_fd_sc_hd__a21oi_1 _1441_ (.A1(\outputs.sample_rate.count[1] ),
    .A2(\outputs.sample_rate.count[0] ),
    .B1(net112),
    .Y(_1085_));
 sky130_fd_sc_hd__nor2_1 _1442_ (.A(_0994_),
    .B(net113),
    .Y(\outputs.sample_rate.next_count[2] ));
 sky130_fd_sc_hd__nor2_1 _1443_ (.A(net145),
    .B(_0994_),
    .Y(_1086_));
 sky130_fd_sc_hd__nor2_1 _1444_ (.A(_0995_),
    .B(_1086_),
    .Y(\outputs.sample_rate.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _1445_ (.A(net141),
    .B(_0995_),
    .X(\outputs.sample_rate.next_count[4] ));
 sky130_fd_sc_hd__a21oi_1 _1446_ (.A1(\outputs.sample_rate.count[4] ),
    .A2(_0995_),
    .B1(net131),
    .Y(_1087_));
 sky130_fd_sc_hd__nor2_1 _1447_ (.A(_0996_),
    .B(net132),
    .Y(\outputs.sample_rate.next_count[5] ));
 sky130_fd_sc_hd__nor2_1 _1448_ (.A(net180),
    .B(_0996_),
    .Y(_1088_));
 sky130_fd_sc_hd__nor2_1 _1449_ (.A(_0997_),
    .B(_1088_),
    .Y(\outputs.sample_rate.next_count[6] ));
 sky130_fd_sc_hd__clkbuf_4 _1450_ (.A(_1081_),
    .X(_1089_));
 sky130_fd_sc_hd__clkbuf_4 _1451_ (.A(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__nor2_1 _1452_ (.A(net204),
    .B(_0997_),
    .Y(_1091_));
 sky130_fd_sc_hd__nor2_1 _1453_ (.A(_1090_),
    .B(_1091_),
    .Y(\outputs.sample_rate.next_count[7] ));
 sky130_fd_sc_hd__inv_2 _1454_ (.A(\outputs.divider_buffer[1] ),
    .Y(_1092_));
 sky130_fd_sc_hd__inv_2 _1455_ (.A(\outputs.sig_gen.count[13] ),
    .Y(_1093_));
 sky130_fd_sc_hd__a2bb2o_1 _1456_ (.A1_N(_1092_),
    .A2_N(\outputs.sig_gen.count[1] ),
    .B1(\outputs.divider_buffer[13] ),
    .B2(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__inv_2 _1457_ (.A(\outputs.divider_buffer[9] ),
    .Y(_1095_));
 sky130_fd_sc_hd__inv_2 _1458_ (.A(\outputs.divider_buffer[17] ),
    .Y(_1096_));
 sky130_fd_sc_hd__xor2_1 _1459_ (.A(\outputs.divider_buffer[12] ),
    .B(\outputs.sig_gen.count[12] ),
    .X(_1097_));
 sky130_fd_sc_hd__a221o_1 _1460_ (.A1(_1095_),
    .A2(\outputs.sig_gen.count[9] ),
    .B1(_1096_),
    .B2(\outputs.sig_gen.count[17] ),
    .C1(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__inv_2 _1461_ (.A(\outputs.sig_gen.count[3] ),
    .Y(_1099_));
 sky130_fd_sc_hd__inv_2 _1462_ (.A(\outputs.sig_gen.count[9] ),
    .Y(_1100_));
 sky130_fd_sc_hd__xor2_1 _1463_ (.A(\outputs.divider_buffer[4] ),
    .B(\outputs.sig_gen.count[4] ),
    .X(_1101_));
 sky130_fd_sc_hd__a221o_1 _1464_ (.A1(\outputs.divider_buffer[3] ),
    .A2(_1099_),
    .B1(\outputs.divider_buffer[9] ),
    .B2(_1100_),
    .C1(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__inv_2 _1465_ (.A(\outputs.divider_buffer[10] ),
    .Y(_1103_));
 sky130_fd_sc_hd__a2bb2o_1 _1466_ (.A1_N(_1103_),
    .A2_N(\outputs.sig_gen.count[10] ),
    .B1(_1092_),
    .B2(\outputs.sig_gen.count[1] ),
    .X(_1104_));
 sky130_fd_sc_hd__or4_1 _1467_ (.A(_1094_),
    .B(_1098_),
    .C(_1102_),
    .D(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__inv_2 _1468_ (.A(\outputs.divider_buffer[3] ),
    .Y(_1106_));
 sky130_fd_sc_hd__inv_2 _1469_ (.A(\outputs.divider_buffer[15] ),
    .Y(_1107_));
 sky130_fd_sc_hd__inv_2 _1470_ (.A(\outputs.divider_buffer[5] ),
    .Y(_1108_));
 sky130_fd_sc_hd__o22ai_1 _1471_ (.A1(_1108_),
    .A2(\outputs.sig_gen.count[5] ),
    .B1(_1096_),
    .B2(\outputs.sig_gen.count[17] ),
    .Y(_1109_));
 sky130_fd_sc_hd__a221o_1 _1472_ (.A1(_1106_),
    .A2(\outputs.sig_gen.count[3] ),
    .B1(_1107_),
    .B2(\outputs.sig_gen.count[15] ),
    .C1(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__inv_2 _1473_ (.A(\outputs.divider_buffer[14] ),
    .Y(_1111_));
 sky130_fd_sc_hd__inv_2 _1474_ (.A(\outputs.sig_gen.count[16] ),
    .Y(_1112_));
 sky130_fd_sc_hd__xor2_1 _1475_ (.A(\outputs.divider_buffer[2] ),
    .B(\outputs.sig_gen.count[2] ),
    .X(_1113_));
 sky130_fd_sc_hd__a221o_1 _1476_ (.A1(_1111_),
    .A2(\outputs.sig_gen.count[14] ),
    .B1(\outputs.divider_buffer[16] ),
    .B2(_1112_),
    .C1(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__inv_2 _1477_ (.A(\outputs.sig_gen.count[7] ),
    .Y(_1115_));
 sky130_fd_sc_hd__inv_2 _1478_ (.A(\outputs.sig_gen.count[11] ),
    .Y(_1116_));
 sky130_fd_sc_hd__xor2_1 _1479_ (.A(\outputs.divider_buffer[8] ),
    .B(\outputs.sig_gen.count[8] ),
    .X(_1117_));
 sky130_fd_sc_hd__a221o_1 _1480_ (.A1(\outputs.divider_buffer[7] ),
    .A2(_1115_),
    .B1(\outputs.divider_buffer[11] ),
    .B2(_1116_),
    .C1(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__inv_2 _1481_ (.A(\outputs.divider_buffer[6] ),
    .Y(_1119_));
 sky130_fd_sc_hd__o22a_1 _1482_ (.A1(_1119_),
    .A2(\outputs.sig_gen.count[6] ),
    .B1(\outputs.divider_buffer[16] ),
    .B2(_1112_),
    .X(_1120_));
 sky130_fd_sc_hd__o221ai_1 _1483_ (.A1(\outputs.divider_buffer[13] ),
    .A2(_1093_),
    .B1(_1111_),
    .B2(\outputs.sig_gen.count[14] ),
    .C1(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__inv_2 _1484_ (.A(\outputs.divider_buffer[0] ),
    .Y(_1122_));
 sky130_fd_sc_hd__inv_2 _1485_ (.A(\outputs.divider_buffer[11] ),
    .Y(_1123_));
 sky130_fd_sc_hd__a2bb2o_1 _1486_ (.A1_N(_1122_),
    .A2_N(\outputs.sig_gen.count[0] ),
    .B1(_1108_),
    .B2(\outputs.sig_gen.count[5] ),
    .X(_1124_));
 sky130_fd_sc_hd__a221o_1 _1487_ (.A1(_1122_),
    .A2(\outputs.sig_gen.count[0] ),
    .B1(_1123_),
    .B2(\outputs.sig_gen.count[11] ),
    .C1(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__inv_2 _1488_ (.A(\outputs.divider_buffer[7] ),
    .Y(_1126_));
 sky130_fd_sc_hd__a2bb2o_1 _1489_ (.A1_N(_1107_),
    .A2_N(\outputs.sig_gen.count[15] ),
    .B1(_1119_),
    .B2(\outputs.sig_gen.count[6] ),
    .X(_1127_));
 sky130_fd_sc_hd__a221o_1 _1490_ (.A1(_1126_),
    .A2(\outputs.sig_gen.count[7] ),
    .B1(_1103_),
    .B2(\outputs.sig_gen.count[10] ),
    .C1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__or4_1 _1491_ (.A(_1118_),
    .B(_1121_),
    .C(_1125_),
    .D(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__or4_4 _1492_ (.A(_1105_),
    .B(_1110_),
    .C(_1114_),
    .D(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__buf_2 _1493_ (.A(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(net193),
    .B(_1131_),
    .Y(\outputs.sig_gen.next_count[0] ));
 sky130_fd_sc_hd__or2_1 _1495_ (.A(\outputs.sig_gen.count[0] ),
    .B(\outputs.sig_gen.count[1] ),
    .X(_1132_));
 sky130_fd_sc_hd__nand2_1 _1496_ (.A(\outputs.sig_gen.count[0] ),
    .B(\outputs.sig_gen.count[1] ),
    .Y(_1133_));
 sky130_fd_sc_hd__and3_1 _1497_ (.A(_1131_),
    .B(_1132_),
    .C(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _1498_ (.A(_1134_),
    .X(\outputs.sig_gen.next_count[1] ));
 sky130_fd_sc_hd__a21o_1 _1499_ (.A1(\outputs.sig_gen.count[0] ),
    .A2(\outputs.sig_gen.count[1] ),
    .B1(\outputs.sig_gen.count[2] ),
    .X(_1135_));
 sky130_fd_sc_hd__nand3_1 _1500_ (.A(\outputs.sig_gen.count[0] ),
    .B(\outputs.sig_gen.count[1] ),
    .C(\outputs.sig_gen.count[2] ),
    .Y(_1136_));
 sky130_fd_sc_hd__and3_1 _1501_ (.A(_1130_),
    .B(_1135_),
    .C(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _1502_ (.A(_1137_),
    .X(\outputs.sig_gen.next_count[2] ));
 sky130_fd_sc_hd__nor2_1 _1503_ (.A(_1099_),
    .B(_1136_),
    .Y(_1138_));
 sky130_fd_sc_hd__inv_2 _1504_ (.A(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__nand2_1 _1505_ (.A(_1099_),
    .B(_1136_),
    .Y(_1140_));
 sky130_fd_sc_hd__and3_1 _1506_ (.A(_1130_),
    .B(_1139_),
    .C(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _1507_ (.A(_1141_),
    .X(\outputs.sig_gen.next_count[3] ));
 sky130_fd_sc_hd__and2_1 _1508_ (.A(\outputs.sig_gen.count[4] ),
    .B(_1138_),
    .X(_1142_));
 sky130_fd_sc_hd__o21ai_1 _1509_ (.A1(net290),
    .A2(_1138_),
    .B1(_1131_),
    .Y(_1143_));
 sky130_fd_sc_hd__nor2_1 _1510_ (.A(_1142_),
    .B(_1143_),
    .Y(\outputs.sig_gen.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1511_ (.A(\outputs.sig_gen.count[4] ),
    .B(\outputs.sig_gen.count[5] ),
    .C(_1138_),
    .X(_1144_));
 sky130_fd_sc_hd__o21ai_1 _1512_ (.A1(\outputs.sig_gen.count[5] ),
    .A2(_1142_),
    .B1(_1131_),
    .Y(_1145_));
 sky130_fd_sc_hd__nor2_1 _1513_ (.A(_1144_),
    .B(_1145_),
    .Y(\outputs.sig_gen.next_count[5] ));
 sky130_fd_sc_hd__or2_1 _1514_ (.A(\outputs.sig_gen.count[6] ),
    .B(_1144_),
    .X(_1146_));
 sky130_fd_sc_hd__and2_1 _1515_ (.A(\outputs.sig_gen.count[6] ),
    .B(_1144_),
    .X(_1147_));
 sky130_fd_sc_hd__inv_2 _1516_ (.A(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__and3_1 _1517_ (.A(_1130_),
    .B(_1146_),
    .C(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__clkbuf_1 _1518_ (.A(_1149_),
    .X(\outputs.sig_gen.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _1519_ (.A(\outputs.sig_gen.count[6] ),
    .B(\outputs.sig_gen.count[7] ),
    .C(_1144_),
    .X(_1150_));
 sky130_fd_sc_hd__o21ai_1 _1520_ (.A1(\outputs.sig_gen.count[7] ),
    .A2(_1147_),
    .B1(_1131_),
    .Y(_1151_));
 sky130_fd_sc_hd__nor2_1 _1521_ (.A(_1150_),
    .B(_1151_),
    .Y(\outputs.sig_gen.next_count[7] ));
 sky130_fd_sc_hd__or2_1 _1522_ (.A(\outputs.sig_gen.count[8] ),
    .B(_1150_),
    .X(_1152_));
 sky130_fd_sc_hd__and2_1 _1523_ (.A(\outputs.sig_gen.count[8] ),
    .B(_1150_),
    .X(_1153_));
 sky130_fd_sc_hd__inv_2 _1524_ (.A(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__and3_1 _1525_ (.A(_1130_),
    .B(_1152_),
    .C(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__clkbuf_1 _1526_ (.A(_1155_),
    .X(\outputs.sig_gen.next_count[8] ));
 sky130_fd_sc_hd__or2_1 _1527_ (.A(\outputs.sig_gen.count[9] ),
    .B(_1153_),
    .X(_1156_));
 sky130_fd_sc_hd__o211a_1 _1528_ (.A1(_1100_),
    .A2(_1154_),
    .B1(_1156_),
    .C1(_1131_),
    .X(\outputs.sig_gen.next_count[9] ));
 sky130_fd_sc_hd__nor2_1 _1529_ (.A(_1100_),
    .B(_1154_),
    .Y(_1157_));
 sky130_fd_sc_hd__or2_1 _1530_ (.A(\outputs.sig_gen.count[10] ),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__nand2_1 _1531_ (.A(\outputs.sig_gen.count[10] ),
    .B(_1157_),
    .Y(_1159_));
 sky130_fd_sc_hd__and3_1 _1532_ (.A(_1130_),
    .B(_1158_),
    .C(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__clkbuf_1 _1533_ (.A(_1160_),
    .X(\outputs.sig_gen.next_count[10] ));
 sky130_fd_sc_hd__nand2_1 _1534_ (.A(_1116_),
    .B(_1159_),
    .Y(_1161_));
 sky130_fd_sc_hd__o211a_1 _1535_ (.A1(_1116_),
    .A2(_1159_),
    .B1(_1161_),
    .C1(_1131_),
    .X(\outputs.sig_gen.next_count[11] ));
 sky130_fd_sc_hd__nor2_1 _1536_ (.A(_1116_),
    .B(_1159_),
    .Y(_1162_));
 sky130_fd_sc_hd__or2_1 _1537_ (.A(\outputs.sig_gen.count[12] ),
    .B(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__and2_1 _1538_ (.A(\outputs.sig_gen.count[12] ),
    .B(_1162_),
    .X(_1164_));
 sky130_fd_sc_hd__inv_2 _1539_ (.A(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__and3_1 _1540_ (.A(_1130_),
    .B(_1163_),
    .C(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_1166_),
    .X(\outputs.sig_gen.next_count[12] ));
 sky130_fd_sc_hd__or2_1 _1542_ (.A(\outputs.sig_gen.count[13] ),
    .B(_1164_),
    .X(_1167_));
 sky130_fd_sc_hd__nand2_1 _1543_ (.A(\outputs.sig_gen.count[13] ),
    .B(_1164_),
    .Y(_1168_));
 sky130_fd_sc_hd__and3_1 _1544_ (.A(_1130_),
    .B(_1167_),
    .C(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__clkbuf_1 _1545_ (.A(_1169_),
    .X(\outputs.sig_gen.next_count[13] ));
 sky130_fd_sc_hd__inv_2 _1546_ (.A(\outputs.sig_gen.count[14] ),
    .Y(_1170_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(_1170_),
    .B(_1168_),
    .Y(_1171_));
 sky130_fd_sc_hd__o211a_1 _1548_ (.A1(_1170_),
    .A2(_1168_),
    .B1(_1171_),
    .C1(_1131_),
    .X(\outputs.sig_gen.next_count[14] ));
 sky130_fd_sc_hd__nor2_1 _1549_ (.A(_1170_),
    .B(_1168_),
    .Y(_1172_));
 sky130_fd_sc_hd__or2_1 _1550_ (.A(\outputs.sig_gen.count[15] ),
    .B(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__nand2_1 _1551_ (.A(\outputs.sig_gen.count[15] ),
    .B(_1172_),
    .Y(_1174_));
 sky130_fd_sc_hd__and3_1 _1552_ (.A(_1130_),
    .B(_1173_),
    .C(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _1553_ (.A(_1175_),
    .X(\outputs.sig_gen.next_count[15] ));
 sky130_fd_sc_hd__nand2_1 _1554_ (.A(_1112_),
    .B(_1174_),
    .Y(_1176_));
 sky130_fd_sc_hd__o211a_1 _1555_ (.A1(_1112_),
    .A2(_1174_),
    .B1(_1176_),
    .C1(_1131_),
    .X(\outputs.sig_gen.next_count[16] ));
 sky130_fd_sc_hd__nor2_1 _1556_ (.A(_1112_),
    .B(_1174_),
    .Y(_1177_));
 sky130_fd_sc_hd__o21ai_1 _1557_ (.A1(net186),
    .A2(_1177_),
    .B1(_1131_),
    .Y(_1178_));
 sky130_fd_sc_hd__a21oi_1 _1558_ (.A1(net186),
    .A2(_1177_),
    .B1(_1178_),
    .Y(\outputs.sig_gen.next_count[17] ));
 sky130_fd_sc_hd__nand2_1 _1559_ (.A(\inputs.wavetype_fsm.state[0] ),
    .B(\inputs.mode_edge.det_edge ),
    .Y(_1179_));
 sky130_fd_sc_hd__or2_1 _1560_ (.A(\inputs.wavetype_fsm.state[0] ),
    .B(\inputs.mode_edge.det_edge ),
    .X(_1180_));
 sky130_fd_sc_hd__and2_1 _1561_ (.A(_1179_),
    .B(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__clkbuf_1 _1562_ (.A(_1181_),
    .X(\inputs.wavetype_fsm.next_state[0] ));
 sky130_fd_sc_hd__xnor2_1 _1563_ (.A(net183),
    .B(_1179_),
    .Y(\inputs.wavetype_fsm.next_state[1] ));
 sky130_fd_sc_hd__buf_2 _1564_ (.A(\inputs.random_note_generator.out[15] ),
    .X(_1182_));
 sky130_fd_sc_hd__xor2_1 _1565_ (.A(_1182_),
    .B(\inputs.random_note_generator.out[13] ),
    .X(_1183_));
 sky130_fd_sc_hd__xor2_1 _1566_ (.A(net319),
    .B(\inputs.random_note_generator.out[10] ),
    .X(_1184_));
 sky130_fd_sc_hd__xnor2_1 _1567_ (.A(_1183_),
    .B(_1184_),
    .Y(\inputs.random_note_generator.feedback ));
 sky130_fd_sc_hd__or2b_1 _1568_ (.A(net115),
    .B_N(\inputs.key_encoder.mode_key ),
    .X(_1185_));
 sky130_fd_sc_hd__inv_2 _1569_ (.A(_1185_),
    .Y(\inputs.mode_edge.ff_in ));
 sky130_fd_sc_hd__and2b_1 _1570_ (.A_N(net296),
    .B(\inputs.down.in ),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_1 _1571_ (.A(_1186_),
    .X(\inputs.down.ff_in ));
 sky130_fd_sc_hd__and2b_1 _1572_ (.A_N(net305),
    .B(\inputs.key_encoder.octave_key_up ),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_1 _1573_ (.A(_1187_),
    .X(\inputs.up.ff_in ));
 sky130_fd_sc_hd__or4_2 _1574_ (.A(\outputs.scaled_buffer[0] ),
    .B(\outputs.scaled_buffer[1] ),
    .C(\outputs.scaled_buffer[3] ),
    .D(\outputs.scaled_buffer[2] ),
    .X(_1188_));
 sky130_fd_sc_hd__and2_1 _1575_ (.A(_1111_),
    .B(\outputs.shaper.count[13] ),
    .X(_1189_));
 sky130_fd_sc_hd__inv_2 _1576_ (.A(\outputs.shaper.count[14] ),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _1577_ (.A(\outputs.divider_buffer[15] ),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__inv_2 _1578_ (.A(\outputs.divider_buffer[16] ),
    .Y(_1192_));
 sky130_fd_sc_hd__a2bb2o_1 _1579_ (.A1_N(_1192_),
    .A2_N(\outputs.shaper.count[15] ),
    .B1(_1190_),
    .B2(\outputs.divider_buffer[15] ),
    .X(_1193_));
 sky130_fd_sc_hd__nand2_1 _1580_ (.A(_1192_),
    .B(\outputs.shaper.count[15] ),
    .Y(_1194_));
 sky130_fd_sc_hd__or3b_1 _1581_ (.A(_1191_),
    .B(_1193_),
    .C_N(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__inv_2 _1582_ (.A(\outputs.shaper.count[9] ),
    .Y(_1196_));
 sky130_fd_sc_hd__a2bb2o_1 _1583_ (.A1_N(_1095_),
    .A2_N(\outputs.shaper.count[8] ),
    .B1(\outputs.divider_buffer[10] ),
    .B2(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__a21o_1 _1584_ (.A1(_1095_),
    .A2(\outputs.shaper.count[8] ),
    .B1(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__inv_2 _1585_ (.A(\outputs.shaper.count[12] ),
    .Y(_1199_));
 sky130_fd_sc_hd__a2bb2o_1 _1586_ (.A1_N(_1111_),
    .A2_N(\outputs.shaper.count[13] ),
    .B1(_1199_),
    .B2(\outputs.divider_buffer[13] ),
    .X(_1200_));
 sky130_fd_sc_hd__inv_2 _1587_ (.A(\outputs.shaper.count[11] ),
    .Y(_1201_));
 sky130_fd_sc_hd__inv_2 _1588_ (.A(\outputs.shaper.count[10] ),
    .Y(_1202_));
 sky130_fd_sc_hd__a22o_1 _1589_ (.A1(\outputs.divider_buffer[12] ),
    .A2(_1201_),
    .B1(_1202_),
    .B2(\outputs.divider_buffer[11] ),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_1 _1590_ (.A(\outputs.divider_buffer[10] ),
    .B(_1196_),
    .Y(_1204_));
 sky130_fd_sc_hd__nor2_1 _1591_ (.A(\outputs.divider_buffer[11] ),
    .B(_1202_),
    .Y(_1205_));
 sky130_fd_sc_hd__nor2_1 _1592_ (.A(\outputs.divider_buffer[12] ),
    .B(_1201_),
    .Y(_1206_));
 sky130_fd_sc_hd__nor2_1 _1593_ (.A(\outputs.divider_buffer[13] ),
    .B(_1199_),
    .Y(_1207_));
 sky130_fd_sc_hd__or4_1 _1594_ (.A(_1204_),
    .B(_1205_),
    .C(_1206_),
    .D(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__or4_1 _1595_ (.A(_1198_),
    .B(_1200_),
    .C(_1203_),
    .D(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__or3_1 _1596_ (.A(_1189_),
    .B(_1195_),
    .C(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__inv_2 _1597_ (.A(\outputs.shaper.count[7] ),
    .Y(_1211_));
 sky130_fd_sc_hd__or2_1 _1598_ (.A(\outputs.divider_buffer[8] ),
    .B(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__inv_2 _1599_ (.A(\outputs.shaper.count[3] ),
    .Y(_1213_));
 sky130_fd_sc_hd__inv_2 _1600_ (.A(\outputs.shaper.count[2] ),
    .Y(_1214_));
 sky130_fd_sc_hd__a22o_1 _1601_ (.A1(\outputs.divider_buffer[4] ),
    .A2(_1213_),
    .B1(_1214_),
    .B2(\outputs.divider_buffer[3] ),
    .X(_1215_));
 sky130_fd_sc_hd__or2b_1 _1602_ (.A(\outputs.shaper.count[1] ),
    .B_N(\outputs.divider_buffer[2] ),
    .X(_1216_));
 sky130_fd_sc_hd__inv_2 _1603_ (.A(\outputs.shaper.count[0] ),
    .Y(_1217_));
 sky130_fd_sc_hd__or2b_1 _1604_ (.A(\outputs.divider_buffer[2] ),
    .B_N(\outputs.shaper.count[1] ),
    .X(_1218_));
 sky130_fd_sc_hd__o211ai_1 _1605_ (.A1(\outputs.divider_buffer[1] ),
    .A2(_1217_),
    .B1(_1216_),
    .C1(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__nor2_1 _1606_ (.A(\outputs.divider_buffer[3] ),
    .B(_1214_),
    .Y(_1220_));
 sky130_fd_sc_hd__a21oi_1 _1607_ (.A1(_1216_),
    .A2(_1219_),
    .B1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__or2_1 _1608_ (.A(_1215_),
    .B(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__or2_1 _1609_ (.A(\outputs.divider_buffer[4] ),
    .B(_1213_),
    .X(_1223_));
 sky130_fd_sc_hd__nand2_1 _1610_ (.A(_1108_),
    .B(\outputs.shaper.count[4] ),
    .Y(_1224_));
 sky130_fd_sc_hd__o22ai_1 _1611_ (.A1(_1119_),
    .A2(\outputs.shaper.count[5] ),
    .B1(\outputs.shaper.count[4] ),
    .B2(_1108_),
    .Y(_1225_));
 sky130_fd_sc_hd__a31o_1 _1612_ (.A1(_1222_),
    .A2(_1223_),
    .A3(_1224_),
    .B1(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__nand2_1 _1613_ (.A(_1119_),
    .B(\outputs.shaper.count[5] ),
    .Y(_1227_));
 sky130_fd_sc_hd__nand2_1 _1614_ (.A(_1126_),
    .B(\outputs.shaper.count[6] ),
    .Y(_1228_));
 sky130_fd_sc_hd__a2bb2o_1 _1615_ (.A1_N(_1126_),
    .A2_N(\outputs.shaper.count[6] ),
    .B1(\outputs.divider_buffer[8] ),
    .B2(_1211_),
    .X(_1229_));
 sky130_fd_sc_hd__a31o_1 _1616_ (.A1(_1226_),
    .A2(_1227_),
    .A3(_1228_),
    .B1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__and3b_1 _1617_ (.A_N(_1210_),
    .B(_1212_),
    .C(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__nor2_1 _1618_ (.A(_1204_),
    .B(_1205_),
    .Y(_1232_));
 sky130_fd_sc_hd__a21oi_1 _1619_ (.A1(_1197_),
    .A2(_1232_),
    .B1(_1203_),
    .Y(_1233_));
 sky130_fd_sc_hd__inv_2 _1620_ (.A(_1200_),
    .Y(_1234_));
 sky130_fd_sc_hd__o31a_1 _1621_ (.A1(_1206_),
    .A2(_1207_),
    .A3(_1233_),
    .B1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__o2bb2a_1 _1622_ (.A1_N(_1193_),
    .A2_N(_1194_),
    .B1(_1096_),
    .B2(\outputs.shaper.count[16] ),
    .X(_1236_));
 sky130_fd_sc_hd__o31ai_1 _1623_ (.A1(_1189_),
    .A2(_1195_),
    .A3(_1235_),
    .B1(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__a21oi_1 _1624_ (.A1(_1096_),
    .A2(\outputs.shaper.count[16] ),
    .B1(\outputs.shaper.count[17] ),
    .Y(_1238_));
 sky130_fd_sc_hd__or4b_1 _1625_ (.A(_1229_),
    .B(_1225_),
    .C(_1215_),
    .D_N(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__o22a_1 _1626_ (.A1(_1096_),
    .A2(\outputs.shaper.count[16] ),
    .B1(\outputs.shaper.count[0] ),
    .B2(_1092_),
    .X(_1240_));
 sky130_fd_sc_hd__and4b_1 _1627_ (.A_N(_1220_),
    .B(_1223_),
    .C(_1228_),
    .D(_1212_),
    .X(_1241_));
 sky130_fd_sc_hd__and4_1 _1628_ (.A(_1224_),
    .B(_1227_),
    .C(_1240_),
    .D(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__or4b_1 _1629_ (.A(_1219_),
    .B(_1210_),
    .C(_1239_),
    .D_N(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__o211ai_1 _1630_ (.A1(_1231_),
    .A2(_1237_),
    .B1(_1238_),
    .C1(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__a21oi_1 _1631_ (.A1(_1188_),
    .A2(net21),
    .B1(\outputs.scaled_buffer[4] ),
    .Y(_1245_));
 sky130_fd_sc_hd__nor2b_4 _1632_ (.A(\inputs.wavetype_fsm.state[1] ),
    .B_N(\inputs.wavetype_fsm.state[0] ),
    .Y(_1246_));
 sky130_fd_sc_hd__inv_2 _1633_ (.A(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__a31o_1 _1634_ (.A1(\outputs.scaled_buffer[4] ),
    .A2(_1188_),
    .A3(net21),
    .B1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__and2b_1 _1635_ (.A_N(\inputs.wavetype_fsm.state[0] ),
    .B(\inputs.wavetype_fsm.state[1] ),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_4 _1636_ (.A(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__nand2_1 _1637_ (.A(\inputs.wavetype_fsm.state[0] ),
    .B(\inputs.wavetype_fsm.state[1] ),
    .Y(_1251_));
 sky130_fd_sc_hd__or3_1 _1638_ (.A(\outputs.scaled_buffer[5] ),
    .B(\outputs.scaled_buffer[4] ),
    .C(_1188_),
    .X(_1252_));
 sky130_fd_sc_hd__or4b_2 _1639_ (.A(\outputs.scaled_buffer[6] ),
    .B(_1247_),
    .C(_1252_),
    .D_N(\outputs.scaled_buffer[7] ),
    .X(_1253_));
 sky130_fd_sc_hd__o21ai_4 _1640_ (.A1(net21),
    .A2(_1251_),
    .B1(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__a21oi_1 _1641_ (.A1(\outputs.scaled_buffer[5] ),
    .A2(_1250_),
    .B1(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__o21a_1 _1642_ (.A1(_1245_),
    .A2(_1248_),
    .B1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__o21ai_1 _1643_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(\outputs.scaled_buffer[1] ),
    .B1(net21),
    .Y(_1257_));
 sky130_fd_sc_hd__xnor2_1 _1644_ (.A(\outputs.scaled_buffer[2] ),
    .B(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__a221oi_2 _1645_ (.A1(\outputs.scaled_buffer[3] ),
    .A2(_1250_),
    .B1(_1258_),
    .B2(_1246_),
    .C1(_1254_),
    .Y(_1259_));
 sky130_fd_sc_hd__a21oi_1 _1646_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(net21),
    .B1(\outputs.scaled_buffer[1] ),
    .Y(_1260_));
 sky130_fd_sc_hd__a31o_1 _1647_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(\outputs.scaled_buffer[1] ),
    .A3(net21),
    .B1(_1247_),
    .X(_1261_));
 sky130_fd_sc_hd__a21oi_1 _1648_ (.A1(\outputs.scaled_buffer[2] ),
    .A2(_1250_),
    .B1(_1254_),
    .Y(_1262_));
 sky130_fd_sc_hd__o21a_1 _1649_ (.A1(_1260_),
    .A2(_1261_),
    .B1(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__a221oi_2 _1650_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(_1246_),
    .B1(_1250_),
    .B2(\outputs.scaled_buffer[1] ),
    .C1(_1254_),
    .Y(_1264_));
 sky130_fd_sc_hd__or2_1 _1651_ (.A(\outputs.output_gen.count[1] ),
    .B(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__a21oi_1 _1652_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(_1250_),
    .B1(_1254_),
    .Y(_1266_));
 sky130_fd_sc_hd__a211o_1 _1653_ (.A1(\outputs.output_gen.count[1] ),
    .A2(_1264_),
    .B1(_1266_),
    .C1(\outputs.output_gen.count[0] ),
    .X(_1267_));
 sky130_fd_sc_hd__a22o_1 _1654_ (.A1(\outputs.output_gen.count[2] ),
    .A2(_1263_),
    .B1(_1265_),
    .B2(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__o221a_1 _1655_ (.A1(\outputs.output_gen.count[3] ),
    .A2(_1259_),
    .B1(_1263_),
    .B2(\outputs.output_gen.count[2] ),
    .C1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__o31a_1 _1656_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(\outputs.scaled_buffer[1] ),
    .A3(\outputs.scaled_buffer[2] ),
    .B1(net21),
    .X(_1270_));
 sky130_fd_sc_hd__xor2_1 _1657_ (.A(\outputs.scaled_buffer[3] ),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a221oi_2 _1658_ (.A1(\outputs.scaled_buffer[4] ),
    .A2(_1250_),
    .B1(_1271_),
    .B2(_1246_),
    .C1(_1254_),
    .Y(_1272_));
 sky130_fd_sc_hd__a22o_1 _1659_ (.A1(\outputs.output_gen.count[4] ),
    .A2(_1272_),
    .B1(_1259_),
    .B2(\outputs.output_gen.count[3] ),
    .X(_1273_));
 sky130_fd_sc_hd__or2_1 _1660_ (.A(\outputs.output_gen.count[4] ),
    .B(_1272_),
    .X(_1274_));
 sky130_fd_sc_hd__o221a_1 _1661_ (.A1(\outputs.output_gen.count[5] ),
    .A2(_1256_),
    .B1(_1269_),
    .B2(_1273_),
    .C1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__o21ai_1 _1662_ (.A1(\outputs.scaled_buffer[4] ),
    .A2(_1188_),
    .B1(net21),
    .Y(_1276_));
 sky130_fd_sc_hd__xnor2_1 _1663_ (.A(\outputs.scaled_buffer[5] ),
    .B(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__a221oi_2 _1664_ (.A1(\outputs.scaled_buffer[6] ),
    .A2(_1250_),
    .B1(_1277_),
    .B2(_1246_),
    .C1(_1254_),
    .Y(_1278_));
 sky130_fd_sc_hd__a22o_1 _1665_ (.A1(\outputs.output_gen.count[5] ),
    .A2(_1256_),
    .B1(_1278_),
    .B2(\outputs.output_gen.count[6] ),
    .X(_1279_));
 sky130_fd_sc_hd__a21oi_1 _1666_ (.A1(net21),
    .A2(_1252_),
    .B1(\outputs.scaled_buffer[6] ),
    .Y(_1280_));
 sky130_fd_sc_hd__a31o_1 _1667_ (.A1(\outputs.scaled_buffer[6] ),
    .A2(net21),
    .A3(_1252_),
    .B1(_1247_),
    .X(_1281_));
 sky130_fd_sc_hd__a21oi_1 _1668_ (.A1(\outputs.scaled_buffer[7] ),
    .A2(_1250_),
    .B1(_1254_),
    .Y(_1282_));
 sky130_fd_sc_hd__o21a_1 _1669_ (.A1(_1280_),
    .A2(_1281_),
    .B1(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__or2_1 _1670_ (.A(\outputs.output_gen.count[6] ),
    .B(_1278_),
    .X(_1284_));
 sky130_fd_sc_hd__o221a_1 _1671_ (.A1(_1275_),
    .A2(_1279_),
    .B1(_1283_),
    .B2(\outputs.output_gen.count[7] ),
    .C1(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__nand2_1 _1672_ (.A(\outputs.output_gen.count[7] ),
    .B(_1283_),
    .Y(_1286_));
 sky130_fd_sc_hd__nor3_2 _1673_ (.A(\inputs.key_encoder.sync_keys[14] ),
    .B(\inputs.key_encoder.sync_keys[15] ),
    .C(\inputs.key_encoder.octave_key_up ),
    .Y(_1287_));
 sky130_fd_sc_hd__or4_4 _1674_ (.A(\inputs.key_encoder.sync_keys[11] ),
    .B(\inputs.key_encoder.sync_keys[8] ),
    .C(\inputs.key_encoder.sync_keys[9] ),
    .D(\inputs.key_encoder.sync_keys[10] ),
    .X(_1288_));
 sky130_fd_sc_hd__or2_1 _1675_ (.A(\inputs.key_encoder.sync_keys[2] ),
    .B(\inputs.key_encoder.sync_keys[3] ),
    .X(_1289_));
 sky130_fd_sc_hd__or4_1 _1676_ (.A(\inputs.key_encoder.sync_keys[13] ),
    .B(\inputs.key_encoder.sync_keys[1] ),
    .C(\inputs.key_encoder.sync_keys[0] ),
    .D(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__or4_1 _1677_ (.A(\inputs.key_encoder.sync_keys[4] ),
    .B(\inputs.key_encoder.sync_keys[5] ),
    .C(\inputs.key_encoder.sync_keys[6] ),
    .D(\inputs.key_encoder.sync_keys[7] ),
    .X(_1291_));
 sky130_fd_sc_hd__or4_1 _1678_ (.A(\inputs.key_encoder.sync_keys[12] ),
    .B(_1288_),
    .C(_1290_),
    .D(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__and4b_1 _1679_ (.A_N(_1285_),
    .B(_1286_),
    .C(_1287_),
    .D(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _1680_ (.A(_1293_),
    .X(\outputs.output_gen.pwm_unff ));
 sky130_fd_sc_hd__buf_4 _1681_ (.A(_1081_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _1682_ (.A0(\outputs.div.m[0] ),
    .A1(net297),
    .S(_1294_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _1683_ (.A(_0209_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(\outputs.div.m[1] ),
    .A1(\outputs.div.divisor[1] ),
    .S(_1294_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _1685_ (.A(_0210_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(\outputs.div.m[2] ),
    .A1(net315),
    .S(_1294_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _1687_ (.A(_0211_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _1688_ (.A0(\outputs.div.m[3] ),
    .A1(net292),
    .S(_1294_),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _1689_ (.A(_0212_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _1690_ (.A0(\outputs.div.m[4] ),
    .A1(\outputs.div.divisor[4] ),
    .S(_1294_),
    .X(_0213_));
 sky130_fd_sc_hd__clkbuf_1 _1691_ (.A(_0213_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _1692_ (.A0(\outputs.div.m[5] ),
    .A1(\outputs.div.divisor[5] ),
    .S(_1294_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _1693_ (.A(_0214_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _1694_ (.A0(\outputs.div.m[6] ),
    .A1(net316),
    .S(_1294_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_1 _1695_ (.A(_0215_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(\outputs.div.m[7] ),
    .A1(\outputs.div.divisor[7] ),
    .S(_1294_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _1697_ (.A(_0216_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _1698_ (.A0(\outputs.div.m[8] ),
    .A1(net308),
    .S(_1294_),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_1 _1699_ (.A(_0217_),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_4 _1700_ (.A(_1089_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1701_ (.A0(\outputs.div.m[9] ),
    .A1(net217),
    .S(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_1 _1702_ (.A(_0219_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(\outputs.div.m[10] ),
    .A1(\outputs.div.divisor[10] ),
    .S(_0218_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _1704_ (.A(_0220_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(\outputs.div.m[11] ),
    .A1(net278),
    .S(_0218_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_1 _1706_ (.A(_0221_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _1707_ (.A0(\outputs.div.m[12] ),
    .A1(net276),
    .S(_0218_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _1708_ (.A(_0222_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _1709_ (.A0(\outputs.div.m[13] ),
    .A1(\outputs.div.divisor[13] ),
    .S(_0218_),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_1 _1710_ (.A(_0223_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _1711_ (.A0(\outputs.div.m[14] ),
    .A1(net269),
    .S(_0218_),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_1 _1712_ (.A(_0224_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _1713_ (.A0(\outputs.div.m[15] ),
    .A1(net313),
    .S(_0218_),
    .X(_0225_));
 sky130_fd_sc_hd__clkbuf_1 _1714_ (.A(_0225_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _1715_ (.A0(\outputs.div.m[16] ),
    .A1(net298),
    .S(_0218_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _1716_ (.A(_0226_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _1717_ (.A0(\outputs.div.m[17] ),
    .A1(\outputs.div.divisor[17] ),
    .S(_0218_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_1 _1718_ (.A(_0227_),
    .X(_0017_));
 sky130_fd_sc_hd__nor2_1 _1719_ (.A(\inputs.octave_fsm.state[1] ),
    .B(\inputs.octave_fsm.state[0] ),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_1 _1720_ (.A(\inputs.octave_fsm.state[2] ),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__clkbuf_4 _1721_ (.A(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__clkbuf_4 _1722_ (.A(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__or2b_1 _1723_ (.A(\inputs.octave_fsm.state[2] ),
    .B_N(\inputs.octave_fsm.state[1] ),
    .X(_0232_));
 sky130_fd_sc_hd__and2b_1 _1724_ (.A_N(\inputs.down.det_edge ),
    .B(\inputs.octave_fsm.octave_key_up ),
    .X(_0233_));
 sky130_fd_sc_hd__or2b_1 _1725_ (.A(\inputs.octave_fsm.octave_key_up ),
    .B_N(\inputs.down.det_edge ),
    .X(_0234_));
 sky130_fd_sc_hd__or2b_1 _1726_ (.A(_0233_),
    .B_N(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__a21oi_1 _1727_ (.A1(_0231_),
    .A2(_0232_),
    .B1(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2b_2 _1728_ (.A(\inputs.octave_fsm.state[2] ),
    .B_N(\inputs.octave_fsm.state[0] ),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _1729_ (.A(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__nor2_1 _1730_ (.A(\inputs.octave_fsm.state[1] ),
    .B(_0233_),
    .Y(_0239_));
 sky130_fd_sc_hd__o32a_1 _1731_ (.A1(\inputs.octave_fsm.state[0] ),
    .A2(\inputs.octave_fsm.state[2] ),
    .A3(_0239_),
    .B1(_0231_),
    .B2(_0233_),
    .X(_0240_));
 sky130_fd_sc_hd__o31a_1 _1732_ (.A1(\inputs.octave_fsm.state[1] ),
    .A2(_0235_),
    .A3(_0238_),
    .B1(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__xnor2_1 _1733_ (.A(_0236_),
    .B(_0241_),
    .Y(_0018_));
 sky130_fd_sc_hd__a21o_1 _1734_ (.A1(\inputs.octave_fsm.state[1] ),
    .A2(\inputs.octave_fsm.state[0] ),
    .B1(\inputs.octave_fsm.state[2] ),
    .X(_0242_));
 sky130_fd_sc_hd__and3b_1 _1735_ (.A_N(\inputs.octave_fsm.state[2] ),
    .B(\inputs.octave_fsm.state[0] ),
    .C(\inputs.octave_fsm.state[1] ),
    .X(_0243_));
 sky130_fd_sc_hd__nor2_1 _1736_ (.A(_0228_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__mux2_1 _1737_ (.A0(_0242_),
    .A1(_0244_),
    .S(_0233_),
    .X(_0245_));
 sky130_fd_sc_hd__o22a_1 _1738_ (.A1(_0235_),
    .A2(_0231_),
    .B1(_0236_),
    .B2(_0245_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _1739_ (.A(\inputs.octave_fsm.state[2] ),
    .B(_0228_),
    .X(_0246_));
 sky130_fd_sc_hd__buf_2 _1740_ (.A(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__a22o_1 _1741_ (.A1(_0234_),
    .A2(_0247_),
    .B1(_0243_),
    .B2(_0233_),
    .X(_0020_));
 sky130_fd_sc_hd__buf_2 _1742_ (.A(_1082_),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_4 _1743_ (.A(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _1744_ (.A(\outputs.div.m[0] ),
    .B(\outputs.div.q[26] ),
    .Y(_0250_));
 sky130_fd_sc_hd__or2_1 _1745_ (.A(\outputs.div.m[0] ),
    .B(\outputs.div.q[26] ),
    .X(_0251_));
 sky130_fd_sc_hd__buf_4 _1746_ (.A(_1003_),
    .X(_0252_));
 sky130_fd_sc_hd__a32o_1 _1747_ (.A1(_0249_),
    .A2(_0250_),
    .A3(_0251_),
    .B1(_0252_),
    .B2(net140),
    .X(_0021_));
 sky130_fd_sc_hd__inv_2 _1748_ (.A(\outputs.div.a[25] ),
    .Y(_0253_));
 sky130_fd_sc_hd__a21o_1 _1749_ (.A1(\outputs.div.m[0] ),
    .A2(_0253_),
    .B1(\outputs.div.m[1] ),
    .X(_0254_));
 sky130_fd_sc_hd__nand3_1 _1750_ (.A(\outputs.div.m[0] ),
    .B(\outputs.div.m[1] ),
    .C(_0253_),
    .Y(_0255_));
 sky130_fd_sc_hd__and3_1 _1751_ (.A(\outputs.div.a[0] ),
    .B(_0254_),
    .C(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__a21oi_1 _1752_ (.A1(_0254_),
    .A2(_0255_),
    .B1(\outputs.div.a[0] ),
    .Y(_0257_));
 sky130_fd_sc_hd__or2_1 _1753_ (.A(_0256_),
    .B(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__xor2_1 _1754_ (.A(_0250_),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__a22o_1 _1755_ (.A1(net181),
    .A2(_1004_),
    .B1(\outputs.div.next_div ),
    .B2(_0259_),
    .X(_0022_));
 sky130_fd_sc_hd__o21ba_1 _1756_ (.A1(_0250_),
    .A2(_0257_),
    .B1_N(_0256_),
    .X(_0260_));
 sky130_fd_sc_hd__inv_2 _1757_ (.A(\outputs.div.a[1] ),
    .Y(_0261_));
 sky130_fd_sc_hd__o21ba_1 _1758_ (.A1(\outputs.div.m[0] ),
    .A2(\outputs.div.m[1] ),
    .B1_N(\outputs.div.a[25] ),
    .X(_0262_));
 sky130_fd_sc_hd__xnor2_1 _1759_ (.A(\outputs.div.m[2] ),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__or2_1 _1760_ (.A(_0261_),
    .B(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_1 _1761_ (.A(_0261_),
    .B(_0263_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _1762_ (.A(_0264_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__or2_1 _1763_ (.A(_0260_),
    .B(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _1764_ (.A(_0260_),
    .B(_0266_),
    .Y(_0268_));
 sky130_fd_sc_hd__a32o_1 _1765_ (.A1(_0249_),
    .A2(_0267_),
    .A3(_0268_),
    .B1(_0252_),
    .B2(net203),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_1 _1766_ (.A(_0264_),
    .B(_0267_),
    .Y(_0269_));
 sky130_fd_sc_hd__a21o_1 _1767_ (.A1(\outputs.div.m[2] ),
    .A2(_0253_),
    .B1(_0262_),
    .X(_0270_));
 sky130_fd_sc_hd__xor2_1 _1768_ (.A(\outputs.div.m[3] ),
    .B(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__and2_1 _1769_ (.A(\outputs.div.a[2] ),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _1770_ (.A(\outputs.div.a[2] ),
    .B(_0271_),
    .Y(_0273_));
 sky130_fd_sc_hd__nor2_1 _1771_ (.A(_0272_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nand2_1 _1772_ (.A(_0269_),
    .B(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__o21a_1 _1773_ (.A1(_0269_),
    .A2(_0274_),
    .B1(_1084_),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _1774_ (.A1(net299),
    .A2(_1004_),
    .B1(_0275_),
    .B2(_0276_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_4 _1775_ (.A(_1084_),
    .X(_0277_));
 sky130_fd_sc_hd__nand2_1 _1776_ (.A(\outputs.div.a[2] ),
    .B(_0271_),
    .Y(_0278_));
 sky130_fd_sc_hd__o211a_1 _1777_ (.A1(_0260_),
    .A2(_0266_),
    .B1(_0278_),
    .C1(_0264_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_1 _1778_ (.A(_0273_),
    .B(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__or4_2 _1779_ (.A(\outputs.div.m[3] ),
    .B(\outputs.div.m[2] ),
    .C(\outputs.div.m[0] ),
    .D(\outputs.div.m[1] ),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _1780_ (.A(_0253_),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__xor2_2 _1781_ (.A(\outputs.div.m[4] ),
    .B(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__xnor2_1 _1782_ (.A(\outputs.div.a[3] ),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__or2_1 _1783_ (.A(_0280_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__nand2_1 _1784_ (.A(_0280_),
    .B(_0284_),
    .Y(_0286_));
 sky130_fd_sc_hd__a32o_1 _1785_ (.A1(_0277_),
    .A2(_0285_),
    .A3(_0286_),
    .B1(_0252_),
    .B2(net154),
    .X(_0025_));
 sky130_fd_sc_hd__inv_2 _1786_ (.A(\outputs.div.a[3] ),
    .Y(_0287_));
 sky130_fd_sc_hd__or2_1 _1787_ (.A(_0287_),
    .B(_0283_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _1788_ (.A(\outputs.div.a[4] ),
    .Y(_0289_));
 sky130_fd_sc_hd__o21a_1 _1789_ (.A1(\outputs.div.m[4] ),
    .A2(_0281_),
    .B1(_0253_),
    .X(_0290_));
 sky130_fd_sc_hd__xnor2_2 _1790_ (.A(\outputs.div.m[5] ),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__xnor2_1 _1791_ (.A(_0289_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__nand3_1 _1792_ (.A(_0288_),
    .B(_0286_),
    .C(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__a21o_1 _1793_ (.A1(_0288_),
    .A2(_0286_),
    .B1(_0292_),
    .X(_0294_));
 sky130_fd_sc_hd__a32o_1 _1794_ (.A1(_0277_),
    .A2(_0293_),
    .A3(_0294_),
    .B1(_0252_),
    .B2(net173),
    .X(_0026_));
 sky130_fd_sc_hd__inv_2 _1795_ (.A(\outputs.div.a[5] ),
    .Y(_0295_));
 sky130_fd_sc_hd__or2_1 _1796_ (.A(\outputs.div.m[5] ),
    .B(\outputs.div.m[4] ),
    .X(_0296_));
 sky130_fd_sc_hd__o21a_1 _1797_ (.A1(_0281_),
    .A2(_0296_),
    .B1(_0253_),
    .X(_0297_));
 sky130_fd_sc_hd__xnor2_1 _1798_ (.A(\outputs.div.m[6] ),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__or2_1 _1799_ (.A(_0295_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _1800_ (.A(_0295_),
    .B(_0298_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _1801_ (.A(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand2_1 _1802_ (.A(_0287_),
    .B(_0283_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _1803_ (.A(_0288_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__o22a_1 _1804_ (.A1(_0287_),
    .A2(_0283_),
    .B1(_0291_),
    .B2(_0289_),
    .X(_0304_));
 sky130_fd_sc_hd__a21o_1 _1805_ (.A1(_0289_),
    .A2(_0291_),
    .B1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__o41a_1 _1806_ (.A1(_0273_),
    .A2(_0279_),
    .A3(_0303_),
    .A4(_0292_),
    .B1(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _1807_ (.A(_0301_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__or2_1 _1808_ (.A(_0301_),
    .B(_0306_),
    .X(_0308_));
 sky130_fd_sc_hd__a32o_1 _1809_ (.A1(_0277_),
    .A2(_0307_),
    .A3(_0308_),
    .B1(_0252_),
    .B2(net169),
    .X(_0027_));
 sky130_fd_sc_hd__inv_2 _1810_ (.A(\outputs.div.a[6] ),
    .Y(_0309_));
 sky130_fd_sc_hd__o31a_1 _1811_ (.A1(\outputs.div.m[6] ),
    .A2(_0281_),
    .A3(_0296_),
    .B1(_0253_),
    .X(_0310_));
 sky130_fd_sc_hd__xnor2_1 _1812_ (.A(\outputs.div.m[7] ),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__nor2_1 _1813_ (.A(_0309_),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__and2_1 _1814_ (.A(_0309_),
    .B(_0311_),
    .X(_0313_));
 sky130_fd_sc_hd__or2_1 _1815_ (.A(_0312_),
    .B(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__o21a_1 _1816_ (.A1(_0301_),
    .A2(_0306_),
    .B1(_0299_),
    .X(_0315_));
 sky130_fd_sc_hd__xor2_1 _1817_ (.A(_0314_),
    .B(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _1818_ (.A1(net185),
    .A2(_1004_),
    .B1(\outputs.div.next_div ),
    .B2(_0316_),
    .X(_0028_));
 sky130_fd_sc_hd__o21a_1 _1819_ (.A1(_0309_),
    .A2(_0311_),
    .B1(_0299_),
    .X(_0317_));
 sky130_fd_sc_hd__o32a_2 _1820_ (.A1(_0301_),
    .A2(_0306_),
    .A3(_0314_),
    .B1(_0317_),
    .B2(_0313_),
    .X(_0318_));
 sky130_fd_sc_hd__inv_2 _1821_ (.A(\outputs.div.a[7] ),
    .Y(_0319_));
 sky130_fd_sc_hd__buf_2 _1822_ (.A(_0253_),
    .X(_0320_));
 sky130_fd_sc_hd__or4_2 _1823_ (.A(\outputs.div.m[7] ),
    .B(\outputs.div.m[6] ),
    .C(_0281_),
    .D(_0296_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2_1 _1824_ (.A(_0320_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__xor2_1 _1825_ (.A(\outputs.div.m[8] ),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_1 _1826_ (.A(_0319_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__and2_1 _1827_ (.A(_0319_),
    .B(_0323_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_2 _1828_ (.A(_0324_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_1 _1829_ (.A(_0318_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21bo_1 _1830_ (.A1(_0318_),
    .A2(_0326_),
    .B1_N(_1084_),
    .X(_0328_));
 sky130_fd_sc_hd__a2bb2o_1 _1831_ (.A1_N(_0327_),
    .A2_N(_0328_),
    .B1(net161),
    .B2(_1004_),
    .X(_0029_));
 sky130_fd_sc_hd__o21a_1 _1832_ (.A1(\outputs.div.m[8] ),
    .A2(_0321_),
    .B1(_0253_),
    .X(_0329_));
 sky130_fd_sc_hd__xor2_1 _1833_ (.A(\outputs.div.m[9] ),
    .B(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__and2_1 _1834_ (.A(\outputs.div.a[8] ),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__or2_1 _1835_ (.A(\outputs.div.a[8] ),
    .B(_0330_),
    .X(_0332_));
 sky130_fd_sc_hd__and2b_1 _1836_ (.A_N(_0331_),
    .B(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _1837_ (.A1(_0324_),
    .A2(_0327_),
    .B1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__o31a_1 _1838_ (.A1(_0324_),
    .A2(_0327_),
    .A3(_0333_),
    .B1(_1084_),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _1839_ (.A1(net288),
    .A2(_1004_),
    .B1(_0334_),
    .B2(_0335_),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _1840_ (.A(\outputs.div.m[9] ),
    .B(\outputs.div.m[8] ),
    .X(_0336_));
 sky130_fd_sc_hd__o21a_1 _1841_ (.A1(_0321_),
    .A2(_0336_),
    .B1(_0320_),
    .X(_0337_));
 sky130_fd_sc_hd__xnor2_2 _1842_ (.A(\outputs.div.m[10] ),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__xnor2_2 _1843_ (.A(\outputs.div.a[9] ),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _1844_ (.A(_0333_),
    .Y(_0340_));
 sky130_fd_sc_hd__o21ai_1 _1845_ (.A1(_0324_),
    .A2(_0331_),
    .B1(_0332_),
    .Y(_0341_));
 sky130_fd_sc_hd__o31ai_4 _1846_ (.A1(_0318_),
    .A2(_0326_),
    .A3(_0340_),
    .B1(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__or2_1 _1847_ (.A(_0339_),
    .B(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__nand2_1 _1848_ (.A(_0339_),
    .B(_0342_),
    .Y(_0344_));
 sky130_fd_sc_hd__a32o_1 _1849_ (.A1(_0277_),
    .A2(_0343_),
    .A3(_0344_),
    .B1(_0252_),
    .B2(net175),
    .X(_0031_));
 sky130_fd_sc_hd__o31a_1 _1850_ (.A1(\outputs.div.m[10] ),
    .A2(_0321_),
    .A3(_0336_),
    .B1(_0320_),
    .X(_0345_));
 sky130_fd_sc_hd__xnor2_1 _1851_ (.A(\outputs.div.m[11] ),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _1852_ (.A(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_2 _1853_ (.A(\outputs.div.a[10] ),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__nor2_1 _1854_ (.A(\outputs.div.a[10] ),
    .B(_0347_),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _1855_ (.A(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _1856_ (.A(_0348_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _1857_ (.A(\outputs.div.a[9] ),
    .Y(_0352_));
 sky130_fd_sc_hd__or2_1 _1858_ (.A(_0352_),
    .B(_0338_),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_1 _1859_ (.A(_0353_),
    .B(_0344_),
    .Y(_0354_));
 sky130_fd_sc_hd__xnor2_1 _1860_ (.A(_0351_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__a22o_1 _1861_ (.A1(net179),
    .A2(_1004_),
    .B1(\outputs.div.next_div ),
    .B2(_0355_),
    .X(_0032_));
 sky130_fd_sc_hd__inv_2 _1862_ (.A(\outputs.div.a[11] ),
    .Y(_0356_));
 sky130_fd_sc_hd__or4_2 _1863_ (.A(\outputs.div.m[11] ),
    .B(\outputs.div.m[10] ),
    .C(_0321_),
    .D(_0336_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_1 _1864_ (.A(_0320_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__xor2_1 _1865_ (.A(\outputs.div.m[12] ),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _1866_ (.A(_0356_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__nand2_1 _1867_ (.A(_0356_),
    .B(_0359_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _1868_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__a21oi_1 _1869_ (.A1(_0353_),
    .A2(_0348_),
    .B1(_0349_),
    .Y(_0363_));
 sky130_fd_sc_hd__a41oi_4 _1870_ (.A1(_0339_),
    .A2(_0342_),
    .A3(_0348_),
    .A4(_0350_),
    .B1(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2_1 _1871_ (.A(_0362_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__or2_1 _1872_ (.A(_0362_),
    .B(_0364_),
    .X(_0366_));
 sky130_fd_sc_hd__a32o_1 _1873_ (.A1(_0277_),
    .A2(_0365_),
    .A3(_0366_),
    .B1(_0252_),
    .B2(net165),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _1874_ (.A(\outputs.div.a[12] ),
    .Y(_0367_));
 sky130_fd_sc_hd__o21a_1 _1875_ (.A1(\outputs.div.m[12] ),
    .A2(_0357_),
    .B1(_0320_),
    .X(_0368_));
 sky130_fd_sc_hd__xnor2_1 _1876_ (.A(\outputs.div.m[13] ),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _1877_ (.A(_0367_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__and2_1 _1878_ (.A(_0367_),
    .B(_0369_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _1879_ (.A(_0370_),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__o21ai_1 _1880_ (.A1(_0362_),
    .A2(_0364_),
    .B1(_0360_),
    .Y(_0373_));
 sky130_fd_sc_hd__xnor2_1 _1881_ (.A(_0372_),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__a22o_1 _1882_ (.A1(net182),
    .A2(_1004_),
    .B1(\outputs.div.next_div ),
    .B2(_0374_),
    .X(_0034_));
 sky130_fd_sc_hd__inv_2 _1883_ (.A(\outputs.div.a[13] ),
    .Y(_0375_));
 sky130_fd_sc_hd__o31a_1 _1884_ (.A1(\outputs.div.m[13] ),
    .A2(\outputs.div.m[12] ),
    .A3(_0357_),
    .B1(_0320_),
    .X(_0376_));
 sky130_fd_sc_hd__xnor2_1 _1885_ (.A(\outputs.div.m[14] ),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__or2_1 _1886_ (.A(_0375_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _1887_ (.A(_0375_),
    .B(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _1888_ (.A(_0378_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _1889_ (.A(_0370_),
    .Y(_0381_));
 sky130_fd_sc_hd__a21o_1 _1890_ (.A1(_0360_),
    .A2(_0381_),
    .B1(_0371_),
    .X(_0382_));
 sky130_fd_sc_hd__o31a_1 _1891_ (.A1(_0362_),
    .A2(_0364_),
    .A3(_0372_),
    .B1(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _1892_ (.A(_0380_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__or2_1 _1893_ (.A(_0380_),
    .B(_0383_),
    .X(_0385_));
 sky130_fd_sc_hd__a32o_1 _1894_ (.A1(_0277_),
    .A2(_0384_),
    .A3(_0385_),
    .B1(_0252_),
    .B2(net126),
    .X(_0035_));
 sky130_fd_sc_hd__or4_1 _1895_ (.A(\outputs.div.m[14] ),
    .B(\outputs.div.m[13] ),
    .C(\outputs.div.m[12] ),
    .D(_0357_),
    .X(_0386_));
 sky130_fd_sc_hd__nand2_1 _1896_ (.A(_0320_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__xor2_1 _1897_ (.A(\outputs.div.m[15] ),
    .B(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__inv_2 _1898_ (.A(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_1 _1899_ (.A(\outputs.div.a[14] ),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__or2_1 _1900_ (.A(\outputs.div.a[14] ),
    .B(_0389_),
    .X(_0391_));
 sky130_fd_sc_hd__nand2_1 _1901_ (.A(_0390_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__o21ai_1 _1902_ (.A1(_0380_),
    .A2(_0383_),
    .B1(_0378_),
    .Y(_0393_));
 sky130_fd_sc_hd__xnor2_1 _1903_ (.A(_0392_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__a22o_1 _1904_ (.A1(net192),
    .A2(_1004_),
    .B1(\outputs.div.next_div ),
    .B2(_0394_),
    .X(_0036_));
 sky130_fd_sc_hd__inv_2 _1905_ (.A(\outputs.div.a[15] ),
    .Y(_0395_));
 sky130_fd_sc_hd__o21a_1 _1906_ (.A1(\outputs.div.m[15] ),
    .A2(_0386_),
    .B1(_0320_),
    .X(_0396_));
 sky130_fd_sc_hd__xnor2_1 _1907_ (.A(\outputs.div.m[16] ),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__or2_1 _1908_ (.A(_0395_),
    .B(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _1909_ (.A(_0395_),
    .B(_0397_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _1910_ (.A(_0398_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__a21bo_1 _1911_ (.A1(_0378_),
    .A2(_0390_),
    .B1_N(_0391_),
    .X(_0401_));
 sky130_fd_sc_hd__o31a_2 _1912_ (.A1(_0380_),
    .A2(_0383_),
    .A3(_0392_),
    .B1(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _1913_ (.A(_0400_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__or2_1 _1914_ (.A(_0400_),
    .B(_0402_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_4 _1915_ (.A(_1002_),
    .X(_0405_));
 sky130_fd_sc_hd__a32o_1 _1916_ (.A1(_0277_),
    .A2(_0403_),
    .A3(_0404_),
    .B1(_0405_),
    .B2(net158),
    .X(_0037_));
 sky130_fd_sc_hd__inv_2 _1917_ (.A(\outputs.div.a[16] ),
    .Y(_0406_));
 sky130_fd_sc_hd__or3_1 _1918_ (.A(\outputs.div.m[16] ),
    .B(\outputs.div.m[15] ),
    .C(_0386_),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _1919_ (.A(_0320_),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__xnor2_2 _1920_ (.A(\outputs.div.m[17] ),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__xnor2_1 _1921_ (.A(_0406_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__o21ai_1 _1922_ (.A1(_0400_),
    .A2(_0402_),
    .B1(_0398_),
    .Y(_0411_));
 sky130_fd_sc_hd__xnor2_1 _1923_ (.A(_0410_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__a22o_1 _1924_ (.A1(net260),
    .A2(_1004_),
    .B1(\outputs.div.next_div ),
    .B2(_0412_),
    .X(_0038_));
 sky130_fd_sc_hd__clkbuf_4 _1925_ (.A(_1003_),
    .X(_0413_));
 sky130_fd_sc_hd__o21a_2 _1926_ (.A1(\outputs.div.m[17] ),
    .A2(_0407_),
    .B1(_0320_),
    .X(_0414_));
 sky130_fd_sc_hd__nand2_1 _1927_ (.A(\outputs.div.a[17] ),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__or2_1 _1928_ (.A(\outputs.div.a[17] ),
    .B(_0414_),
    .X(_0416_));
 sky130_fd_sc_hd__nand2_1 _1929_ (.A(_0415_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__or2_1 _1930_ (.A(_0400_),
    .B(_0410_),
    .X(_0418_));
 sky130_fd_sc_hd__o21a_1 _1931_ (.A1(_0406_),
    .A2(_0409_),
    .B1(_0398_),
    .X(_0419_));
 sky130_fd_sc_hd__a21oi_1 _1932_ (.A1(_0406_),
    .A2(_0409_),
    .B1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__o21ba_1 _1933_ (.A1(_0402_),
    .A2(_0418_),
    .B1_N(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__xor2_1 _1934_ (.A(_0417_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_1 _1935_ (.A1(net256),
    .A2(_0413_),
    .B1(\outputs.div.next_div ),
    .B2(_0422_),
    .X(_0039_));
 sky130_fd_sc_hd__xnor2_2 _1936_ (.A(\outputs.div.a[18] ),
    .B(_0414_),
    .Y(_0423_));
 sky130_fd_sc_hd__o21ai_1 _1937_ (.A1(_0417_),
    .A2(_0421_),
    .B1(_0415_),
    .Y(_0424_));
 sky130_fd_sc_hd__xnor2_1 _1938_ (.A(_0423_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a22o_1 _1939_ (.A1(net295),
    .A2(_0413_),
    .B1(\outputs.div.next_div ),
    .B2(_0425_),
    .X(_0040_));
 sky130_fd_sc_hd__or3_1 _1940_ (.A(_0417_),
    .B(_0418_),
    .C(_0423_),
    .X(_0426_));
 sky130_fd_sc_hd__buf_2 _1941_ (.A(_0414_),
    .X(_0427_));
 sky130_fd_sc_hd__o21ai_1 _1942_ (.A1(\outputs.div.a[18] ),
    .A2(\outputs.div.a[17] ),
    .B1(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__a2111o_1 _1943_ (.A1(_0406_),
    .A2(_0409_),
    .B1(_0417_),
    .C1(_0419_),
    .D1(_0423_),
    .X(_0429_));
 sky130_fd_sc_hd__o211a_1 _1944_ (.A1(_0402_),
    .A2(_0426_),
    .B1(_0428_),
    .C1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _1945_ (.A(\outputs.div.a[19] ),
    .B(_0414_),
    .Y(_0431_));
 sky130_fd_sc_hd__or2_1 _1946_ (.A(\outputs.div.a[19] ),
    .B(_0414_),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_1 _1947_ (.A(_0431_),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2_1 _1948_ (.A(_0430_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__or2_1 _1949_ (.A(_0430_),
    .B(_0433_),
    .X(_0435_));
 sky130_fd_sc_hd__a32o_1 _1950_ (.A1(_0277_),
    .A2(_0434_),
    .A3(_0435_),
    .B1(_0405_),
    .B2(net281),
    .X(_0041_));
 sky130_fd_sc_hd__xnor2_1 _1951_ (.A(\outputs.div.a[20] ),
    .B(_0427_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand3_1 _1952_ (.A(_0431_),
    .B(_0435_),
    .C(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21o_1 _1953_ (.A1(_0431_),
    .A2(_0435_),
    .B1(_0436_),
    .X(_0438_));
 sky130_fd_sc_hd__a32o_1 _1954_ (.A1(_0277_),
    .A2(_0437_),
    .A3(_0438_),
    .B1(_0405_),
    .B2(net222),
    .X(_0042_));
 sky130_fd_sc_hd__o21ai_1 _1955_ (.A1(\outputs.div.a[20] ),
    .A2(\outputs.div.a[19] ),
    .B1(_0427_),
    .Y(_0439_));
 sky130_fd_sc_hd__o211ai_1 _1956_ (.A1(_0402_),
    .A2(_0426_),
    .B1(_0428_),
    .C1(_0429_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _1957_ (.A(_0433_),
    .B(_0436_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_1 _1958_ (.A(_0440_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _1959_ (.A(\outputs.div.a[21] ),
    .B(_0427_),
    .Y(_0443_));
 sky130_fd_sc_hd__or2_1 _1960_ (.A(\outputs.div.a[21] ),
    .B(_0414_),
    .X(_0444_));
 sky130_fd_sc_hd__nand2_1 _1961_ (.A(_0443_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__a21o_1 _1962_ (.A1(_0439_),
    .A2(_0442_),
    .B1(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__a311oi_1 _1963_ (.A1(_0445_),
    .A2(_0439_),
    .A3(_0442_),
    .B1(_1001_),
    .C1(_1294_),
    .Y(_0447_));
 sky130_fd_sc_hd__a22o_1 _1964_ (.A1(net283),
    .A2(_0413_),
    .B1(_0446_),
    .B2(_0447_),
    .X(_0043_));
 sky130_fd_sc_hd__xnor2_1 _1965_ (.A(\outputs.div.a[22] ),
    .B(_0427_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand3_1 _1966_ (.A(_0443_),
    .B(_0446_),
    .C(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__a21o_1 _1967_ (.A1(_0443_),
    .A2(_0446_),
    .B1(_0448_),
    .X(_0450_));
 sky130_fd_sc_hd__a32o_1 _1968_ (.A1(_0277_),
    .A2(_0449_),
    .A3(_0450_),
    .B1(_0405_),
    .B2(net170),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_1 _1969_ (.A(_0445_),
    .B(_0448_),
    .Y(_0451_));
 sky130_fd_sc_hd__o41a_1 _1970_ (.A1(\outputs.div.a[22] ),
    .A2(\outputs.div.a[21] ),
    .A3(\outputs.div.a[20] ),
    .A4(\outputs.div.a[19] ),
    .B1(_0427_),
    .X(_0452_));
 sky130_fd_sc_hd__a31o_1 _1971_ (.A1(_0440_),
    .A2(_0441_),
    .A3(_0451_),
    .B1(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__nand2_1 _1972_ (.A(\outputs.div.a[23] ),
    .B(_0427_),
    .Y(_0454_));
 sky130_fd_sc_hd__or2_1 _1973_ (.A(\outputs.div.a[23] ),
    .B(_0427_),
    .X(_0455_));
 sky130_fd_sc_hd__and2_1 _1974_ (.A(_0454_),
    .B(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__nand2_1 _1975_ (.A(_0453_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__or2_1 _1976_ (.A(_0453_),
    .B(_0456_),
    .X(_0458_));
 sky130_fd_sc_hd__a32o_1 _1977_ (.A1(_1084_),
    .A2(_0457_),
    .A3(_0458_),
    .B1(_0405_),
    .B2(net133),
    .X(_0045_));
 sky130_fd_sc_hd__nand2_1 _1978_ (.A(\outputs.div.a[24] ),
    .B(_0427_),
    .Y(_0459_));
 sky130_fd_sc_hd__or2_1 _1979_ (.A(\outputs.div.a[24] ),
    .B(_0427_),
    .X(_0460_));
 sky130_fd_sc_hd__nand2_1 _1980_ (.A(_0459_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand3_1 _1981_ (.A(_0454_),
    .B(_0457_),
    .C(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21o_1 _1982_ (.A1(_0454_),
    .A2(_0457_),
    .B1(_0461_),
    .X(_0463_));
 sky130_fd_sc_hd__a32o_1 _1983_ (.A1(_1084_),
    .A2(_0462_),
    .A3(_0463_),
    .B1(_0405_),
    .B2(net274),
    .X(_0046_));
 sky130_fd_sc_hd__o311a_1 _1984_ (.A1(\outputs.div.m[17] ),
    .A2(\outputs.div.a[25] ),
    .A3(_0407_),
    .B1(_0454_),
    .C1(_0459_),
    .X(_0464_));
 sky130_fd_sc_hd__o21ai_1 _1985_ (.A1(_0457_),
    .A2(_0461_),
    .B1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a22o_1 _1986_ (.A1(net261),
    .A2(_0413_),
    .B1(\outputs.div.next_div ),
    .B2(_0465_),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_1 _1987_ (.A1(net213),
    .A2(_0413_),
    .B1(_0249_),
    .B2(net261),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _1988_ (.A1(\outputs.div.q[2] ),
    .A2(_0413_),
    .B1(_0249_),
    .B2(net213),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _1989_ (.A1(net210),
    .A2(_0413_),
    .B1(_0249_),
    .B2(net250),
    .X(_0050_));
 sky130_fd_sc_hd__a22o_1 _1990_ (.A1(net122),
    .A2(_0413_),
    .B1(_0249_),
    .B2(net210),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_1 _1991_ (.A1(net197),
    .A2(_0413_),
    .B1(_0249_),
    .B2(net122),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _1992_ (.A1(net199),
    .A2(_0413_),
    .B1(_0249_),
    .B2(net197),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_1 _1993_ (.A1(\outputs.div.q[7] ),
    .A2(_0252_),
    .B1(_0249_),
    .B2(net199),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _1994_ (.A(\outputs.div.q[7] ),
    .B(_0248_),
    .X(_0466_));
 sky130_fd_sc_hd__a221o_1 _1995_ (.A1(net155),
    .A2(_1090_),
    .B1(_0405_),
    .B2(\outputs.div.q[8] ),
    .C1(_0466_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _1996_ (.A(\outputs.div.q[8] ),
    .B(_0248_),
    .X(_0467_));
 sky130_fd_sc_hd__a221o_1 _1997_ (.A1(\outputs.div.oscillator_out[1] ),
    .A2(_1090_),
    .B1(_0405_),
    .B2(net136),
    .C1(_0467_),
    .X(_0056_));
 sky130_fd_sc_hd__clkbuf_4 _1998_ (.A(_1002_),
    .X(_0468_));
 sky130_fd_sc_hd__and2_1 _1999_ (.A(\outputs.div.q[9] ),
    .B(_0248_),
    .X(_0469_));
 sky130_fd_sc_hd__a221o_1 _2000_ (.A1(\outputs.div.oscillator_out[2] ),
    .A2(_1090_),
    .B1(_0468_),
    .B2(net120),
    .C1(_0469_),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _2001_ (.A(\outputs.div.q[10] ),
    .B(_0248_),
    .X(_0470_));
 sky130_fd_sc_hd__a221o_1 _2002_ (.A1(net92),
    .A2(_1090_),
    .B1(_0468_),
    .B2(\outputs.div.q[11] ),
    .C1(_0470_),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _2003_ (.A(\outputs.div.q[11] ),
    .B(_0248_),
    .X(_0471_));
 sky130_fd_sc_hd__a221o_1 _2004_ (.A1(net98),
    .A2(_1090_),
    .B1(_0468_),
    .B2(\outputs.div.q[12] ),
    .C1(_0471_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _2005_ (.A(\outputs.div.q[12] ),
    .B(_0248_),
    .X(_0472_));
 sky130_fd_sc_hd__a221o_1 _2006_ (.A1(net150),
    .A2(_1090_),
    .B1(_0468_),
    .B2(\outputs.div.q[13] ),
    .C1(_0472_),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _2007_ (.A(\outputs.div.q[13] ),
    .B(_0248_),
    .X(_0473_));
 sky130_fd_sc_hd__a221o_1 _2008_ (.A1(net107),
    .A2(_1090_),
    .B1(_0468_),
    .B2(\outputs.div.q[14] ),
    .C1(_0473_),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _2009_ (.A(\outputs.div.q[14] ),
    .B(_0248_),
    .X(_0474_));
 sky130_fd_sc_hd__a221o_1 _2010_ (.A1(\outputs.div.oscillator_out[7] ),
    .A2(_1090_),
    .B1(_0468_),
    .B2(net116),
    .C1(_0474_),
    .X(_0062_));
 sky130_fd_sc_hd__clkbuf_4 _2011_ (.A(_1089_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _2012_ (.A(net116),
    .B(_0248_),
    .X(_0476_));
 sky130_fd_sc_hd__a221o_1 _2013_ (.A1(\outputs.div.oscillator_out[8] ),
    .A2(_0475_),
    .B1(_0468_),
    .B2(net124),
    .C1(_0476_),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _2014_ (.A(net124),
    .B(_1083_),
    .X(_0477_));
 sky130_fd_sc_hd__a221o_1 _2015_ (.A1(\outputs.div.oscillator_out[9] ),
    .A2(_0475_),
    .B1(_0468_),
    .B2(net134),
    .C1(_0477_),
    .X(_0064_));
 sky130_fd_sc_hd__and2_1 _2016_ (.A(net134),
    .B(_1083_),
    .X(_0478_));
 sky130_fd_sc_hd__a221o_1 _2017_ (.A1(\outputs.div.oscillator_out[10] ),
    .A2(_0475_),
    .B1(_0468_),
    .B2(net146),
    .C1(_0478_),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _2018_ (.A(\outputs.div.q[18] ),
    .B(_1083_),
    .X(_0479_));
 sky130_fd_sc_hd__a221o_1 _2019_ (.A1(\outputs.div.oscillator_out[11] ),
    .A2(_0475_),
    .B1(_0468_),
    .B2(net118),
    .C1(_0479_),
    .X(_0066_));
 sky130_fd_sc_hd__and2_1 _2020_ (.A(net118),
    .B(_1083_),
    .X(_0480_));
 sky130_fd_sc_hd__a221o_1 _2021_ (.A1(net127),
    .A2(_0475_),
    .B1(_1003_),
    .B2(\outputs.div.q[20] ),
    .C1(_0480_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _2022_ (.A(\outputs.div.q[20] ),
    .B(_1083_),
    .X(_0481_));
 sky130_fd_sc_hd__a221o_1 _2023_ (.A1(\outputs.div.oscillator_out[13] ),
    .A2(_0475_),
    .B1(_1003_),
    .B2(net152),
    .C1(_0481_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _2024_ (.A(\outputs.div.q[21] ),
    .B(_1083_),
    .X(_0482_));
 sky130_fd_sc_hd__a221o_1 _2025_ (.A1(net101),
    .A2(_0475_),
    .B1(_1003_),
    .B2(\outputs.div.q[22] ),
    .C1(_0482_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _2026_ (.A(\outputs.div.q[22] ),
    .B(_1083_),
    .X(_0483_));
 sky130_fd_sc_hd__a221o_1 _2027_ (.A1(net103),
    .A2(_0475_),
    .B1(_1003_),
    .B2(\outputs.div.q[23] ),
    .C1(_0483_),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _2028_ (.A(\outputs.div.q[23] ),
    .B(_1083_),
    .X(_0484_));
 sky130_fd_sc_hd__a221o_1 _2029_ (.A1(net109),
    .A2(_0475_),
    .B1(_1003_),
    .B2(\outputs.div.q[24] ),
    .C1(_0484_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _2030_ (.A(\outputs.div.q[24] ),
    .B(_1083_),
    .X(_0485_));
 sky130_fd_sc_hd__a221o_1 _2031_ (.A1(net159),
    .A2(_0475_),
    .B1(_1003_),
    .B2(\outputs.div.q[25] ),
    .C1(_0485_),
    .X(_0072_));
 sky130_fd_sc_hd__a22o_1 _2032_ (.A1(\outputs.div.q[26] ),
    .A2(_0252_),
    .B1(_0249_),
    .B2(net264),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2033_ (.A0(_1084_),
    .A1(_1003_),
    .S(\outputs.div.count[0] ),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _2034_ (.A(_0486_),
    .X(_0074_));
 sky130_fd_sc_hd__nand2_1 _2035_ (.A(\outputs.div.count[1] ),
    .B(\outputs.div.count[0] ),
    .Y(_0487_));
 sky130_fd_sc_hd__or2_1 _2036_ (.A(\outputs.div.count[1] ),
    .B(\outputs.div.count[0] ),
    .X(_0488_));
 sky130_fd_sc_hd__a32o_1 _2037_ (.A1(_0487_),
    .A2(_1084_),
    .A3(_0488_),
    .B1(_0405_),
    .B2(net263),
    .X(_0075_));
 sky130_fd_sc_hd__and3_1 _2038_ (.A(\outputs.div.count[2] ),
    .B(\outputs.div.count[1] ),
    .C(\outputs.div.count[0] ),
    .X(_0489_));
 sky130_fd_sc_hd__inv_2 _2039_ (.A(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__a32o_1 _2040_ (.A1(_0999_),
    .A2(_1084_),
    .A3(_0490_),
    .B1(_0405_),
    .B2(net162),
    .X(_0076_));
 sky130_fd_sc_hd__inv_2 _2041_ (.A(\outputs.div.count[3] ),
    .Y(_0491_));
 sky130_fd_sc_hd__or3_1 _2042_ (.A(_0491_),
    .B(_1001_),
    .C(_0490_),
    .X(_0492_));
 sky130_fd_sc_hd__a21o_1 _2043_ (.A1(\outputs.div.start ),
    .A2(_0489_),
    .B1(\outputs.div.count[3] ),
    .X(_0493_));
 sky130_fd_sc_hd__and3_1 _2044_ (.A(_0998_),
    .B(_0492_),
    .C(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _2045_ (.A(_0494_),
    .X(_0077_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(net211),
    .Y(_0495_));
 sky130_fd_sc_hd__a21oi_1 _2047_ (.A1(_0495_),
    .A2(_0492_),
    .B1(_1090_),
    .Y(_0078_));
 sky130_fd_sc_hd__mux2_1 _2048_ (.A0(\outputs.scaled_buffer[0] ),
    .A1(net129),
    .S(_0218_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _2049_ (.A(_0496_),
    .X(_0079_));
 sky130_fd_sc_hd__buf_4 _2050_ (.A(_1089_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _2051_ (.A0(\outputs.scaled_buffer[1] ),
    .A1(net105),
    .S(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _2052_ (.A(_0498_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2053_ (.A0(\outputs.scaled_buffer[2] ),
    .A1(net201),
    .S(_0497_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _2054_ (.A(_0499_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2055_ (.A0(\outputs.scaled_buffer[3] ),
    .A1(net163),
    .S(_0497_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _2056_ (.A(_0500_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2057_ (.A0(\outputs.scaled_buffer[4] ),
    .A1(net289),
    .S(_0497_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _2058_ (.A(_0501_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2059_ (.A0(\outputs.scaled_buffer[5] ),
    .A1(net143),
    .S(_0497_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _2060_ (.A(_0502_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2061_ (.A0(\outputs.scaled_buffer[6] ),
    .A1(net138),
    .S(_0497_),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _2062_ (.A(_0503_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2063_ (.A0(net303),
    .A1(net171),
    .S(_0497_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _2064_ (.A(_0504_),
    .X(_0086_));
 sky130_fd_sc_hd__and3_1 _2065_ (.A(\outputs.div.div ),
    .B(_0998_),
    .C(_1001_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_4 _2066_ (.A(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__or3b_1 _2067_ (.A(\outputs.div.q[7] ),
    .B(\outputs.div.q[6] ),
    .C_N(\outputs.div.q[8] ),
    .X(_0507_));
 sky130_fd_sc_hd__or4_1 _2068_ (.A(\outputs.div.q[3] ),
    .B(\outputs.div.q[2] ),
    .C(\outputs.div.q[5] ),
    .D(\outputs.div.q[4] ),
    .X(_0508_));
 sky130_fd_sc_hd__or4_1 _2069_ (.A(\outputs.div.q[1] ),
    .B(\outputs.div.q[0] ),
    .C(_0507_),
    .D(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_2 _2070_ (.A(_0506_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__o22a_1 _2071_ (.A1(net129),
    .A2(_0506_),
    .B1(_0510_),
    .B2(\outputs.div.q[0] ),
    .X(_0087_));
 sky130_fd_sc_hd__o22a_1 _2072_ (.A1(net105),
    .A2(_0506_),
    .B1(_0510_),
    .B2(\outputs.div.q[1] ),
    .X(_0088_));
 sky130_fd_sc_hd__o22a_1 _2073_ (.A1(net201),
    .A2(_0506_),
    .B1(_0510_),
    .B2(\outputs.div.q[2] ),
    .X(_0089_));
 sky130_fd_sc_hd__o22a_1 _2074_ (.A1(net163),
    .A2(_0506_),
    .B1(_0510_),
    .B2(\outputs.div.q[3] ),
    .X(_0090_));
 sky130_fd_sc_hd__o22a_1 _2075_ (.A1(\outputs.div.q_out[4] ),
    .A2(_0506_),
    .B1(_0510_),
    .B2(net122),
    .X(_0091_));
 sky130_fd_sc_hd__o22a_1 _2076_ (.A1(net143),
    .A2(_0506_),
    .B1(_0510_),
    .B2(\outputs.div.q[5] ),
    .X(_0092_));
 sky130_fd_sc_hd__o22a_1 _2077_ (.A1(net138),
    .A2(_0506_),
    .B1(_0510_),
    .B2(\outputs.div.q[6] ),
    .X(_0093_));
 sky130_fd_sc_hd__o22a_1 _2078_ (.A1(net171),
    .A2(_0506_),
    .B1(_0510_),
    .B2(\outputs.div.q[7] ),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _2079_ (.A(net43),
    .B(_1081_),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_4 _2080_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_4 _2081_ (.A(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _2082_ (.A0(net255),
    .A1(net317),
    .S(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _2083_ (.A(_0514_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _2084_ (.A0(net241),
    .A1(\outputs.div.divisor[1] ),
    .S(_0513_),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_1 _2085_ (.A(net242),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2086_ (.A0(\outputs.divider_buffer2[2] ),
    .A1(net279),
    .S(_0513_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _2087_ (.A(net280),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2088_ (.A0(net251),
    .A1(\outputs.div.divisor[3] ),
    .S(_0513_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _2089_ (.A(net252),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2090_ (.A0(net239),
    .A1(\outputs.div.divisor[4] ),
    .S(_0513_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _2091_ (.A(net240),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2092_ (.A0(net257),
    .A1(\outputs.div.divisor[5] ),
    .S(_0513_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_1 _2093_ (.A(net258),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(net224),
    .A1(net208),
    .S(_0513_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _2095_ (.A(_0520_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(net231),
    .A1(\outputs.div.divisor[7] ),
    .S(_0513_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _2097_ (.A(_0521_),
    .X(_0102_));
 sky130_fd_sc_hd__buf_4 _2098_ (.A(_0512_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _2099_ (.A0(net245),
    .A1(\outputs.div.divisor[8] ),
    .S(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_1 _2100_ (.A(_0523_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2101_ (.A0(net111),
    .A1(net253),
    .S(_0522_),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_1 _2102_ (.A(_0524_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2103_ (.A0(net275),
    .A1(\outputs.div.divisor[10] ),
    .S(_0522_),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _2104_ (.A(_0525_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2105_ (.A0(net246),
    .A1(\outputs.div.divisor[11] ),
    .S(_0522_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _2106_ (.A(net247),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(net226),
    .A1(net276),
    .S(_0522_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _2108_ (.A(_0527_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(net272),
    .A1(\outputs.div.divisor[13] ),
    .S(_0522_),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _2110_ (.A(_0528_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2111_ (.A0(\outputs.divider_buffer2[14] ),
    .A1(net269),
    .S(_0522_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _2112_ (.A(net270),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2113_ (.A0(net195),
    .A1(net220),
    .S(_0522_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _2114_ (.A(_0530_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(net266),
    .A1(\outputs.div.divisor[16] ),
    .S(_0522_),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _2116_ (.A(net267),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(net248),
    .A1(\outputs.div.divisor[17] ),
    .S(_0522_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _2118_ (.A(_0532_),
    .X(_0112_));
 sky130_fd_sc_hd__nand2_1 _2119_ (.A(\inputs.key_encoder.sync_keys[13] ),
    .B(_1287_),
    .Y(_0533_));
 sky130_fd_sc_hd__buf_2 _2120_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_4 _2121_ (.A(\inputs.frequency_lut.rng[2] ),
    .X(_0535_));
 sky130_fd_sc_hd__buf_2 _2122_ (.A(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_4 _2123_ (.A(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__inv_2 _2124_ (.A(\inputs.frequency_lut.rng[0] ),
    .Y(_0538_));
 sky130_fd_sc_hd__or2_1 _2125_ (.A(_0538_),
    .B(\inputs.frequency_lut.rng[1] ),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_4 _2126_ (.A(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__nand2_2 _2127_ (.A(_0538_),
    .B(\inputs.frequency_lut.rng[1] ),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_2 _2128_ (.A(_0540_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__buf_2 _2129_ (.A(\inputs.frequency_lut.rng[1] ),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _2130_ (.A(_0543_),
    .B(_0535_),
    .Y(_0544_));
 sky130_fd_sc_hd__o21a_1 _2131_ (.A1(_0537_),
    .A2(_0542_),
    .B1(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _2132_ (.A(_0538_),
    .B(\inputs.frequency_lut.rng[1] ),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_2 _2133_ (.A(_0535_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__and3_1 _2134_ (.A(\inputs.frequency_lut.rng[2] ),
    .B(_0539_),
    .C(_0541_),
    .X(_0548_));
 sky130_fd_sc_hd__buf_2 _2135_ (.A(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__nor2_1 _2136_ (.A(_0547_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__clkbuf_4 _2137_ (.A(\inputs.frequency_lut.rng[3] ),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_4 _2138_ (.A(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _2139_ (.A0(_0545_),
    .A1(_0550_),
    .S(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__inv_2 _2140_ (.A(\inputs.frequency_lut.rng[3] ),
    .Y(_0554_));
 sky130_fd_sc_hd__clkbuf_4 _2141_ (.A(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_4 _2142_ (.A(\inputs.frequency_lut.rng[0] ),
    .X(_0556_));
 sky130_fd_sc_hd__a21o_1 _2143_ (.A1(_0556_),
    .A2(_0543_),
    .B1(_0536_),
    .X(_0557_));
 sky130_fd_sc_hd__nor2_1 _2144_ (.A(_0556_),
    .B(_0543_),
    .Y(_0558_));
 sky130_fd_sc_hd__nand2_2 _2145_ (.A(_0537_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__o21ai_1 _2146_ (.A1(_0555_),
    .A2(_0557_),
    .B1(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__clkbuf_4 _2147_ (.A(_0551_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_4 _2148_ (.A(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__or2_1 _2149_ (.A(_0535_),
    .B(_0540_),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_4 _2150_ (.A(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _2151_ (.A(_0536_),
    .B(_0542_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_1 _2152_ (.A(_0564_),
    .B(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__nand2_2 _2153_ (.A(_0537_),
    .B(_0540_),
    .Y(_0567_));
 sky130_fd_sc_hd__clkbuf_4 _2154_ (.A(\inputs.frequency_lut.rng[3] ),
    .X(_0568_));
 sky130_fd_sc_hd__clkbuf_4 _2155_ (.A(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__a21oi_1 _2156_ (.A1(_0564_),
    .A2(_0567_),
    .B1(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__a21oi_1 _2157_ (.A1(_0562_),
    .A2(_0566_),
    .B1(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__nor2_1 _2158_ (.A(_0543_),
    .B(_0536_),
    .Y(_0572_));
 sky130_fd_sc_hd__nor2_1 _2159_ (.A(_0556_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__a21oi_1 _2160_ (.A1(_0562_),
    .A2(_0547_),
    .B1(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_2 _2161_ (.A(\inputs.frequency_lut.rng[4] ),
    .Y(_0575_));
 sky130_fd_sc_hd__clkbuf_4 _2162_ (.A(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__inv_2 _2163_ (.A(\inputs.frequency_lut.rng[5] ),
    .Y(_0577_));
 sky130_fd_sc_hd__clkbuf_4 _2164_ (.A(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__mux4_1 _2165_ (.A0(_0553_),
    .A1(_0560_),
    .A2(_0571_),
    .A3(_0574_),
    .S0(_0576_),
    .S1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__inv_2 _2166_ (.A(\inputs.key_encoder.sync_keys[2] ),
    .Y(_0580_));
 sky130_fd_sc_hd__a21oi_1 _2167_ (.A1(\inputs.key_encoder.sync_keys[1] ),
    .A2(_0580_),
    .B1(\inputs.key_encoder.sync_keys[3] ),
    .Y(_0581_));
 sky130_fd_sc_hd__o21ba_1 _2168_ (.A1(\inputs.key_encoder.sync_keys[4] ),
    .A2(_0581_),
    .B1_N(\inputs.key_encoder.sync_keys[5] ),
    .X(_0582_));
 sky130_fd_sc_hd__o21ba_1 _2169_ (.A1(\inputs.key_encoder.sync_keys[6] ),
    .A2(_0582_),
    .B1_N(\inputs.key_encoder.sync_keys[7] ),
    .X(_0583_));
 sky130_fd_sc_hd__o21ba_1 _2170_ (.A1(\inputs.key_encoder.sync_keys[8] ),
    .A2(_0583_),
    .B1_N(\inputs.key_encoder.sync_keys[9] ),
    .X(_0584_));
 sky130_fd_sc_hd__o21bai_4 _2171_ (.A1(\inputs.key_encoder.sync_keys[10] ),
    .A2(_0584_),
    .B1_N(\inputs.key_encoder.sync_keys[11] ),
    .Y(_0585_));
 sky130_fd_sc_hd__and2b_1 _2172_ (.A_N(\inputs.key_encoder.sync_keys[13] ),
    .B(_1287_),
    .X(_0586_));
 sky130_fd_sc_hd__o31a_1 _2173_ (.A1(\inputs.key_encoder.sync_keys[12] ),
    .A2(_1288_),
    .A3(_1291_),
    .B1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__nor2_1 _2174_ (.A(\inputs.key_encoder.sync_keys[8] ),
    .B(\inputs.key_encoder.sync_keys[9] ),
    .Y(_0588_));
 sky130_fd_sc_hd__nor2_1 _2175_ (.A(\inputs.key_encoder.sync_keys[4] ),
    .B(\inputs.key_encoder.sync_keys[5] ),
    .Y(_0589_));
 sky130_fd_sc_hd__a211o_1 _2176_ (.A1(_1289_),
    .A2(_0589_),
    .B1(\inputs.key_encoder.sync_keys[6] ),
    .C1(\inputs.key_encoder.sync_keys[7] ),
    .X(_0590_));
 sky130_fd_sc_hd__a211o_2 _2177_ (.A1(_0588_),
    .A2(_0590_),
    .B1(\inputs.key_encoder.sync_keys[11] ),
    .C1(\inputs.key_encoder.sync_keys[10] ),
    .X(_0591_));
 sky130_fd_sc_hd__nor2b_2 _2178_ (.A(\inputs.key_encoder.sync_keys[12] ),
    .B_N(_0586_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _2179_ (.A(_0591_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__or2_1 _2180_ (.A(_0587_),
    .B(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__inv_2 _2181_ (.A(_1288_),
    .Y(_0595_));
 sky130_fd_sc_hd__and2_1 _2182_ (.A(_0595_),
    .B(_1291_),
    .X(_0596_));
 sky130_fd_sc_hd__nand2_2 _2183_ (.A(_0596_),
    .B(_0592_),
    .Y(_0597_));
 sky130_fd_sc_hd__or2_2 _2184_ (.A(_0591_),
    .B(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__or3_1 _2185_ (.A(_0595_),
    .B(_0585_),
    .C(_0593_),
    .X(_0599_));
 sky130_fd_sc_hd__nand2_1 _2186_ (.A(_0585_),
    .B(_0592_),
    .Y(_0600_));
 sky130_fd_sc_hd__or3_4 _2187_ (.A(_0587_),
    .B(_0591_),
    .C(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__o2111ai_2 _2188_ (.A1(_0585_),
    .A2(_0594_),
    .B1(_0598_),
    .C1(_0599_),
    .D1(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__and2_2 _2189_ (.A(\inputs.key_encoder.sync_keys[13] ),
    .B(_1287_),
    .X(_0603_));
 sky130_fd_sc_hd__or2_1 _2190_ (.A(_0603_),
    .B(_0587_),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_1 _2191_ (.A(_0600_),
    .B(_0593_),
    .Y(_0605_));
 sky130_fd_sc_hd__or2_1 _2192_ (.A(_0604_),
    .B(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__o211a_1 _2193_ (.A1(_0600_),
    .A2(_0598_),
    .B1(_0606_),
    .C1(_0601_),
    .X(_0607_));
 sky130_fd_sc_hd__or3b_1 _2194_ (.A(_0595_),
    .B(_0585_),
    .C_N(_0592_),
    .X(_0608_));
 sky130_fd_sc_hd__nand2b_1 _2195_ (.A_N(_0594_),
    .B(_0585_),
    .Y(_0609_));
 sky130_fd_sc_hd__and3_1 _2196_ (.A(_0607_),
    .B(_0608_),
    .C(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__buf_2 _2197_ (.A(_0237_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _2198_ (.A0(_0602_),
    .A1(_0610_),
    .S(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__o21a_1 _2199_ (.A1(\inputs.key_encoder.sync_keys[12] ),
    .A2(_0596_),
    .B1(_0586_),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_1 _2200_ (.A(_0613_),
    .B(_0598_),
    .Y(_0614_));
 sky130_fd_sc_hd__and2_1 _2201_ (.A(_0601_),
    .B(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__or3_2 _2202_ (.A(_0595_),
    .B(_0591_),
    .C(_0600_),
    .X(_0616_));
 sky130_fd_sc_hd__and3_1 _2203_ (.A(_0599_),
    .B(_0614_),
    .C(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _2204_ (.A(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__nor2_1 _2205_ (.A(_0591_),
    .B(_0608_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_1 _2206_ (.A(_0585_),
    .B(_0598_),
    .Y(_0620_));
 sky130_fd_sc_hd__or4b_1 _2207_ (.A(_0618_),
    .B(_0619_),
    .C(_0620_),
    .D_N(_0604_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(_0615_),
    .A1(_0621_),
    .S(_0238_),
    .X(_0622_));
 sky130_fd_sc_hd__a21o_1 _2209_ (.A1(\inputs.octave_fsm.state[0] ),
    .A2(\inputs.octave_fsm.state[2] ),
    .B1(\inputs.octave_fsm.state[1] ),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_4 _2210_ (.A(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _2211_ (.A0(_0612_),
    .A1(_0622_),
    .S(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__a21oi_4 _2212_ (.A1(\inputs.octave_fsm.state[0] ),
    .A2(\inputs.octave_fsm.state[2] ),
    .B1(\inputs.octave_fsm.state[1] ),
    .Y(_0626_));
 sky130_fd_sc_hd__or2b_1 _2213_ (.A(_0600_),
    .B_N(_0591_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_1 _2214_ (.A(_0604_),
    .B(_0605_),
    .Y(_0628_));
 sky130_fd_sc_hd__a311o_1 _2215_ (.A1(_0596_),
    .A2(_0592_),
    .A3(_0627_),
    .B1(_0619_),
    .C1(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _2216_ (.A(_0597_),
    .B(_0627_),
    .Y(_0630_));
 sky130_fd_sc_hd__or2_1 _2217_ (.A(_0585_),
    .B(_0598_),
    .X(_0631_));
 sky130_fd_sc_hd__nand2_1 _2218_ (.A(_0594_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__or3_1 _2219_ (.A(_0628_),
    .B(_0630_),
    .C(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(_0629_),
    .A1(_0633_),
    .S(_0238_),
    .X(_0634_));
 sky130_fd_sc_hd__inv_2 _2221_ (.A(_0601_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2_1 _2222_ (.A(_0609_),
    .B(_0631_),
    .Y(_0636_));
 sky130_fd_sc_hd__a31o_1 _2223_ (.A1(_0596_),
    .A2(_0591_),
    .A3(_0592_),
    .B1(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__or3b_1 _2224_ (.A(_0635_),
    .B(_0637_),
    .C_N(_0616_),
    .X(_0638_));
 sky130_fd_sc_hd__a31oi_1 _2225_ (.A1(_0607_),
    .A2(_0609_),
    .A3(_0614_),
    .B1(_0611_),
    .Y(_0639_));
 sky130_fd_sc_hd__a211o_1 _2226_ (.A1(_0611_),
    .A2(_0638_),
    .B1(_0639_),
    .C1(_0624_),
    .X(_0640_));
 sky130_fd_sc_hd__o211a_1 _2227_ (.A1(_0626_),
    .A2(_0634_),
    .B1(_0640_),
    .C1(_0230_),
    .X(_0641_));
 sky130_fd_sc_hd__clkbuf_4 _2228_ (.A(_0603_),
    .X(_0642_));
 sky130_fd_sc_hd__a211o_1 _2229_ (.A1(_0247_),
    .A2(_0625_),
    .B1(_0641_),
    .C1(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__o21ai_1 _2230_ (.A1(_0534_),
    .A2(_0579_),
    .B1(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__clkbuf_4 _2231_ (.A(_0512_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(net317),
    .A1(_0644_),
    .S(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(_0646_),
    .X(_0113_));
 sky130_fd_sc_hd__o21ai_1 _2234_ (.A1(_0554_),
    .A2(_0558_),
    .B1(_0540_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_2 _2235_ (.A(_0551_),
    .B(_0544_),
    .Y(_0648_));
 sky130_fd_sc_hd__o22a_1 _2236_ (.A1(_0547_),
    .A2(_0647_),
    .B1(_0648_),
    .B2(_0538_),
    .X(_0649_));
 sky130_fd_sc_hd__nor2_2 _2237_ (.A(_0536_),
    .B(_0558_),
    .Y(_0650_));
 sky130_fd_sc_hd__or2b_1 _2238_ (.A(_0535_),
    .B_N(_0543_),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_2 _2239_ (.A(_0535_),
    .B(_0541_),
    .Y(_0652_));
 sky130_fd_sc_hd__and2_1 _2240_ (.A(_0651_),
    .B(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__nand2_1 _2241_ (.A(_0561_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__o31a_1 _2242_ (.A1(_0561_),
    .A2(_0549_),
    .A3(_0650_),
    .B1(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__and3_2 _2243_ (.A(\inputs.frequency_lut.rng[0] ),
    .B(\inputs.frequency_lut.rng[1] ),
    .C(\inputs.frequency_lut.rng[2] ),
    .X(_0656_));
 sky130_fd_sc_hd__a21oi_4 _2244_ (.A1(_0556_),
    .A2(\inputs.frequency_lut.rng[1] ),
    .B1(\inputs.frequency_lut.rng[2] ),
    .Y(_0657_));
 sky130_fd_sc_hd__nor2_1 _2245_ (.A(_0551_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__and2b_1 _2246_ (.A_N(_0535_),
    .B(_0543_),
    .X(_0659_));
 sky130_fd_sc_hd__nand2_1 _2247_ (.A(_0554_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__o32a_1 _2248_ (.A1(_0650_),
    .A2(_0656_),
    .A3(_0658_),
    .B1(_0660_),
    .B2(_0538_),
    .X(_0661_));
 sky130_fd_sc_hd__nor2_2 _2249_ (.A(_0556_),
    .B(_0535_),
    .Y(_0662_));
 sky130_fd_sc_hd__nor2_1 _2250_ (.A(_0551_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__a21oi_1 _2251_ (.A1(_0564_),
    .A2(_0567_),
    .B1(_0555_),
    .Y(_0664_));
 sky130_fd_sc_hd__a21oi_1 _2252_ (.A1(_0565_),
    .A2(_0663_),
    .B1(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__mux4_1 _2253_ (.A0(_0649_),
    .A1(_0655_),
    .A2(_0661_),
    .A3(_0665_),
    .S0(_0576_),
    .S1(_0578_),
    .X(_0666_));
 sky130_fd_sc_hd__a31o_1 _2254_ (.A1(_0598_),
    .A2(_0599_),
    .A3(_0616_),
    .B1(_0632_),
    .X(_0667_));
 sky130_fd_sc_hd__and3_1 _2255_ (.A(_0601_),
    .B(_0606_),
    .C(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(_0615_),
    .A1(_0668_),
    .S(_0237_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _2257_ (.A0(_0610_),
    .A1(_0621_),
    .S(_0611_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _2258_ (.A0(_0669_),
    .A1(_0670_),
    .S(_0626_),
    .X(_0671_));
 sky130_fd_sc_hd__nor2_1 _2259_ (.A(_0230_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__mux4_1 _2260_ (.A0(_0602_),
    .A1(_0629_),
    .A2(_0633_),
    .A3(_0638_),
    .S0(_0238_),
    .S1(_0626_),
    .X(_0673_));
 sky130_fd_sc_hd__buf_2 _2261_ (.A(_0533_),
    .X(_0674_));
 sky130_fd_sc_hd__o21ai_1 _2262_ (.A1(_0247_),
    .A2(_0673_),
    .B1(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__o22a_1 _2263_ (.A1(_0534_),
    .A2(_0666_),
    .B1(_0672_),
    .B2(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _2264_ (.A0(net310),
    .A1(_0676_),
    .S(_0645_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _2265_ (.A(_0677_),
    .X(_0114_));
 sky130_fd_sc_hd__and4_1 _2266_ (.A(_0601_),
    .B(_0598_),
    .C(_0609_),
    .D(_0617_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _2267_ (.A0(_0668_),
    .A1(_0678_),
    .S(_0237_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _2268_ (.A0(_0622_),
    .A1(_0679_),
    .S(_0624_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _2269_ (.A0(_0612_),
    .A1(_0634_),
    .S(_0626_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _2270_ (.A0(_0680_),
    .A1(_0681_),
    .S(_0230_),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_1 _2271_ (.A(_0555_),
    .B(_0545_),
    .Y(_0683_));
 sky130_fd_sc_hd__a21o_1 _2272_ (.A1(_0559_),
    .A2(_0658_),
    .B1(_0576_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_4 _2273_ (.A(\inputs.frequency_lut.rng[4] ),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_4 _2274_ (.A(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__a211o_1 _2275_ (.A1(_0569_),
    .A2(_0559_),
    .B1(_0566_),
    .C1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__o211a_1 _2276_ (.A1(_0683_),
    .A2(_0684_),
    .B1(_0687_),
    .C1(_0578_),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_1 _2277_ (.A(_0685_),
    .B(_0647_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _2278_ (.A(_0538_),
    .B(_0536_),
    .Y(_0690_));
 sky130_fd_sc_hd__nor2_1 _2279_ (.A(_0568_),
    .B(_0541_),
    .Y(_0691_));
 sky130_fd_sc_hd__a31o_1 _2280_ (.A1(_0552_),
    .A2(_0564_),
    .A3(_0690_),
    .B1(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__o32a_1 _2281_ (.A1(_0657_),
    .A2(_0656_),
    .A3(_0689_),
    .B1(_0692_),
    .B2(_0686_),
    .X(_0693_));
 sky130_fd_sc_hd__o21ai_1 _2282_ (.A1(_0578_),
    .A2(_0693_),
    .B1(_0603_),
    .Y(_0694_));
 sky130_fd_sc_hd__o2bb2a_1 _2283_ (.A1_N(_0534_),
    .A2_N(_0682_),
    .B1(_0688_),
    .B2(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _2284_ (.A0(net279),
    .A1(_0695_),
    .S(_0645_),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_1 _2285_ (.A(_0696_),
    .X(_0115_));
 sky130_fd_sc_hd__o221a_1 _2286_ (.A1(\inputs.key_encoder.sync_keys[12] ),
    .A2(_1288_),
    .B1(_0596_),
    .B2(_0593_),
    .C1(_0586_),
    .X(_0697_));
 sky130_fd_sc_hd__or3_1 _2287_ (.A(_0635_),
    .B(_0620_),
    .C(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _2288_ (.A0(_0678_),
    .A1(_0698_),
    .S(_0237_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _2289_ (.A0(_0669_),
    .A1(_0699_),
    .S(_0623_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _2290_ (.A0(_0602_),
    .A1(_0629_),
    .S(_0238_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(_0670_),
    .A1(_0701_),
    .S(_0626_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _2292_ (.A0(_0700_),
    .A1(_0702_),
    .S(_0230_),
    .X(_0703_));
 sky130_fd_sc_hd__inv_2 _2293_ (.A(_0656_),
    .Y(_0704_));
 sky130_fd_sc_hd__a31o_1 _2294_ (.A1(_0561_),
    .A2(_0564_),
    .A3(_0704_),
    .B1(_0663_),
    .X(_0705_));
 sky130_fd_sc_hd__or2b_1 _2295_ (.A(\inputs.frequency_lut.rng[1] ),
    .B_N(\inputs.frequency_lut.rng[2] ),
    .X(_0706_));
 sky130_fd_sc_hd__nor2_1 _2296_ (.A(_0554_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__a31oi_1 _2297_ (.A1(_0651_),
    .A2(_0663_),
    .A3(_0706_),
    .B1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__and2_1 _2298_ (.A(_0538_),
    .B(_0707_),
    .X(_0709_));
 sky130_fd_sc_hd__nor3_1 _2299_ (.A(_0650_),
    .B(_0656_),
    .C(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o22a_1 _2300_ (.A1(_0573_),
    .A2(_0648_),
    .B1(_0653_),
    .B2(_0561_),
    .X(_0711_));
 sky130_fd_sc_hd__mux4_1 _2301_ (.A0(_0705_),
    .A1(_0708_),
    .A2(_0710_),
    .A3(_0711_),
    .S0(_0685_),
    .S1(_0577_),
    .X(_0712_));
 sky130_fd_sc_hd__or2_1 _2302_ (.A(_0674_),
    .B(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__o21ai_1 _2303_ (.A1(_0642_),
    .A2(_0703_),
    .B1(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__mux2_1 _2304_ (.A0(net318),
    .A1(_0714_),
    .S(_0645_),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_1 _2305_ (.A(_0715_),
    .X(_0116_));
 sky130_fd_sc_hd__nor2_1 _2306_ (.A(_0685_),
    .B(_0550_),
    .Y(_0716_));
 sky130_fd_sc_hd__and3b_2 _2307_ (.A_N(_0543_),
    .B(_0535_),
    .C(_0556_),
    .X(_0717_));
 sky130_fd_sc_hd__nand3_1 _2308_ (.A(_0554_),
    .B(_0564_),
    .C(_0690_),
    .Y(_0718_));
 sky130_fd_sc_hd__o21a_1 _2309_ (.A1(_0555_),
    .A2(_0717_),
    .B1(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__a21oi_1 _2310_ (.A1(_0716_),
    .A2(_0719_),
    .B1(\inputs.frequency_lut.rng[5] ),
    .Y(_0720_));
 sky130_fd_sc_hd__o21a_1 _2311_ (.A1(_0716_),
    .A2(_0719_),
    .B1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__a21oi_2 _2312_ (.A1(_0539_),
    .A2(_0541_),
    .B1(_0535_),
    .Y(_0722_));
 sky130_fd_sc_hd__o21a_1 _2313_ (.A1(_0549_),
    .A2(_0722_),
    .B1(_0569_),
    .X(_0723_));
 sky130_fd_sc_hd__o21a_1 _2314_ (.A1(_0572_),
    .A2(_0717_),
    .B1(_0554_),
    .X(_0724_));
 sky130_fd_sc_hd__a21oi_1 _2315_ (.A1(_0561_),
    .A2(_0659_),
    .B1(_0685_),
    .Y(_0725_));
 sky130_fd_sc_hd__a21bo_1 _2316_ (.A1(_0567_),
    .A2(_0658_),
    .B1_N(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_4 _2317_ (.A(\inputs.frequency_lut.rng[5] ),
    .X(_0727_));
 sky130_fd_sc_hd__o311a_1 _2318_ (.A1(_0576_),
    .A2(_0723_),
    .A3(_0724_),
    .B1(_0726_),
    .C1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _2319_ (.A(_0591_),
    .B(_0597_),
    .Y(_0729_));
 sky130_fd_sc_hd__o21a_1 _2320_ (.A1(_0585_),
    .A2(_0597_),
    .B1(_0616_),
    .X(_0730_));
 sky130_fd_sc_hd__o21ai_1 _2321_ (.A1(_0729_),
    .A2(_0730_),
    .B1(_0604_),
    .Y(_0731_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(_0698_),
    .A1(_0731_),
    .S(_0611_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _2323_ (.A0(_0679_),
    .A1(_0732_),
    .S(_0624_),
    .X(_0733_));
 sky130_fd_sc_hd__nor2_1 _2324_ (.A(_0230_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__o21ai_1 _2325_ (.A1(_0247_),
    .A2(_0625_),
    .B1(_0674_),
    .Y(_0735_));
 sky130_fd_sc_hd__o32a_1 _2326_ (.A1(_0674_),
    .A2(_0721_),
    .A3(_0728_),
    .B1(_0734_),
    .B2(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _2327_ (.A0(net311),
    .A1(_0736_),
    .S(_0645_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_1 _2328_ (.A(_0737_),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _2329_ (.A(_0556_),
    .B(_0537_),
    .X(_0738_));
 sky130_fd_sc_hd__a31o_1 _2330_ (.A1(_0568_),
    .A2(_0538_),
    .A3(_0659_),
    .B1(_0663_),
    .X(_0739_));
 sky130_fd_sc_hd__a211o_1 _2331_ (.A1(_0738_),
    .A2(_0653_),
    .B1(_0739_),
    .C1(_0575_),
    .X(_0740_));
 sky130_fd_sc_hd__nor2_1 _2332_ (.A(_0561_),
    .B(_0706_),
    .Y(_0741_));
 sky130_fd_sc_hd__a211o_1 _2333_ (.A1(_0569_),
    .A2(_0566_),
    .B1(_0741_),
    .C1(_0686_),
    .X(_0742_));
 sky130_fd_sc_hd__nor2_1 _2334_ (.A(_0551_),
    .B(_0547_),
    .Y(_0743_));
 sky130_fd_sc_hd__o2bb2a_1 _2335_ (.A1_N(_0565_),
    .A2_N(_0743_),
    .B1(_0555_),
    .B2(_0662_),
    .X(_0744_));
 sky130_fd_sc_hd__or2_1 _2336_ (.A(\inputs.frequency_lut.rng[3] ),
    .B(_0656_),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_1 _2337_ (.A(_0648_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__a31o_1 _2338_ (.A1(_0685_),
    .A2(_0564_),
    .A3(_0746_),
    .B1(\inputs.frequency_lut.rng[5] ),
    .X(_0747_));
 sky130_fd_sc_hd__o21ba_1 _2339_ (.A1(_0686_),
    .A2(_0744_),
    .B1_N(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__a31o_1 _2340_ (.A1(_0727_),
    .A2(_0740_),
    .A3(_0742_),
    .B1(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__nand2_1 _2341_ (.A(_0231_),
    .B(_0671_),
    .Y(_0750_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(_0618_),
    .A1(_0731_),
    .S(_0238_),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(_0699_),
    .A1(_0751_),
    .S(_0624_),
    .X(_0752_));
 sky130_fd_sc_hd__a21oi_1 _2344_ (.A1(_0247_),
    .A2(_0752_),
    .B1(_0642_),
    .Y(_0753_));
 sky130_fd_sc_hd__a22o_1 _2345_ (.A1(_0642_),
    .A2(_0749_),
    .B1(_0750_),
    .B2(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(\outputs.div.divisor[5] ),
    .A1(_0754_),
    .S(_0645_),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_1 _2347_ (.A(_0755_),
    .X(_0118_));
 sky130_fd_sc_hd__o21a_1 _2348_ (.A1(_0585_),
    .A2(_0593_),
    .B1(_0597_),
    .X(_0756_));
 sky130_fd_sc_hd__a31o_1 _2349_ (.A1(_0613_),
    .A2(_0605_),
    .A3(_0627_),
    .B1(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__and2_1 _2350_ (.A(_0606_),
    .B(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(_0617_),
    .A1(_0758_),
    .S(_0611_),
    .X(_0759_));
 sky130_fd_sc_hd__nand2_1 _2352_ (.A(_0626_),
    .B(_0732_),
    .Y(_0760_));
 sky130_fd_sc_hd__o21a_1 _2353_ (.A1(_0626_),
    .A2(_0759_),
    .B1(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__nand2_1 _2354_ (.A(_0231_),
    .B(_0680_),
    .Y(_0762_));
 sky130_fd_sc_hd__o211a_1 _2355_ (.A1(_0231_),
    .A2(_0761_),
    .B1(_0762_),
    .C1(_0534_),
    .X(_0763_));
 sky130_fd_sc_hd__and2_1 _2356_ (.A(\inputs.frequency_lut.rng[0] ),
    .B(\inputs.frequency_lut.rng[2] ),
    .X(_0764_));
 sky130_fd_sc_hd__or3_1 _2357_ (.A(_0568_),
    .B(_0722_),
    .C(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__nand2_1 _2358_ (.A(_0568_),
    .B(_0537_),
    .Y(_0766_));
 sky130_fd_sc_hd__or2_1 _2359_ (.A(_0542_),
    .B(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_4 _2360_ (.A(_0686_),
    .X(_0768_));
 sky130_fd_sc_hd__a41o_1 _2361_ (.A1(_0768_),
    .A2(_0559_),
    .A3(_0564_),
    .A4(_0654_),
    .B1(_0578_),
    .X(_0769_));
 sky130_fd_sc_hd__a31o_1 _2362_ (.A1(_0576_),
    .A2(_0765_),
    .A3(_0767_),
    .B1(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__o21ai_1 _2363_ (.A1(_0572_),
    .A2(_0717_),
    .B1(_0562_),
    .Y(_0771_));
 sky130_fd_sc_hd__a311oi_1 _2364_ (.A1(_0562_),
    .A2(_0557_),
    .A3(_0567_),
    .B1(_0717_),
    .C1(_0768_),
    .Y(_0772_));
 sky130_fd_sc_hd__a31o_1 _2365_ (.A1(_0768_),
    .A2(_0660_),
    .A3(_0771_),
    .B1(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__a21oi_1 _2366_ (.A1(_0578_),
    .A2(_0773_),
    .B1(_0534_),
    .Y(_0774_));
 sky130_fd_sc_hd__a21bo_1 _2367_ (.A1(_0770_),
    .A2(_0774_),
    .B1_N(_0513_),
    .X(_0775_));
 sky130_fd_sc_hd__o22a_1 _2368_ (.A1(net208),
    .A2(_0513_),
    .B1(_0763_),
    .B2(_0775_),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _2369_ (.A(_0536_),
    .B(_0540_),
    .X(_0776_));
 sky130_fd_sc_hd__o32a_1 _2370_ (.A1(_0561_),
    .A2(_0776_),
    .A3(_0722_),
    .B1(_0650_),
    .B2(_0648_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _2371_ (.A(_0561_),
    .B(_0540_),
    .Y(_0778_));
 sky130_fd_sc_hd__a22oi_1 _2372_ (.A1(_0552_),
    .A2(_0764_),
    .B1(_0778_),
    .B2(_0652_),
    .Y(_0779_));
 sky130_fd_sc_hd__a21oi_1 _2373_ (.A1(_0563_),
    .A2(_0704_),
    .B1(_0568_),
    .Y(_0780_));
 sky130_fd_sc_hd__or2_1 _2374_ (.A(_0707_),
    .B(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__o21ba_1 _2375_ (.A1(_0552_),
    .A2(_0542_),
    .B1_N(_0662_),
    .X(_0782_));
 sky130_fd_sc_hd__mux4_1 _2376_ (.A0(_0777_),
    .A1(_0779_),
    .A2(_0781_),
    .A3(_0782_),
    .S0(_0686_),
    .S1(_0578_),
    .X(_0783_));
 sky130_fd_sc_hd__a311o_1 _2377_ (.A1(_1288_),
    .A2(_0592_),
    .A3(_0627_),
    .B1(_0636_),
    .C1(_0628_),
    .X(_0784_));
 sky130_fd_sc_hd__or2_1 _2378_ (.A(_0611_),
    .B(_0758_),
    .X(_0785_));
 sky130_fd_sc_hd__o21ai_1 _2379_ (.A1(_0238_),
    .A2(_0784_),
    .B1(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(_0751_),
    .A1(_0786_),
    .S(_0624_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_1 _2381_ (.A(_0229_),
    .B(_0700_),
    .X(_0788_));
 sky130_fd_sc_hd__a21oi_1 _2382_ (.A1(_0247_),
    .A2(_0787_),
    .B1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(_0783_),
    .A1(_0789_),
    .S(_0674_),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(\outputs.div.divisor[7] ),
    .A1(_0790_),
    .S(_0645_),
    .X(_0791_));
 sky130_fd_sc_hd__clkbuf_1 _2385_ (.A(_0791_),
    .X(_0120_));
 sky130_fd_sc_hd__o21a_1 _2386_ (.A1(_0722_),
    .A2(_0764_),
    .B1(_0551_),
    .X(_0792_));
 sky130_fd_sc_hd__or2_1 _2387_ (.A(_0724_),
    .B(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__nor2_1 _2388_ (.A(_0568_),
    .B(_0549_),
    .Y(_0794_));
 sky130_fd_sc_hd__a31o_1 _2389_ (.A1(_0552_),
    .A2(_0559_),
    .A3(_0564_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__nand3_1 _2390_ (.A(_0551_),
    .B(_0536_),
    .C(_0540_),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _2391_ (.A(_0660_),
    .B(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__a21o_1 _2392_ (.A1(_0552_),
    .A2(_0547_),
    .B1(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__a21o_1 _2393_ (.A1(_0540_),
    .A2(_0547_),
    .B1(_0764_),
    .X(_0799_));
 sky130_fd_sc_hd__and2_1 _2394_ (.A(_0554_),
    .B(_0544_),
    .X(_0800_));
 sky130_fd_sc_hd__a21o_1 _2395_ (.A1(_0552_),
    .A2(_0799_),
    .B1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__mux4_1 _2396_ (.A0(_0793_),
    .A1(_0795_),
    .A2(_0798_),
    .A3(_0801_),
    .S0(_0686_),
    .S1(_0727_),
    .X(_0802_));
 sky130_fd_sc_hd__nand2_1 _2397_ (.A(_0231_),
    .B(_0733_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_1 _2398_ (.A(_0597_),
    .B(_0609_),
    .Y(_0804_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(_0784_),
    .A1(_0804_),
    .S(_0611_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _2400_ (.A0(_0759_),
    .A1(_0805_),
    .S(_0624_),
    .X(_0806_));
 sky130_fd_sc_hd__o21a_1 _2401_ (.A1(_0230_),
    .A2(_0806_),
    .B1(_0674_),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _2402_ (.A1(_0642_),
    .A2(_0802_),
    .B1(_0803_),
    .B2(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(\outputs.div.divisor[8] ),
    .A1(_0808_),
    .S(_0645_),
    .X(_0809_));
 sky130_fd_sc_hd__clkbuf_1 _2404_ (.A(_0809_),
    .X(_0121_));
 sky130_fd_sc_hd__or3_1 _2405_ (.A(_0568_),
    .B(_0549_),
    .C(_0662_),
    .X(_0810_));
 sky130_fd_sc_hd__and2_1 _2406_ (.A(_0538_),
    .B(_0536_),
    .X(_0811_));
 sky130_fd_sc_hd__o21ai_1 _2407_ (.A1(_0547_),
    .A2(_0811_),
    .B1(_0569_),
    .Y(_0812_));
 sky130_fd_sc_hd__a21o_1 _2408_ (.A1(_0810_),
    .A2(_0812_),
    .B1(_0577_),
    .X(_0813_));
 sky130_fd_sc_hd__inv_2 _2409_ (.A(_0650_),
    .Y(_0814_));
 sky130_fd_sc_hd__a221o_1 _2410_ (.A1(_0569_),
    .A2(_0652_),
    .B1(_0800_),
    .B2(_0814_),
    .C1(\inputs.frequency_lut.rng[5] ),
    .X(_0815_));
 sky130_fd_sc_hd__and3_1 _2411_ (.A(_0768_),
    .B(_0813_),
    .C(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__inv_2 _2412_ (.A(_0722_),
    .Y(_0817_));
 sky130_fd_sc_hd__or3_1 _2413_ (.A(_0568_),
    .B(_0549_),
    .C(_0572_),
    .X(_0818_));
 sky130_fd_sc_hd__a311o_1 _2414_ (.A1(_0567_),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0691_),
    .C1(\inputs.frequency_lut.rng[5] ),
    .X(_0819_));
 sky130_fd_sc_hd__or3_1 _2415_ (.A(_0555_),
    .B(_0549_),
    .C(_0572_),
    .X(_0820_));
 sky130_fd_sc_hd__o211ai_1 _2416_ (.A1(_0562_),
    .A2(_0564_),
    .B1(_0820_),
    .C1(_0727_),
    .Y(_0821_));
 sky130_fd_sc_hd__a31o_1 _2417_ (.A1(_0576_),
    .A2(_0819_),
    .A3(_0821_),
    .B1(_0674_),
    .X(_0822_));
 sky130_fd_sc_hd__o211a_2 _2418_ (.A1(_0585_),
    .A2(_0594_),
    .B1(_0606_),
    .C1(_0601_),
    .X(_0823_));
 sky130_fd_sc_hd__o21ai_1 _2419_ (.A1(_0611_),
    .A2(_0804_),
    .B1(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(_0786_),
    .A1(_0824_),
    .S(_0624_),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(_0752_),
    .A1(_0825_),
    .S(_0247_),
    .X(_0826_));
 sky130_fd_sc_hd__o22ai_1 _2422_ (.A1(_0816_),
    .A2(_0822_),
    .B1(_0826_),
    .B2(_0642_),
    .Y(_0827_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(net253),
    .A1(_0827_),
    .S(_0645_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_1 _2424_ (.A(_0828_),
    .X(_0122_));
 sky130_fd_sc_hd__xnor2_1 _2425_ (.A(_0238_),
    .B(_0823_),
    .Y(_0829_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(_0805_),
    .A1(_0829_),
    .S(_0624_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(_0761_),
    .A1(_0830_),
    .S(_0247_),
    .X(_0831_));
 sky130_fd_sc_hd__o21a_1 _2428_ (.A1(_0657_),
    .A2(_0764_),
    .B1(\inputs.frequency_lut.rng[3] ),
    .X(_0832_));
 sky130_fd_sc_hd__a31o_1 _2429_ (.A1(_0540_),
    .A2(_0541_),
    .A3(_0800_),
    .B1(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__a31o_1 _2430_ (.A1(_0551_),
    .A2(_0652_),
    .A3(_0817_),
    .B1(_0685_),
    .X(_0834_));
 sky130_fd_sc_hd__nor2_1 _2431_ (.A(_0561_),
    .B(_0799_),
    .Y(_0835_));
 sky130_fd_sc_hd__o2bb2a_1 _2432_ (.A1_N(_0685_),
    .A2_N(_0833_),
    .B1(_0834_),
    .B2(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__o21ai_1 _2433_ (.A1(_0547_),
    .A2(_0776_),
    .B1(_0555_),
    .Y(_0837_));
 sky130_fd_sc_hd__a32o_1 _2434_ (.A1(_0685_),
    .A2(_0648_),
    .A3(_0837_),
    .B1(_0725_),
    .B2(_0718_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(_0836_),
    .A1(_0838_),
    .S(_0578_),
    .X(_0839_));
 sky130_fd_sc_hd__nor2_1 _2436_ (.A(_0674_),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__a21o_1 _2437_ (.A1(_0534_),
    .A2(_0831_),
    .B1(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(\outputs.div.divisor[10] ),
    .A1(_0841_),
    .S(_0645_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_1 _2439_ (.A(_0842_),
    .X(_0123_));
 sky130_fd_sc_hd__nor2_1 _2440_ (.A(_0658_),
    .B(_0811_),
    .Y(_0843_));
 sky130_fd_sc_hd__or3_1 _2441_ (.A(_0554_),
    .B(_0650_),
    .C(_0656_),
    .X(_0844_));
 sky130_fd_sc_hd__o21a_1 _2442_ (.A1(_0569_),
    .A2(_0550_),
    .B1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__o21ai_1 _2443_ (.A1(_0549_),
    .A2(_0662_),
    .B1(_0562_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _2444_ (.A(_0818_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__a21oi_1 _2445_ (.A1(_0562_),
    .A2(_0540_),
    .B1(_0537_),
    .Y(_0848_));
 sky130_fd_sc_hd__mux4_1 _2446_ (.A0(_0843_),
    .A1(_0845_),
    .A2(_0847_),
    .A3(_0848_),
    .S0(_0576_),
    .S1(_0578_),
    .X(_0849_));
 sky130_fd_sc_hd__or3_1 _2447_ (.A(_0611_),
    .B(_0626_),
    .C(_0823_),
    .X(_0850_));
 sky130_fd_sc_hd__o21ai_1 _2448_ (.A1(_0624_),
    .A2(_0824_),
    .B1(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__nor2_1 _2449_ (.A(_0230_),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__a211o_1 _2450_ (.A1(_0230_),
    .A2(_0787_),
    .B1(_0852_),
    .C1(_0642_),
    .X(_0853_));
 sky130_fd_sc_hd__o21ai_1 _2451_ (.A1(_0534_),
    .A2(_0849_),
    .B1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__buf_4 _2452_ (.A(_0512_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(\outputs.div.divisor[11] ),
    .A1(_0854_),
    .S(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__clkbuf_1 _2454_ (.A(_0856_),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _2455_ (.A(_0652_),
    .B(_0817_),
    .X(_0857_));
 sky130_fd_sc_hd__o22ai_1 _2456_ (.A1(_0542_),
    .A2(_0648_),
    .B1(_0857_),
    .B2(_0562_),
    .Y(_0858_));
 sky130_fd_sc_hd__nor2_1 _2457_ (.A(_0685_),
    .B(_0745_),
    .Y(_0859_));
 sky130_fd_sc_hd__a311o_1 _2458_ (.A1(_0576_),
    .A2(_0569_),
    .A3(_0799_),
    .B1(_0859_),
    .C1(\inputs.frequency_lut.rng[5] ),
    .X(_0860_));
 sky130_fd_sc_hd__a21o_1 _2459_ (.A1(_0768_),
    .A2(_0858_),
    .B1(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__nand2_1 _2460_ (.A(_0555_),
    .B(_0657_),
    .Y(_0862_));
 sky130_fd_sc_hd__o311a_1 _2461_ (.A1(_0552_),
    .A2(_0657_),
    .A3(_0656_),
    .B1(_0766_),
    .C1(_0576_),
    .X(_0863_));
 sky130_fd_sc_hd__a311o_1 _2462_ (.A1(_0768_),
    .A2(_0796_),
    .A3(_0862_),
    .B1(_0863_),
    .C1(_0578_),
    .X(_0864_));
 sky130_fd_sc_hd__or2_1 _2463_ (.A(_0229_),
    .B(_0823_),
    .X(_0865_));
 sky130_fd_sc_hd__o211a_1 _2464_ (.A1(_0247_),
    .A2(_0806_),
    .B1(_0865_),
    .C1(_0533_),
    .X(_0866_));
 sky130_fd_sc_hd__a31o_1 _2465_ (.A1(_0642_),
    .A2(_0861_),
    .A3(_0864_),
    .B1(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _2466_ (.A0(net312),
    .A1(_0867_),
    .S(_0855_),
    .X(_0868_));
 sky130_fd_sc_hd__clkbuf_1 _2467_ (.A(_0868_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2468_ (.A0(_0823_),
    .A1(_0825_),
    .S(_0230_),
    .X(_0869_));
 sky130_fd_sc_hd__a31o_1 _2469_ (.A1(_0686_),
    .A2(_0767_),
    .A3(_0862_),
    .B1(_0859_),
    .X(_0870_));
 sky130_fd_sc_hd__o211ai_1 _2470_ (.A1(_0555_),
    .A2(_0550_),
    .B1(_0810_),
    .C1(_0576_),
    .Y(_0871_));
 sky130_fd_sc_hd__a21oi_1 _2471_ (.A1(_0568_),
    .A2(_0557_),
    .B1(_0575_),
    .Y(_0872_));
 sky130_fd_sc_hd__o21ai_1 _2472_ (.A1(_0650_),
    .A2(_0745_),
    .B1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21oi_1 _2473_ (.A1(_0871_),
    .A2(_0873_),
    .B1(_0727_),
    .Y(_0874_));
 sky130_fd_sc_hd__a211o_1 _2474_ (.A1(_0727_),
    .A2(_0870_),
    .B1(_0874_),
    .C1(_0674_),
    .X(_0875_));
 sky130_fd_sc_hd__o21ai_1 _2475_ (.A1(_0642_),
    .A2(_0869_),
    .B1(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(net306),
    .A1(_0876_),
    .S(_0855_),
    .X(_0877_));
 sky130_fd_sc_hd__clkbuf_1 _2477_ (.A(_0877_),
    .X(_0126_));
 sky130_fd_sc_hd__a41o_1 _2478_ (.A1(_0551_),
    .A2(_0556_),
    .A3(_0543_),
    .A4(_0536_),
    .B1(\inputs.frequency_lut.rng[4] ),
    .X(_0878_));
 sky130_fd_sc_hd__a21oi_1 _2479_ (.A1(_0552_),
    .A2(_0657_),
    .B1(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__o21a_1 _2480_ (.A1(_0552_),
    .A2(_0537_),
    .B1(_0872_),
    .X(_0880_));
 sky130_fd_sc_hd__a21oi_1 _2481_ (.A1(_0765_),
    .A2(_0879_),
    .B1(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__a41o_1 _2482_ (.A1(_0686_),
    .A2(_0569_),
    .A3(_0537_),
    .A4(_0546_),
    .B1(_0577_),
    .X(_0882_));
 sky130_fd_sc_hd__o221a_1 _2483_ (.A1(_0727_),
    .A2(_0881_),
    .B1(_0882_),
    .B2(_0859_),
    .C1(_0603_),
    .X(_0883_));
 sky130_fd_sc_hd__a31o_1 _2484_ (.A1(_0231_),
    .A2(_0534_),
    .A3(_0830_),
    .B1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(net269),
    .A1(_0884_),
    .S(_0855_),
    .X(_0885_));
 sky130_fd_sc_hd__clkbuf_1 _2486_ (.A(_0885_),
    .X(_0127_));
 sky130_fd_sc_hd__and4_1 _2487_ (.A(\inputs.frequency_lut.rng[5] ),
    .B(_0686_),
    .C(_0569_),
    .D(_0717_),
    .X(_0886_));
 sky130_fd_sc_hd__o211a_1 _2488_ (.A1(_0656_),
    .A2(_0800_),
    .B1(_0575_),
    .C1(_0557_),
    .X(_0887_));
 sky130_fd_sc_hd__o21a_1 _2489_ (.A1(_0872_),
    .A2(_0887_),
    .B1(_0577_),
    .X(_0888_));
 sky130_fd_sc_hd__o21a_1 _2490_ (.A1(_0886_),
    .A2(_0888_),
    .B1(_0603_),
    .X(_0889_));
 sky130_fd_sc_hd__a31o_1 _2491_ (.A1(_0231_),
    .A2(_0534_),
    .A3(_0851_),
    .B1(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(net220),
    .A1(_0890_),
    .S(_0855_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_1 _2493_ (.A(_0891_),
    .X(_0128_));
 sky130_fd_sc_hd__nand2_1 _2494_ (.A(\inputs.frequency_lut.rng[5] ),
    .B(_0709_),
    .Y(_0892_));
 sky130_fd_sc_hd__a21o_1 _2495_ (.A1(_0555_),
    .A2(_0657_),
    .B1(_0878_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(\inputs.frequency_lut.rng[5] ),
    .A1(_0892_),
    .S(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__nor2_1 _2497_ (.A(_0674_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__a41o_1 _2498_ (.A1(_0231_),
    .A2(_0534_),
    .A3(_0626_),
    .A4(_0829_),
    .B1(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(net298),
    .A1(_0896_),
    .S(_0855_),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _2500_ (.A(_0897_),
    .X(_0129_));
 sky130_fd_sc_hd__or3b_1 _2501_ (.A(\inputs.octave_fsm.state[2] ),
    .B(_0823_),
    .C_N(_0228_),
    .X(_0898_));
 sky130_fd_sc_hd__or4_1 _2502_ (.A(_0727_),
    .B(_0768_),
    .C(_0533_),
    .D(_0862_),
    .X(_0899_));
 sky130_fd_sc_hd__nand2_1 _2503_ (.A(_0898_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(\outputs.div.divisor[17] ),
    .A1(_0900_),
    .S(_0855_),
    .X(_0901_));
 sky130_fd_sc_hd__clkbuf_1 _2505_ (.A(_0901_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(\outputs.divider_buffer[0] ),
    .A1(net255),
    .S(_0497_),
    .X(_0902_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(_0902_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(\outputs.divider_buffer[1] ),
    .A1(net241),
    .S(_0497_),
    .X(_0903_));
 sky130_fd_sc_hd__clkbuf_1 _2509_ (.A(_0903_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(\outputs.divider_buffer[2] ),
    .A1(net291),
    .S(_0497_),
    .X(_0904_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_0904_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_4 _2512_ (.A(_1089_),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _2513_ (.A0(\outputs.divider_buffer[3] ),
    .A1(net251),
    .S(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__clkbuf_1 _2514_ (.A(_0906_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2515_ (.A0(\outputs.divider_buffer[4] ),
    .A1(net239),
    .S(_0905_),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_1 _2516_ (.A(_0907_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(\outputs.divider_buffer[5] ),
    .A1(net257),
    .S(_0905_),
    .X(_0908_));
 sky130_fd_sc_hd__clkbuf_1 _2518_ (.A(_0908_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(\outputs.divider_buffer[6] ),
    .A1(net224),
    .S(_0905_),
    .X(_0909_));
 sky130_fd_sc_hd__clkbuf_1 _2520_ (.A(_0909_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(\outputs.divider_buffer[7] ),
    .A1(net231),
    .S(_0905_),
    .X(_0910_));
 sky130_fd_sc_hd__clkbuf_1 _2522_ (.A(_0910_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(\outputs.divider_buffer[8] ),
    .A1(net245),
    .S(_0905_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(_0911_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(\outputs.divider_buffer[9] ),
    .A1(net111),
    .S(_0905_),
    .X(_0912_));
 sky130_fd_sc_hd__clkbuf_1 _2526_ (.A(_0912_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(\outputs.divider_buffer[10] ),
    .A1(net275),
    .S(_0905_),
    .X(_0913_));
 sky130_fd_sc_hd__clkbuf_1 _2528_ (.A(_0913_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(\outputs.divider_buffer[11] ),
    .A1(net246),
    .S(_0905_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_1 _2530_ (.A(_0914_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(\outputs.divider_buffer[12] ),
    .A1(net226),
    .S(_0905_),
    .X(_0915_));
 sky130_fd_sc_hd__clkbuf_1 _2532_ (.A(_0915_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_4 _2533_ (.A(_1089_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(\outputs.divider_buffer[13] ),
    .A1(net272),
    .S(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_1 _2535_ (.A(_0917_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(\outputs.divider_buffer[14] ),
    .A1(net286),
    .S(_0916_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _2537_ (.A(net287),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\outputs.divider_buffer[15] ),
    .A1(net195),
    .S(_0916_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(_0919_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(\outputs.divider_buffer[16] ),
    .A1(net266),
    .S(_0916_),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _2541_ (.A(_0920_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(\outputs.divider_buffer[17] ),
    .A1(net248),
    .S(_0916_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(_0921_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(net237),
    .A1(net155),
    .S(_0855_),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_1 _2545_ (.A(_0922_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(net234),
    .A1(\outputs.div.oscillator_out[1] ),
    .S(_0855_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(net235),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(net188),
    .A1(net225),
    .S(_0855_),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_0924_),
    .X(_0151_));
 sky130_fd_sc_hd__buf_4 _2550_ (.A(_0512_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(net262),
    .A1(net92),
    .S(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _2552_ (.A(_0926_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(net249),
    .A1(net98),
    .S(_0925_),
    .X(_0927_));
 sky130_fd_sc_hd__clkbuf_1 _2554_ (.A(_0927_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(net215),
    .A1(net150),
    .S(_0925_),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_1 _2556_ (.A(_0928_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(net206),
    .A1(net107),
    .S(_0925_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_0929_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(net205),
    .A1(net221),
    .S(_0925_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_1 _2560_ (.A(_0930_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(net271),
    .A1(net277),
    .S(_0925_),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_1 _2562_ (.A(_0931_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(net209),
    .A1(\outputs.div.oscillator_out[9] ),
    .S(_0925_),
    .X(_0932_));
 sky130_fd_sc_hd__clkbuf_1 _2564_ (.A(_0932_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(net243),
    .A1(\outputs.div.oscillator_out[10] ),
    .S(_0925_),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_1 _2566_ (.A(net244),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(net228),
    .A1(\outputs.div.oscillator_out[11] ),
    .S(_0925_),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _2568_ (.A(net229),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(net223),
    .A1(net127),
    .S(_0925_),
    .X(_0935_));
 sky130_fd_sc_hd__clkbuf_1 _2570_ (.A(_0935_),
    .X(_0161_));
 sky130_fd_sc_hd__buf_4 _2571_ (.A(_0512_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(net232),
    .A1(\outputs.div.oscillator_out[13] ),
    .S(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__clkbuf_1 _2573_ (.A(net233),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(net254),
    .A1(net101),
    .S(_0936_),
    .X(_0938_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(_0938_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(net238),
    .A1(net103),
    .S(_0936_),
    .X(_0939_));
 sky130_fd_sc_hd__clkbuf_1 _2577_ (.A(_0939_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(net207),
    .A1(net109),
    .S(_0936_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_0940_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(net230),
    .A1(net159),
    .S(_0936_),
    .X(_0941_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(_0941_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(net155),
    .A1(\outputs.sig_gen.count[0] ),
    .S(_0936_),
    .X(_0942_));
 sky130_fd_sc_hd__clkbuf_1 _2583_ (.A(_0942_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(net300),
    .A1(\outputs.sig_gen.count[1] ),
    .S(_0936_),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_1 _2585_ (.A(_0943_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(net225),
    .A1(net294),
    .S(_0936_),
    .X(_0944_));
 sky130_fd_sc_hd__clkbuf_1 _2587_ (.A(_0944_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(net92),
    .A1(\outputs.sig_gen.count[3] ),
    .S(_0936_),
    .X(_0945_));
 sky130_fd_sc_hd__clkbuf_1 _2589_ (.A(_0945_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(net98),
    .A1(\outputs.sig_gen.count[4] ),
    .S(_0936_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_1 _2591_ (.A(_0946_),
    .X(_0171_));
 sky130_fd_sc_hd__buf_4 _2592_ (.A(_0512_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(net150),
    .A1(\outputs.sig_gen.count[5] ),
    .S(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_1 _2594_ (.A(_0948_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(net107),
    .A1(\outputs.sig_gen.count[6] ),
    .S(_0947_),
    .X(_0949_));
 sky130_fd_sc_hd__clkbuf_1 _2596_ (.A(_0949_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(net221),
    .A1(\outputs.sig_gen.count[7] ),
    .S(_0947_),
    .X(_0950_));
 sky130_fd_sc_hd__clkbuf_1 _2598_ (.A(_0950_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(net277),
    .A1(\outputs.sig_gen.count[8] ),
    .S(_0947_),
    .X(_0951_));
 sky130_fd_sc_hd__clkbuf_1 _2600_ (.A(_0951_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(\outputs.div.oscillator_out[9] ),
    .A1(\outputs.sig_gen.count[9] ),
    .S(_0947_),
    .X(_0952_));
 sky130_fd_sc_hd__clkbuf_1 _2602_ (.A(_0952_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(net309),
    .A1(\outputs.sig_gen.count[10] ),
    .S(_0947_),
    .X(_0953_));
 sky130_fd_sc_hd__clkbuf_1 _2604_ (.A(_0953_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2605_ (.A0(net304),
    .A1(\outputs.sig_gen.count[11] ),
    .S(_0947_),
    .X(_0954_));
 sky130_fd_sc_hd__clkbuf_1 _2606_ (.A(_0954_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(net127),
    .A1(\outputs.sig_gen.count[12] ),
    .S(_0947_),
    .X(_0955_));
 sky130_fd_sc_hd__clkbuf_1 _2608_ (.A(_0955_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(net302),
    .A1(\outputs.sig_gen.count[13] ),
    .S(_0947_),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(_0956_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(net101),
    .A1(\outputs.sig_gen.count[14] ),
    .S(_0947_),
    .X(_0957_));
 sky130_fd_sc_hd__clkbuf_1 _2612_ (.A(_0957_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(net103),
    .A1(\outputs.sig_gen.count[15] ),
    .S(_0512_),
    .X(_0958_));
 sky130_fd_sc_hd__clkbuf_1 _2614_ (.A(_0958_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(net109),
    .A1(\outputs.sig_gen.count[16] ),
    .S(_0512_),
    .X(_0959_));
 sky130_fd_sc_hd__clkbuf_1 _2616_ (.A(_0959_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(net159),
    .A1(net301),
    .S(_0512_),
    .X(_0960_));
 sky130_fd_sc_hd__clkbuf_1 _2618_ (.A(_0960_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(\outputs.shaper.count[0] ),
    .A1(net237),
    .S(_0916_),
    .X(_0961_));
 sky130_fd_sc_hd__clkbuf_1 _2620_ (.A(_0961_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2621_ (.A0(\outputs.shaper.count[1] ),
    .A1(net234),
    .S(_0916_),
    .X(_0962_));
 sky130_fd_sc_hd__clkbuf_1 _2622_ (.A(_0962_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2623_ (.A0(\outputs.shaper.count[2] ),
    .A1(net188),
    .S(_0916_),
    .X(_0963_));
 sky130_fd_sc_hd__clkbuf_1 _2624_ (.A(net189),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(\outputs.shaper.count[3] ),
    .A1(net262),
    .S(_0916_),
    .X(_0964_));
 sky130_fd_sc_hd__clkbuf_1 _2626_ (.A(_0964_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(\outputs.shaper.count[4] ),
    .A1(net249),
    .S(_0916_),
    .X(_0965_));
 sky130_fd_sc_hd__clkbuf_1 _2628_ (.A(_0965_),
    .X(_0189_));
 sky130_fd_sc_hd__buf_4 _2629_ (.A(_1089_),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(\outputs.shaper.count[5] ),
    .A1(net215),
    .S(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__clkbuf_1 _2631_ (.A(_0967_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(\outputs.shaper.count[6] ),
    .A1(net206),
    .S(_0966_),
    .X(_0968_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_0968_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(\outputs.shaper.count[7] ),
    .A1(net205),
    .S(_0966_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_0969_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(\outputs.shaper.count[8] ),
    .A1(net271),
    .S(_0966_),
    .X(_0970_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(_0970_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(\outputs.shaper.count[9] ),
    .A1(net209),
    .S(_0966_),
    .X(_0971_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(_0971_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(net282),
    .A1(net243),
    .S(_0966_),
    .X(_0972_));
 sky130_fd_sc_hd__clkbuf_1 _2641_ (.A(_0972_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(net259),
    .A1(net228),
    .S(_0966_),
    .X(_0973_));
 sky130_fd_sc_hd__clkbuf_1 _2643_ (.A(_0973_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(\outputs.shaper.count[12] ),
    .A1(net223),
    .S(_0966_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_1 _2645_ (.A(_0974_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(\outputs.shaper.count[13] ),
    .A1(net232),
    .S(_0966_),
    .X(_0975_));
 sky130_fd_sc_hd__clkbuf_1 _2647_ (.A(_0975_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(net273),
    .A1(net254),
    .S(_0966_),
    .X(_0976_));
 sky130_fd_sc_hd__clkbuf_1 _2649_ (.A(_0976_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(\outputs.shaper.count[15] ),
    .A1(net238),
    .S(_1089_),
    .X(_0977_));
 sky130_fd_sc_hd__clkbuf_1 _2651_ (.A(_0977_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(\outputs.shaper.count[16] ),
    .A1(net207),
    .S(_1089_),
    .X(_0978_));
 sky130_fd_sc_hd__clkbuf_1 _2653_ (.A(_0978_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2654_ (.A0(\outputs.shaper.count[17] ),
    .A1(net230),
    .S(_1089_),
    .X(_0979_));
 sky130_fd_sc_hd__clkbuf_1 _2655_ (.A(_0979_),
    .X(_0202_));
 sky130_fd_sc_hd__xnor2_1 _2656_ (.A(_0727_),
    .B(_0768_),
    .Y(_0980_));
 sky130_fd_sc_hd__xnor2_1 _2657_ (.A(_0562_),
    .B(_1182_),
    .Y(_0981_));
 sky130_fd_sc_hd__xnor2_1 _2658_ (.A(_0980_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_4 _2659_ (.A(_1039_),
    .B(_0642_),
    .Y(_0983_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(_0982_),
    .A1(_0556_),
    .S(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_1 _2661_ (.A(_0984_),
    .X(_0203_));
 sky130_fd_sc_hd__xor2_1 _2662_ (.A(_0556_),
    .B(_1182_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(_0985_),
    .A1(_0543_),
    .S(_0983_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_1 _2664_ (.A(_0986_),
    .X(_0204_));
 sky130_fd_sc_hd__xor2_1 _2665_ (.A(_0543_),
    .B(_1182_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(_0987_),
    .A1(_0537_),
    .S(_0983_),
    .X(_0988_));
 sky130_fd_sc_hd__clkbuf_1 _2667_ (.A(_0988_),
    .X(_0205_));
 sky130_fd_sc_hd__xor2_1 _2668_ (.A(_0537_),
    .B(_1182_),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _2669_ (.A0(_0989_),
    .A1(_0562_),
    .S(_0983_),
    .X(_0990_));
 sky130_fd_sc_hd__clkbuf_1 _2670_ (.A(_0990_),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _2671_ (.A(_0768_),
    .B(_0983_),
    .Y(_0991_));
 sky130_fd_sc_hd__o21ai_1 _2672_ (.A1(_0983_),
    .A2(_0981_),
    .B1(_0991_),
    .Y(_0207_));
 sky130_fd_sc_hd__xor2_1 _2673_ (.A(_0768_),
    .B(_1182_),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(_0992_),
    .A1(_0727_),
    .S(_0983_),
    .X(_0993_));
 sky130_fd_sc_hd__clkbuf_1 _2675_ (.A(_0993_),
    .X(_0208_));
 sky130_fd_sc_hd__dfrtp_1 _2676_ (.CLK(clknet_leaf_16_clk),
    .D(\outputs.sample_rate.next_count[0] ),
    .RESET_B(net51),
    .Q(\outputs.sample_rate.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2677_ (.CLK(clknet_leaf_17_clk),
    .D(\outputs.sample_rate.next_count[1] ),
    .RESET_B(net51),
    .Q(\outputs.sample_rate.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2678_ (.CLK(clknet_leaf_16_clk),
    .D(\outputs.sample_rate.next_count[2] ),
    .RESET_B(net51),
    .Q(\outputs.sample_rate.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2679_ (.CLK(clknet_leaf_16_clk),
    .D(\outputs.sample_rate.next_count[3] ),
    .RESET_B(net51),
    .Q(\outputs.sample_rate.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2680_ (.CLK(clknet_leaf_9_clk),
    .D(net142),
    .RESET_B(net43),
    .Q(\outputs.sample_rate.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2681_ (.CLK(clknet_leaf_9_clk),
    .D(\outputs.sample_rate.next_count[5] ),
    .RESET_B(net43),
    .Q(\outputs.sample_rate.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2682_ (.CLK(clknet_leaf_9_clk),
    .D(\outputs.sample_rate.next_count[6] ),
    .RESET_B(net43),
    .Q(\outputs.sample_rate.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2683_ (.CLK(clknet_leaf_9_clk),
    .D(\outputs.sample_rate.next_count[7] ),
    .RESET_B(net55),
    .Q(\outputs.sample_rate.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2684_ (.CLK(clknet_leaf_26_clk),
    .D(\inputs.wavetype_fsm.next_state[0] ),
    .RESET_B(net35),
    .Q(\inputs.wavetype_fsm.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2685_ (.CLK(clknet_leaf_26_clk),
    .D(net184),
    .RESET_B(net35),
    .Q(\inputs.wavetype_fsm.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2686_ (.CLK(clknet_leaf_23_clk),
    .D(_0000_),
    .RESET_B(net32),
    .Q(\outputs.div.m[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2687_ (.CLK(clknet_leaf_34_clk),
    .D(_0001_),
    .RESET_B(net33),
    .Q(\outputs.div.m[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2688_ (.CLK(clknet_leaf_34_clk),
    .D(_0002_),
    .RESET_B(net33),
    .Q(\outputs.div.m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2689_ (.CLK(clknet_leaf_23_clk),
    .D(_0003_),
    .RESET_B(net33),
    .Q(\outputs.div.m[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2690_ (.CLK(clknet_leaf_34_clk),
    .D(_0004_),
    .RESET_B(net32),
    .Q(\outputs.div.m[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2691_ (.CLK(clknet_leaf_34_clk),
    .D(_0005_),
    .RESET_B(net32),
    .Q(\outputs.div.m[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2692_ (.CLK(clknet_leaf_34_clk),
    .D(_0006_),
    .RESET_B(net33),
    .Q(\outputs.div.m[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2693_ (.CLK(clknet_leaf_34_clk),
    .D(_0007_),
    .RESET_B(net33),
    .Q(\outputs.div.m[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2694_ (.CLK(clknet_leaf_23_clk),
    .D(_0008_),
    .RESET_B(net45),
    .Q(\outputs.div.m[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2695_ (.CLK(clknet_leaf_13_clk),
    .D(_0009_),
    .RESET_B(net45),
    .Q(\outputs.div.m[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2696_ (.CLK(clknet_leaf_23_clk),
    .D(_0010_),
    .RESET_B(net45),
    .Q(\outputs.div.m[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2697_ (.CLK(clknet_leaf_13_clk),
    .D(_0011_),
    .RESET_B(net45),
    .Q(\outputs.div.m[11] ));
 sky130_fd_sc_hd__dfrtp_2 _2698_ (.CLK(clknet_leaf_23_clk),
    .D(_0012_),
    .RESET_B(net45),
    .Q(\outputs.div.m[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2699_ (.CLK(clknet_leaf_13_clk),
    .D(_0013_),
    .RESET_B(net45),
    .Q(\outputs.div.m[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2700_ (.CLK(clknet_leaf_13_clk),
    .D(_0014_),
    .RESET_B(net45),
    .Q(\outputs.div.m[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2701_ (.CLK(clknet_leaf_14_clk),
    .D(_0015_),
    .RESET_B(net45),
    .Q(\outputs.div.m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2702_ (.CLK(clknet_leaf_14_clk),
    .D(_0016_),
    .RESET_B(net46),
    .Q(\outputs.div.m[16] ));
 sky130_fd_sc_hd__dfrtp_2 _2703_ (.CLK(clknet_leaf_14_clk),
    .D(_0017_),
    .RESET_B(net46),
    .Q(\outputs.div.m[17] ));
 sky130_fd_sc_hd__dfstp_1 _2704_ (.CLK(clknet_leaf_37_clk),
    .D(\inputs.random_note_generator.feedback ),
    .SET_B(net22),
    .Q(\inputs.random_note_generator.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2705_ (.CLK(clknet_leaf_37_clk),
    .D(net82),
    .RESET_B(net22),
    .Q(\inputs.random_note_generator.out[1] ));
 sky130_fd_sc_hd__dfstp_1 _2706_ (.CLK(clknet_leaf_37_clk),
    .D(net76),
    .SET_B(net22),
    .Q(\inputs.random_note_generator.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2707_ (.CLK(clknet_leaf_37_clk),
    .D(net84),
    .RESET_B(net22),
    .Q(\inputs.random_note_generator.out[3] ));
 sky130_fd_sc_hd__dfstp_1 _2708_ (.CLK(clknet_leaf_37_clk),
    .D(net73),
    .SET_B(net22),
    .Q(\inputs.random_note_generator.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2709_ (.CLK(clknet_leaf_37_clk),
    .D(net83),
    .RESET_B(net22),
    .Q(\inputs.random_note_generator.out[5] ));
 sky130_fd_sc_hd__dfstp_1 _2710_ (.CLK(clknet_leaf_37_clk),
    .D(net70),
    .SET_B(net22),
    .Q(\inputs.random_note_generator.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2711_ (.CLK(clknet_leaf_37_clk),
    .D(net81),
    .RESET_B(net22),
    .Q(\inputs.random_note_generator.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2712_ (.CLK(clknet_leaf_37_clk),
    .D(net71),
    .RESET_B(net23),
    .Q(\inputs.random_note_generator.out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2713_ (.CLK(clknet_leaf_37_clk),
    .D(net68),
    .RESET_B(net23),
    .Q(\inputs.random_note_generator.out[9] ));
 sky130_fd_sc_hd__dfstp_1 _2714_ (.CLK(clknet_leaf_37_clk),
    .D(net75),
    .SET_B(net23),
    .Q(\inputs.random_note_generator.out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2715_ (.CLK(clknet_leaf_37_clk),
    .D(net89),
    .RESET_B(net22),
    .Q(\inputs.random_note_generator.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2716_ (.CLK(clknet_leaf_37_clk),
    .D(net67),
    .RESET_B(net22),
    .Q(\inputs.random_note_generator.out[12] ));
 sky130_fd_sc_hd__dfstp_1 _2717_ (.CLK(clknet_leaf_37_clk),
    .D(net85),
    .SET_B(net23),
    .Q(\inputs.random_note_generator.out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2718_ (.CLK(clknet_leaf_37_clk),
    .D(net87),
    .RESET_B(net23),
    .Q(\inputs.random_note_generator.out[14] ));
 sky130_fd_sc_hd__dfstp_1 _2719_ (.CLK(clknet_leaf_37_clk),
    .D(net72),
    .SET_B(net23),
    .Q(\inputs.random_note_generator.out[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2720_ (.CLK(clknet_leaf_32_clk),
    .D(_0018_),
    .RESET_B(net27),
    .Q(\inputs.octave_fsm.state[0] ));
 sky130_fd_sc_hd__dfstp_2 _2721_ (.CLK(clknet_leaf_35_clk),
    .D(_0019_),
    .SET_B(net24),
    .Q(\inputs.octave_fsm.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2722_ (.CLK(clknet_leaf_32_clk),
    .D(_0020_),
    .RESET_B(net27),
    .Q(\inputs.octave_fsm.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _2723_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.random_update_clock.next_count[0] ),
    .SET_B(net27),
    .Q(\inputs.random_update_clock.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2724_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.random_update_clock.next_count[1] ),
    .RESET_B(net27),
    .Q(\inputs.random_update_clock.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2725_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.random_update_clock.next_count[2] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2726_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.random_update_clock.next_count[3] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2727_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[4] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2728_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[5] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2729_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[6] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2730_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[7] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2731_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[8] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2732_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[9] ),
    .RESET_B(net30),
    .Q(\inputs.random_update_clock.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2733_ (.CLK(clknet_leaf_29_clk),
    .D(\inputs.random_update_clock.next_count[10] ),
    .RESET_B(net30),
    .Q(\inputs.random_update_clock.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2734_ (.CLK(clknet_leaf_29_clk),
    .D(\inputs.random_update_clock.next_count[11] ),
    .RESET_B(net30),
    .Q(\inputs.random_update_clock.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2735_ (.CLK(clknet_leaf_29_clk),
    .D(\inputs.random_update_clock.next_count[12] ),
    .RESET_B(net30),
    .Q(\inputs.random_update_clock.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2736_ (.CLK(clknet_leaf_29_clk),
    .D(\inputs.random_update_clock.next_count[13] ),
    .RESET_B(net31),
    .Q(\inputs.random_update_clock.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2737_ (.CLK(clknet_leaf_29_clk),
    .D(\inputs.random_update_clock.next_count[14] ),
    .RESET_B(net30),
    .Q(\inputs.random_update_clock.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2738_ (.CLK(clknet_leaf_29_clk),
    .D(\inputs.random_update_clock.next_count[15] ),
    .RESET_B(net30),
    .Q(\inputs.random_update_clock.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2739_ (.CLK(clknet_leaf_31_clk),
    .D(\inputs.random_update_clock.next_count[16] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2740_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[17] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2741_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.random_update_clock.next_count[18] ),
    .RESET_B(net29),
    .Q(\inputs.random_update_clock.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2742_ (.CLK(clknet_leaf_31_clk),
    .D(\inputs.random_update_clock.next_count[19] ),
    .RESET_B(net31),
    .Q(\inputs.random_update_clock.count[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2743_ (.CLK(clknet_leaf_31_clk),
    .D(\inputs.random_update_clock.next_count[20] ),
    .RESET_B(net31),
    .Q(\inputs.random_update_clock.count[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2744_ (.CLK(clknet_leaf_28_clk),
    .D(\inputs.random_update_clock.next_count[21] ),
    .RESET_B(net31),
    .Q(\inputs.random_update_clock.count[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2745_ (.CLK(clknet_leaf_29_clk),
    .D(net97),
    .RESET_B(net31),
    .Q(\inputs.random_update_clock.count[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2746_ (.CLK(clknet_leaf_25_clk),
    .D(net95),
    .RESET_B(net34),
    .Q(\inputs.mode_edge.ff_out ));
 sky130_fd_sc_hd__dfrtp_1 _2747_ (.CLK(clknet_leaf_25_clk),
    .D(\inputs.mode_edge.ff_in ),
    .RESET_B(net34),
    .Q(\inputs.mode_edge.det_edge ));
 sky130_fd_sc_hd__dfrtp_1 _2748_ (.CLK(clknet_leaf_31_clk),
    .D(\inputs.down.in ),
    .RESET_B(net31),
    .Q(\inputs.down.ff_out ));
 sky130_fd_sc_hd__dfrtp_1 _2749_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.down.ff_in ),
    .RESET_B(net27),
    .Q(\inputs.down.det_edge ));
 sky130_fd_sc_hd__dfrtp_1 _2750_ (.CLK(clknet_leaf_31_clk),
    .D(net88),
    .RESET_B(net31),
    .Q(\inputs.up.ff_out ));
 sky130_fd_sc_hd__dfrtp_1 _2751_ (.CLK(clknet_leaf_30_clk),
    .D(\inputs.up.ff_in ),
    .RESET_B(net27),
    .Q(\inputs.octave_fsm.octave_key_up ));
 sky130_fd_sc_hd__dfrtp_1 _2752_ (.CLK(clknet_leaf_28_clk),
    .D(net58),
    .RESET_B(net34),
    .Q(\inputs.key_encoder.sync_keys[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2753_ (.CLK(clknet_leaf_32_clk),
    .D(net66),
    .RESET_B(net27),
    .Q(\inputs.key_encoder.sync_keys[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2754_ (.CLK(clknet_leaf_32_clk),
    .D(net69),
    .RESET_B(net28),
    .Q(\inputs.key_encoder.sync_keys[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2755_ (.CLK(clknet_leaf_32_clk),
    .D(net65),
    .RESET_B(net28),
    .Q(\inputs.key_encoder.sync_keys[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2756_ (.CLK(clknet_leaf_33_clk),
    .D(net61),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2757_ (.CLK(clknet_leaf_28_clk),
    .D(net57),
    .RESET_B(net34),
    .Q(\inputs.key_encoder.sync_keys[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2758_ (.CLK(clknet_leaf_33_clk),
    .D(net79),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2759_ (.CLK(clknet_leaf_25_clk),
    .D(net56),
    .RESET_B(net34),
    .Q(\inputs.key_encoder.sync_keys[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2760_ (.CLK(clknet_leaf_32_clk),
    .D(net64),
    .RESET_B(net28),
    .Q(\inputs.key_encoder.sync_keys[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2761_ (.CLK(clknet_leaf_0_clk),
    .D(net63),
    .RESET_B(net25),
    .Q(\inputs.key_encoder.sync_keys[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2762_ (.CLK(clknet_leaf_33_clk),
    .D(net86),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2763_ (.CLK(clknet_leaf_38_clk),
    .D(net59),
    .RESET_B(net25),
    .Q(\inputs.key_encoder.sync_keys[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2764_ (.CLK(clknet_leaf_38_clk),
    .D(net60),
    .RESET_B(net25),
    .Q(\inputs.key_encoder.sync_keys[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2765_ (.CLK(clknet_leaf_35_clk),
    .D(net78),
    .RESET_B(net28),
    .Q(\inputs.key_encoder.sync_keys[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2766_ (.CLK(clknet_leaf_28_clk),
    .D(net77),
    .RESET_B(net31),
    .Q(\inputs.key_encoder.sync_keys[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2767_ (.CLK(clknet_leaf_33_clk),
    .D(net80),
    .RESET_B(net34),
    .Q(\inputs.key_encoder.sync_keys[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2768_ (.CLK(clknet_leaf_28_clk),
    .D(net74),
    .RESET_B(net36),
    .Q(\inputs.key_encoder.octave_key_up ));
 sky130_fd_sc_hd__dfrtp_1 _2769_ (.CLK(clknet_leaf_25_clk),
    .D(\inputs.keypad[0] ),
    .RESET_B(net34),
    .Q(\inputs.keypad_synchronizer.half_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2770_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.keypad[1] ),
    .RESET_B(net27),
    .Q(\inputs.keypad_synchronizer.half_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2771_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.keypad[2] ),
    .RESET_B(net28),
    .Q(\inputs.keypad_synchronizer.half_sync[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2772_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.keypad[3] ),
    .RESET_B(net27),
    .Q(\inputs.keypad_synchronizer.half_sync[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2773_ (.CLK(clknet_leaf_33_clk),
    .D(\inputs.keypad[4] ),
    .RESET_B(net32),
    .Q(\inputs.keypad_synchronizer.half_sync[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2774_ (.CLK(clknet_leaf_25_clk),
    .D(\inputs.keypad[5] ),
    .RESET_B(net34),
    .Q(\inputs.keypad_synchronizer.half_sync[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2775_ (.CLK(clknet_leaf_0_clk),
    .D(\inputs.keypad[6] ),
    .RESET_B(net25),
    .Q(\inputs.keypad_synchronizer.half_sync[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2776_ (.CLK(clknet_leaf_24_clk),
    .D(\inputs.keypad[7] ),
    .RESET_B(net32),
    .Q(\inputs.keypad_synchronizer.half_sync[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2777_ (.CLK(clknet_leaf_32_clk),
    .D(\inputs.keypad[8] ),
    .RESET_B(net27),
    .Q(\inputs.keypad_synchronizer.half_sync[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2778_ (.CLK(clknet_leaf_0_clk),
    .D(\inputs.keypad[9] ),
    .RESET_B(net25),
    .Q(\inputs.keypad_synchronizer.half_sync[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2779_ (.CLK(clknet_leaf_16_clk),
    .D(\inputs.keypad[10] ),
    .RESET_B(net51),
    .Q(\inputs.keypad_synchronizer.half_sync[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2780_ (.CLK(clknet_leaf_38_clk),
    .D(\inputs.keypad[11] ),
    .RESET_B(net25),
    .Q(\inputs.keypad_synchronizer.half_sync[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2781_ (.CLK(clknet_leaf_38_clk),
    .D(\inputs.keypad[12] ),
    .RESET_B(net25),
    .Q(\inputs.keypad_synchronizer.half_sync[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2782_ (.CLK(clknet_leaf_38_clk),
    .D(\inputs.keypad[13] ),
    .RESET_B(net24),
    .Q(\inputs.keypad_synchronizer.half_sync[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2783_ (.CLK(clknet_leaf_28_clk),
    .D(\inputs.keypad[14] ),
    .RESET_B(net36),
    .Q(\inputs.keypad_synchronizer.half_sync[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2784_ (.CLK(clknet_leaf_38_clk),
    .D(\inputs.keypad[15] ),
    .RESET_B(net25),
    .Q(\inputs.keypad_synchronizer.half_sync[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2785_ (.CLK(clknet_leaf_28_clk),
    .D(\inputs.keypad[16] ),
    .RESET_B(net34),
    .Q(\inputs.keypad_synchronizer.half_sync[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2786_ (.CLK(clknet_leaf_28_clk),
    .D(\outputs.output_gen.pwm_unff ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.pwm_ff ));
 sky130_fd_sc_hd__dfrtp_1 _2787_ (.CLK(clknet_leaf_23_clk),
    .D(_0021_),
    .RESET_B(net33),
    .Q(\outputs.div.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2788_ (.CLK(clknet_leaf_24_clk),
    .D(_0022_),
    .RESET_B(net33),
    .Q(\outputs.div.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2789_ (.CLK(clknet_leaf_26_clk),
    .D(_0023_),
    .RESET_B(net35),
    .Q(\outputs.div.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2790_ (.CLK(clknet_leaf_26_clk),
    .D(_0024_),
    .RESET_B(net35),
    .Q(\outputs.div.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2791_ (.CLK(clknet_leaf_25_clk),
    .D(_0025_),
    .RESET_B(net34),
    .Q(\outputs.div.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2792_ (.CLK(clknet_leaf_25_clk),
    .D(_0026_),
    .RESET_B(net32),
    .Q(\outputs.div.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2793_ (.CLK(clknet_leaf_24_clk),
    .D(_0027_),
    .RESET_B(net32),
    .Q(\outputs.div.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2794_ (.CLK(clknet_leaf_25_clk),
    .D(_0028_),
    .RESET_B(net33),
    .Q(\outputs.div.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2795_ (.CLK(clknet_leaf_23_clk),
    .D(_0029_),
    .RESET_B(net45),
    .Q(\outputs.div.a[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2796_ (.CLK(clknet_leaf_22_clk),
    .D(_0030_),
    .RESET_B(net49),
    .Q(\outputs.div.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2797_ (.CLK(clknet_leaf_21_clk),
    .D(_0031_),
    .RESET_B(net49),
    .Q(\outputs.div.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2798_ (.CLK(clknet_leaf_22_clk),
    .D(_0032_),
    .RESET_B(net47),
    .Q(\outputs.div.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2799_ (.CLK(clknet_leaf_22_clk),
    .D(_0033_),
    .RESET_B(net45),
    .Q(\outputs.div.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2800_ (.CLK(clknet_leaf_22_clk),
    .D(_0034_),
    .RESET_B(net47),
    .Q(\outputs.div.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2801_ (.CLK(clknet_leaf_14_clk),
    .D(_0035_),
    .RESET_B(net46),
    .Q(\outputs.div.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2802_ (.CLK(clknet_leaf_20_clk),
    .D(_0036_),
    .RESET_B(net47),
    .Q(\outputs.div.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2803_ (.CLK(clknet_leaf_15_clk),
    .D(_0037_),
    .RESET_B(net50),
    .Q(\outputs.div.a[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2804_ (.CLK(clknet_leaf_18_clk),
    .D(_0038_),
    .RESET_B(net52),
    .Q(\outputs.div.a[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2805_ (.CLK(clknet_leaf_18_clk),
    .D(_0039_),
    .RESET_B(net53),
    .Q(\outputs.div.a[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2806_ (.CLK(clknet_leaf_18_clk),
    .D(_0040_),
    .RESET_B(net53),
    .Q(\outputs.div.a[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2807_ (.CLK(clknet_leaf_17_clk),
    .D(_0041_),
    .RESET_B(net53),
    .Q(\outputs.div.a[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2808_ (.CLK(clknet_leaf_17_clk),
    .D(_0042_),
    .RESET_B(net51),
    .Q(\outputs.div.a[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2809_ (.CLK(clknet_leaf_17_clk),
    .D(_0043_),
    .RESET_B(net51),
    .Q(\outputs.div.a[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2810_ (.CLK(clknet_leaf_16_clk),
    .D(_0044_),
    .RESET_B(net54),
    .Q(\outputs.div.a[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2811_ (.CLK(clknet_leaf_15_clk),
    .D(_0045_),
    .RESET_B(net50),
    .Q(\outputs.div.a[24] ));
 sky130_fd_sc_hd__dfrtp_2 _2812_ (.CLK(clknet_leaf_15_clk),
    .D(_0046_),
    .RESET_B(net50),
    .Q(\outputs.div.a[25] ));
 sky130_fd_sc_hd__dfrtp_1 _2813_ (.CLK(clknet_leaf_18_clk),
    .D(_0047_),
    .RESET_B(net52),
    .Q(\outputs.div.q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2814_ (.CLK(clknet_leaf_18_clk),
    .D(_0048_),
    .RESET_B(net52),
    .Q(\outputs.div.q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2815_ (.CLK(clknet_leaf_19_clk),
    .D(net214),
    .RESET_B(net52),
    .Q(\outputs.div.q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2816_ (.CLK(clknet_leaf_19_clk),
    .D(_0050_),
    .RESET_B(net52),
    .Q(\outputs.div.q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2817_ (.CLK(clknet_leaf_18_clk),
    .D(_0051_),
    .RESET_B(net52),
    .Q(\outputs.div.q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2818_ (.CLK(clknet_leaf_19_clk),
    .D(_0052_),
    .RESET_B(net52),
    .Q(\outputs.div.q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2819_ (.CLK(clknet_leaf_19_clk),
    .D(_0053_),
    .RESET_B(net52),
    .Q(\outputs.div.q[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2820_ (.CLK(clknet_leaf_20_clk),
    .D(net200),
    .RESET_B(net52),
    .Q(\outputs.div.q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2821_ (.CLK(clknet_leaf_15_clk),
    .D(net156),
    .RESET_B(net50),
    .Q(\outputs.div.q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2822_ (.CLK(clknet_leaf_10_clk),
    .D(net137),
    .RESET_B(net50),
    .Q(\outputs.div.q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2823_ (.CLK(clknet_leaf_10_clk),
    .D(net121),
    .RESET_B(net44),
    .Q(\outputs.div.q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2824_ (.CLK(clknet_leaf_9_clk),
    .D(net93),
    .RESET_B(net44),
    .Q(\outputs.div.q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2825_ (.CLK(clknet_leaf_9_clk),
    .D(net99),
    .RESET_B(net43),
    .Q(\outputs.div.q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2826_ (.CLK(clknet_leaf_7_clk),
    .D(net151),
    .RESET_B(net41),
    .Q(\outputs.div.q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2827_ (.CLK(clknet_leaf_6_clk),
    .D(net108),
    .RESET_B(net41),
    .Q(\outputs.div.q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2828_ (.CLK(clknet_leaf_6_clk),
    .D(net117),
    .RESET_B(net41),
    .Q(\outputs.div.q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2829_ (.CLK(clknet_leaf_6_clk),
    .D(net125),
    .RESET_B(net41),
    .Q(\outputs.div.q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2830_ (.CLK(clknet_leaf_6_clk),
    .D(net135),
    .RESET_B(net41),
    .Q(\outputs.div.q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2831_ (.CLK(clknet_leaf_6_clk),
    .D(net147),
    .RESET_B(net41),
    .Q(\outputs.div.q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2832_ (.CLK(clknet_leaf_6_clk),
    .D(net119),
    .RESET_B(net41),
    .Q(\outputs.div.q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2833_ (.CLK(clknet_leaf_7_clk),
    .D(net128),
    .RESET_B(net41),
    .Q(\outputs.div.q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2834_ (.CLK(clknet_leaf_7_clk),
    .D(net153),
    .RESET_B(net41),
    .Q(\outputs.div.q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2835_ (.CLK(clknet_leaf_8_clk),
    .D(net102),
    .RESET_B(net41),
    .Q(\outputs.div.q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2836_ (.CLK(clknet_leaf_8_clk),
    .D(net104),
    .RESET_B(net43),
    .Q(\outputs.div.q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2837_ (.CLK(clknet_leaf_9_clk),
    .D(net110),
    .RESET_B(net43),
    .Q(\outputs.div.q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _2838_ (.CLK(clknet_leaf_9_clk),
    .D(net160),
    .RESET_B(net44),
    .Q(\outputs.div.q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _2839_ (.CLK(clknet_leaf_15_clk),
    .D(net265),
    .RESET_B(net50),
    .Q(\outputs.div.q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _2840_ (.CLK(clknet_leaf_16_clk),
    .D(_0074_),
    .RESET_B(net51),
    .Q(\outputs.div.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2841_ (.CLK(clknet_leaf_16_clk),
    .D(_0075_),
    .RESET_B(net51),
    .Q(\outputs.div.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2842_ (.CLK(clknet_leaf_16_clk),
    .D(_0076_),
    .RESET_B(net51),
    .Q(\outputs.div.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2843_ (.CLK(clknet_leaf_16_clk),
    .D(_0077_),
    .RESET_B(net50),
    .Q(\outputs.div.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2844_ (.CLK(clknet_leaf_16_clk),
    .D(_0078_),
    .RESET_B(net50),
    .Q(\outputs.div.count[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2845_ (.CLK(clknet_leaf_22_clk),
    .D(_0079_),
    .RESET_B(net47),
    .Q(\outputs.scaled_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2846_ (.CLK(clknet_leaf_20_clk),
    .D(_0080_),
    .RESET_B(net47),
    .Q(\outputs.scaled_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2847_ (.CLK(clknet_leaf_21_clk),
    .D(_0081_),
    .RESET_B(net48),
    .Q(\outputs.scaled_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2848_ (.CLK(clknet_leaf_20_clk),
    .D(_0082_),
    .RESET_B(net48),
    .Q(\outputs.scaled_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2849_ (.CLK(clknet_leaf_20_clk),
    .D(_0083_),
    .RESET_B(net48),
    .Q(\outputs.scaled_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2850_ (.CLK(clknet_leaf_20_clk),
    .D(_0084_),
    .RESET_B(net48),
    .Q(\outputs.scaled_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2851_ (.CLK(clknet_leaf_20_clk),
    .D(_0085_),
    .RESET_B(net47),
    .Q(\outputs.scaled_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2852_ (.CLK(clknet_leaf_22_clk),
    .D(_0086_),
    .RESET_B(net47),
    .Q(\outputs.scaled_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2853_ (.CLK(clknet_leaf_22_clk),
    .D(net130),
    .RESET_B(net47),
    .Q(\outputs.div.q_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2854_ (.CLK(clknet_leaf_19_clk),
    .D(net106),
    .RESET_B(net52),
    .Q(\outputs.div.q_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2855_ (.CLK(clknet_leaf_19_clk),
    .D(net202),
    .RESET_B(net53),
    .Q(\outputs.div.q_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2856_ (.CLK(clknet_leaf_19_clk),
    .D(net164),
    .RESET_B(net53),
    .Q(\outputs.div.q_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2857_ (.CLK(clknet_leaf_19_clk),
    .D(net123),
    .RESET_B(net53),
    .Q(\outputs.div.q_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2858_ (.CLK(clknet_leaf_20_clk),
    .D(net144),
    .RESET_B(net48),
    .Q(\outputs.div.q_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2859_ (.CLK(clknet_leaf_20_clk),
    .D(net139),
    .RESET_B(net47),
    .Q(\outputs.div.q_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2860_ (.CLK(clknet_leaf_20_clk),
    .D(net172),
    .RESET_B(net47),
    .Q(\outputs.div.q_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2861_ (.CLK(clknet_leaf_17_clk),
    .D(\outputs.div.next_div ),
    .RESET_B(net54),
    .Q(\outputs.div.div ));
 sky130_fd_sc_hd__dfrtp_1 _2862_ (.CLK(clknet_leaf_15_clk),
    .D(\outputs.div.next_start ),
    .RESET_B(net50),
    .Q(\outputs.div.start ));
 sky130_fd_sc_hd__dfrtp_1 _2863_ (.CLK(clknet_leaf_27_clk),
    .D(\outputs.output_gen.next_count[0] ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2864_ (.CLK(clknet_leaf_21_clk),
    .D(net91),
    .RESET_B(net49),
    .Q(\outputs.output_gen.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2865_ (.CLK(clknet_leaf_27_clk),
    .D(\outputs.output_gen.next_count[2] ),
    .RESET_B(net49),
    .Q(\outputs.output_gen.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2866_ (.CLK(clknet_leaf_26_clk),
    .D(\outputs.output_gen.next_count[3] ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2867_ (.CLK(clknet_leaf_26_clk),
    .D(\outputs.output_gen.next_count[4] ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2868_ (.CLK(clknet_leaf_26_clk),
    .D(\outputs.output_gen.next_count[5] ),
    .RESET_B(net36),
    .Q(\outputs.output_gen.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2869_ (.CLK(clknet_leaf_26_clk),
    .D(\outputs.output_gen.next_count[6] ),
    .RESET_B(net49),
    .Q(\outputs.output_gen.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2870_ (.CLK(clknet_leaf_22_clk),
    .D(net149),
    .RESET_B(net49),
    .Q(\outputs.output_gen.count[7] ));
 sky130_fd_sc_hd__dfstp_2 _2871_ (.CLK(clknet_leaf_1_clk),
    .D(\outputs.sig_gen.next_count[0] ),
    .SET_B(net38),
    .Q(\outputs.sig_gen.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2872_ (.CLK(clknet_leaf_12_clk),
    .D(\outputs.sig_gen.next_count[1] ),
    .RESET_B(net38),
    .Q(\outputs.sig_gen.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2873_ (.CLK(clknet_leaf_11_clk),
    .D(\outputs.sig_gen.next_count[2] ),
    .RESET_B(net38),
    .Q(\outputs.sig_gen.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2874_ (.CLK(clknet_leaf_2_clk),
    .D(\outputs.sig_gen.next_count[3] ),
    .RESET_B(net38),
    .Q(\outputs.sig_gen.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2875_ (.CLK(clknet_leaf_2_clk),
    .D(\outputs.sig_gen.next_count[4] ),
    .RESET_B(net38),
    .Q(\outputs.sig_gen.count[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2876_ (.CLK(clknet_leaf_2_clk),
    .D(\outputs.sig_gen.next_count[5] ),
    .RESET_B(net38),
    .Q(\outputs.sig_gen.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2877_ (.CLK(clknet_leaf_2_clk),
    .D(\outputs.sig_gen.next_count[6] ),
    .RESET_B(net37),
    .Q(\outputs.sig_gen.count[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2878_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[7] ),
    .RESET_B(net37),
    .Q(\outputs.sig_gen.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2879_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[8] ),
    .RESET_B(net37),
    .Q(\outputs.sig_gen.count[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2880_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[9] ),
    .RESET_B(net37),
    .Q(\outputs.sig_gen.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2881_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[10] ),
    .RESET_B(net37),
    .Q(\outputs.sig_gen.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2882_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[11] ),
    .RESET_B(net37),
    .Q(\outputs.sig_gen.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2883_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[12] ),
    .RESET_B(net42),
    .Q(\outputs.sig_gen.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2884_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[13] ),
    .RESET_B(net42),
    .Q(\outputs.sig_gen.count[13] ));
 sky130_fd_sc_hd__dfrtp_2 _2885_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[14] ),
    .RESET_B(net42),
    .Q(\outputs.sig_gen.count[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2886_ (.CLK(clknet_leaf_8_clk),
    .D(\outputs.sig_gen.next_count[15] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2887_ (.CLK(clknet_leaf_8_clk),
    .D(\outputs.sig_gen.next_count[16] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2888_ (.CLK(clknet_leaf_11_clk),
    .D(\outputs.sig_gen.next_count[17] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2889_ (.CLK(clknet_leaf_1_clk),
    .D(_0095_),
    .Q(\outputs.divider_buffer2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2890_ (.CLK(clknet_leaf_1_clk),
    .D(_0096_),
    .Q(\outputs.divider_buffer2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2891_ (.CLK(clknet_leaf_1_clk),
    .D(_0097_),
    .Q(\outputs.divider_buffer2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2892_ (.CLK(clknet_leaf_1_clk),
    .D(_0098_),
    .Q(\outputs.divider_buffer2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2893_ (.CLK(clknet_leaf_0_clk),
    .D(_0099_),
    .Q(\outputs.divider_buffer2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2894_ (.CLK(clknet_leaf_0_clk),
    .D(_0100_),
    .Q(\outputs.divider_buffer2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2895_ (.CLK(clknet_leaf_0_clk),
    .D(_0101_),
    .Q(\outputs.divider_buffer2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2896_ (.CLK(clknet_leaf_0_clk),
    .D(_0102_),
    .Q(\outputs.divider_buffer2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2897_ (.CLK(clknet_leaf_0_clk),
    .D(_0103_),
    .Q(\outputs.divider_buffer2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2898_ (.CLK(clknet_leaf_1_clk),
    .D(_0104_),
    .Q(\outputs.divider_buffer2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2899_ (.CLK(clknet_leaf_0_clk),
    .D(_0105_),
    .Q(\outputs.divider_buffer2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2900_ (.CLK(clknet_leaf_3_clk),
    .D(_0106_),
    .Q(\outputs.divider_buffer2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2901_ (.CLK(clknet_leaf_2_clk),
    .D(_0107_),
    .Q(\outputs.divider_buffer2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2902_ (.CLK(clknet_leaf_12_clk),
    .D(_0108_),
    .Q(\outputs.divider_buffer2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2903_ (.CLK(clknet_leaf_12_clk),
    .D(_0109_),
    .Q(\outputs.divider_buffer2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2904_ (.CLK(clknet_leaf_13_clk),
    .D(_0110_),
    .Q(\outputs.divider_buffer2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2905_ (.CLK(clknet_leaf_13_clk),
    .D(_0111_),
    .Q(\outputs.divider_buffer2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2906_ (.CLK(clknet_leaf_12_clk),
    .D(_0112_),
    .Q(\outputs.divider_buffer2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2907_ (.CLK(clknet_leaf_1_clk),
    .D(_0113_),
    .Q(\outputs.div.divisor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2908_ (.CLK(clknet_leaf_34_clk),
    .D(_0114_),
    .Q(\outputs.div.divisor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2909_ (.CLK(clknet_leaf_34_clk),
    .D(_0115_),
    .Q(\outputs.div.divisor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2910_ (.CLK(clknet_leaf_34_clk),
    .D(_0116_),
    .Q(\outputs.div.divisor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2911_ (.CLK(clknet_leaf_34_clk),
    .D(_0117_),
    .Q(\outputs.div.divisor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2912_ (.CLK(clknet_leaf_34_clk),
    .D(_0118_),
    .Q(\outputs.div.divisor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2913_ (.CLK(clknet_leaf_34_clk),
    .D(_0119_),
    .Q(\outputs.div.divisor[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2914_ (.CLK(clknet_leaf_34_clk),
    .D(_0120_),
    .Q(\outputs.div.divisor[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2915_ (.CLK(clknet_leaf_1_clk),
    .D(_0121_),
    .Q(\outputs.div.divisor[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2916_ (.CLK(clknet_leaf_1_clk),
    .D(_0122_),
    .Q(\outputs.div.divisor[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2917_ (.CLK(clknet_leaf_1_clk),
    .D(_0123_),
    .Q(\outputs.div.divisor[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2918_ (.CLK(clknet_leaf_1_clk),
    .D(_0124_),
    .Q(\outputs.div.divisor[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2919_ (.CLK(clknet_leaf_1_clk),
    .D(_0125_),
    .Q(\outputs.div.divisor[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2920_ (.CLK(clknet_leaf_12_clk),
    .D(_0126_),
    .Q(\outputs.div.divisor[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2921_ (.CLK(clknet_leaf_13_clk),
    .D(_0127_),
    .Q(\outputs.div.divisor[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2922_ (.CLK(clknet_leaf_13_clk),
    .D(_0128_),
    .Q(\outputs.div.divisor[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2923_ (.CLK(clknet_leaf_13_clk),
    .D(_0129_),
    .Q(\outputs.div.divisor[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2924_ (.CLK(clknet_leaf_12_clk),
    .D(_0130_),
    .Q(\outputs.div.divisor[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2925_ (.CLK(clknet_leaf_1_clk),
    .D(_0131_),
    .RESET_B(net38),
    .Q(\outputs.divider_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2926_ (.CLK(clknet_leaf_1_clk),
    .D(_0132_),
    .RESET_B(net38),
    .Q(\outputs.divider_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2927_ (.CLK(clknet_leaf_1_clk),
    .D(_0133_),
    .RESET_B(net38),
    .Q(\outputs.divider_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2928_ (.CLK(clknet_leaf_1_clk),
    .D(_0134_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2929_ (.CLK(clknet_leaf_0_clk),
    .D(_0135_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2930_ (.CLK(clknet_leaf_0_clk),
    .D(_0136_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2931_ (.CLK(clknet_leaf_0_clk),
    .D(_0137_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2932_ (.CLK(clknet_leaf_0_clk),
    .D(_0138_),
    .RESET_B(net25),
    .Q(\outputs.divider_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2933_ (.CLK(clknet_leaf_39_clk),
    .D(_0139_),
    .RESET_B(net25),
    .Q(\outputs.divider_buffer[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2934_ (.CLK(clknet_leaf_2_clk),
    .D(_0140_),
    .RESET_B(net38),
    .Q(\outputs.divider_buffer[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2935_ (.CLK(clknet_leaf_39_clk),
    .D(_0141_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2936_ (.CLK(clknet_leaf_3_clk),
    .D(_0142_),
    .RESET_B(net37),
    .Q(\outputs.divider_buffer[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2937_ (.CLK(clknet_leaf_3_clk),
    .D(_0143_),
    .RESET_B(net37),
    .Q(\outputs.divider_buffer[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2938_ (.CLK(clknet_leaf_12_clk),
    .D(_0144_),
    .RESET_B(net39),
    .Q(\outputs.divider_buffer[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2939_ (.CLK(clknet_leaf_12_clk),
    .D(_0145_),
    .RESET_B(net39),
    .Q(\outputs.divider_buffer[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2940_ (.CLK(clknet_leaf_12_clk),
    .D(_0146_),
    .RESET_B(net46),
    .Q(\outputs.divider_buffer[15] ));
 sky130_fd_sc_hd__dfrtp_2 _2941_ (.CLK(clknet_leaf_14_clk),
    .D(_0147_),
    .RESET_B(net46),
    .Q(\outputs.divider_buffer[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2942_ (.CLK(clknet_leaf_12_clk),
    .D(_0148_),
    .RESET_B(net39),
    .Q(\outputs.divider_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2943_ (.CLK(clknet_leaf_15_clk),
    .D(_0149_),
    .Q(\outputs.signal_buffer2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2944_ (.CLK(clknet_leaf_12_clk),
    .D(_0150_),
    .Q(\outputs.signal_buffer2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2945_ (.CLK(clknet_leaf_10_clk),
    .D(_0151_),
    .Q(\outputs.signal_buffer2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2946_ (.CLK(clknet_leaf_10_clk),
    .D(_0152_),
    .Q(\outputs.signal_buffer2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2947_ (.CLK(clknet_leaf_8_clk),
    .D(_0153_),
    .Q(\outputs.signal_buffer2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2948_ (.CLK(clknet_leaf_8_clk),
    .D(_0154_),
    .Q(\outputs.signal_buffer2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2949_ (.CLK(clknet_leaf_5_clk),
    .D(_0155_),
    .Q(\outputs.signal_buffer2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2950_ (.CLK(clknet_leaf_4_clk),
    .D(_0156_),
    .Q(\outputs.signal_buffer2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2951_ (.CLK(clknet_leaf_5_clk),
    .D(_0157_),
    .Q(\outputs.signal_buffer2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2952_ (.CLK(clknet_leaf_4_clk),
    .D(_0158_),
    .Q(\outputs.signal_buffer2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2953_ (.CLK(clknet_leaf_4_clk),
    .D(_0159_),
    .Q(\outputs.signal_buffer2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2954_ (.CLK(clknet_leaf_6_clk),
    .D(_0160_),
    .Q(\outputs.signal_buffer2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2955_ (.CLK(clknet_leaf_5_clk),
    .D(_0161_),
    .Q(\outputs.signal_buffer2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2956_ (.CLK(clknet_leaf_7_clk),
    .D(_0162_),
    .Q(\outputs.signal_buffer2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2957_ (.CLK(clknet_leaf_7_clk),
    .D(_0163_),
    .Q(\outputs.signal_buffer2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2958_ (.CLK(clknet_leaf_8_clk),
    .D(_0164_),
    .Q(\outputs.signal_buffer2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2959_ (.CLK(clknet_leaf_8_clk),
    .D(_0165_),
    .Q(\outputs.signal_buffer2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2960_ (.CLK(clknet_leaf_9_clk),
    .D(_0166_),
    .Q(\outputs.signal_buffer2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2961_ (.CLK(clknet_leaf_10_clk),
    .D(_0167_),
    .Q(\outputs.div.oscillator_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2962_ (.CLK(clknet_leaf_10_clk),
    .D(_0168_),
    .Q(\outputs.div.oscillator_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2963_ (.CLK(clknet_leaf_10_clk),
    .D(_0169_),
    .Q(\outputs.div.oscillator_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2964_ (.CLK(clknet_leaf_10_clk),
    .D(_0170_),
    .Q(\outputs.div.oscillator_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2965_ (.CLK(clknet_leaf_8_clk),
    .D(_0171_),
    .Q(\outputs.div.oscillator_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2966_ (.CLK(clknet_leaf_7_clk),
    .D(_0172_),
    .Q(\outputs.div.oscillator_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2967_ (.CLK(clknet_leaf_5_clk),
    .D(_0173_),
    .Q(\outputs.div.oscillator_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2968_ (.CLK(clknet_leaf_4_clk),
    .D(_0174_),
    .Q(\outputs.div.oscillator_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2969_ (.CLK(clknet_leaf_5_clk),
    .D(_0175_),
    .Q(\outputs.div.oscillator_out[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2970_ (.CLK(clknet_leaf_4_clk),
    .D(_0176_),
    .Q(\outputs.div.oscillator_out[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2971_ (.CLK(clknet_leaf_4_clk),
    .D(_0177_),
    .Q(\outputs.div.oscillator_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2972_ (.CLK(clknet_leaf_6_clk),
    .D(_0178_),
    .Q(\outputs.div.oscillator_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2973_ (.CLK(clknet_leaf_5_clk),
    .D(_0179_),
    .Q(\outputs.div.oscillator_out[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2974_ (.CLK(clknet_leaf_7_clk),
    .D(_0180_),
    .Q(\outputs.div.oscillator_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2975_ (.CLK(clknet_leaf_7_clk),
    .D(_0181_),
    .Q(\outputs.div.oscillator_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2976_ (.CLK(clknet_leaf_7_clk),
    .D(_0182_),
    .Q(\outputs.div.oscillator_out[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2977_ (.CLK(clknet_leaf_8_clk),
    .D(_0183_),
    .Q(\outputs.div.oscillator_out[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2978_ (.CLK(clknet_leaf_9_clk),
    .D(_0184_),
    .Q(\outputs.div.oscillator_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2979_ (.CLK(clknet_leaf_15_clk),
    .D(_0185_),
    .RESET_B(net50),
    .Q(\outputs.shaper.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2980_ (.CLK(clknet_leaf_12_clk),
    .D(_0186_),
    .RESET_B(net39),
    .Q(\outputs.shaper.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2981_ (.CLK(clknet_leaf_12_clk),
    .D(_0187_),
    .RESET_B(net39),
    .Q(\outputs.shaper.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2982_ (.CLK(clknet_leaf_10_clk),
    .D(_0188_),
    .RESET_B(net44),
    .Q(\outputs.shaper.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2983_ (.CLK(clknet_leaf_10_clk),
    .D(_0189_),
    .RESET_B(net44),
    .Q(\outputs.shaper.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2984_ (.CLK(clknet_leaf_8_clk),
    .D(_0190_),
    .RESET_B(net43),
    .Q(\outputs.shaper.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2985_ (.CLK(clknet_leaf_7_clk),
    .D(_0191_),
    .RESET_B(net42),
    .Q(\outputs.shaper.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2986_ (.CLK(clknet_leaf_5_clk),
    .D(_0192_),
    .RESET_B(net37),
    .Q(\outputs.shaper.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2987_ (.CLK(clknet_leaf_4_clk),
    .D(_0193_),
    .RESET_B(net37),
    .Q(\outputs.shaper.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2988_ (.CLK(clknet_leaf_4_clk),
    .D(_0194_),
    .RESET_B(net40),
    .Q(\outputs.shaper.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2989_ (.CLK(clknet_leaf_4_clk),
    .D(_0195_),
    .RESET_B(net40),
    .Q(\outputs.shaper.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2990_ (.CLK(clknet_leaf_6_clk),
    .D(_0196_),
    .RESET_B(net42),
    .Q(\outputs.shaper.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2991_ (.CLK(clknet_leaf_5_clk),
    .D(_0197_),
    .RESET_B(net42),
    .Q(\outputs.shaper.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2992_ (.CLK(clknet_leaf_7_clk),
    .D(_0198_),
    .RESET_B(net42),
    .Q(\outputs.shaper.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2993_ (.CLK(clknet_leaf_7_clk),
    .D(_0199_),
    .RESET_B(net42),
    .Q(\outputs.shaper.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2994_ (.CLK(clknet_leaf_8_clk),
    .D(_0200_),
    .RESET_B(net43),
    .Q(\outputs.shaper.count[15] ));
 sky130_fd_sc_hd__dfrtp_2 _2995_ (.CLK(clknet_leaf_9_clk),
    .D(_0201_),
    .RESET_B(net43),
    .Q(\outputs.shaper.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2996_ (.CLK(clknet_leaf_9_clk),
    .D(_0202_),
    .RESET_B(net44),
    .Q(\outputs.shaper.count[17] ));
 sky130_fd_sc_hd__dfstp_1 _2997_ (.CLK(clknet_leaf_36_clk),
    .D(_0203_),
    .SET_B(net24),
    .Q(\inputs.frequency_lut.rng[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2998_ (.CLK(clknet_leaf_36_clk),
    .D(_0204_),
    .RESET_B(net24),
    .Q(\inputs.frequency_lut.rng[1] ));
 sky130_fd_sc_hd__dfstp_1 _2999_ (.CLK(clknet_leaf_37_clk),
    .D(_0205_),
    .SET_B(net23),
    .Q(\inputs.frequency_lut.rng[2] ));
 sky130_fd_sc_hd__dfstp_1 _3000_ (.CLK(clknet_leaf_37_clk),
    .D(_0206_),
    .SET_B(net23),
    .Q(\inputs.frequency_lut.rng[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3001_ (.CLK(clknet_leaf_36_clk),
    .D(_0207_),
    .RESET_B(net24),
    .Q(\inputs.frequency_lut.rng[4] ));
 sky130_fd_sc_hd__dfstp_2 _3002_ (.CLK(clknet_leaf_35_clk),
    .D(_0208_),
    .SET_B(net24),
    .Q(\inputs.frequency_lut.rng[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3003_ (.CLK(clknet_leaf_28_clk),
    .D(net62),
    .RESET_B(net35),
    .Q(\outputs.pwm_output ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(net24),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net19),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net19),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net36),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(net31),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net36),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net36),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net36),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net19),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net40),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net55),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net55),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net55),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net55),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(net55),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net49),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net55),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net54),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net54),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net19),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\inputs.keypad_synchronizer.half_sync[7] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\inputs.keypad_synchronizer.half_sync[3] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\outputs.div.oscillator_out[0] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0055_),
    .X(net156));
 sky130_fd_sc_hd__buf_1 hold102 (.A(\inputs.random_update_clock.count[0] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\outputs.div.a[16] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\outputs.div.oscillator_out[17] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0072_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\outputs.div.a[8] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\outputs.div.count[2] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\outputs.div.q_out[3] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0090_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\inputs.keypad_synchronizer.half_sync[1] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\outputs.div.a[12] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\inputs.random_update_clock.count[14] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_1059_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\inputs.random_update_clock.count[16] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\outputs.div.a[6] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\outputs.div.a[23] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\outputs.div.q_out[7] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0094_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\outputs.div.a[5] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\inputs.random_update_clock.count[1] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\inputs.random_note_generator.out[11] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\outputs.div.a[10] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\inputs.random_update_clock.count[4] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\inputs.random_update_clock.count[20] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_1067_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\outputs.div.a[11] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\outputs.sample_rate.count[6] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\outputs.div.a[1] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\outputs.div.a[13] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\inputs.wavetype_fsm.state[1] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\inputs.wavetype_fsm.next_state[1] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\inputs.random_note_generator.out[8] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\outputs.div.a[7] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\outputs.sig_gen.count[17] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\inputs.random_update_clock.count[15] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\outputs.signal_buffer2[2] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0963_),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\inputs.random_update_clock.count[19] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\inputs.random_update_clock.count[11] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\outputs.div.a[15] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\outputs.sig_gen.count[0] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\inputs.random_update_clock.count[2] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\inputs.keypad_synchronizer.half_sync[2] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\outputs.divider_buffer2[15] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\inputs.random_update_clock.count[9] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\outputs.div.q[5] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\inputs.random_update_clock.count[3] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\outputs.div.q[6] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0054_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\outputs.div.q_out[2] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0089_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\outputs.div.a[2] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\outputs.sample_rate.count[7] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\inputs.random_note_generator.out[5] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\outputs.signal_buffer2[7] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\outputs.signal_buffer2[6] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\outputs.signal_buffer2[16] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\outputs.div.divisor[6] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\outputs.signal_buffer2[9] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\outputs.div.q[3] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\outputs.div.count[4] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\inputs.random_update_clock.count[7] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\outputs.div.q[1] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0049_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\inputs.random_note_generator.out[7] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\outputs.signal_buffer2[5] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\inputs.random_update_clock.count[6] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\outputs.div.divisor[9] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\outputs.output_gen.count[2] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_1073_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\outputs.div.divisor[15] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\outputs.div.oscillator_out[7] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\outputs.div.a[21] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\outputs.signal_buffer2[12] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\outputs.divider_buffer2[6] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\inputs.random_note_generator.out[14] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\outputs.div.oscillator_out[2] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\outputs.divider_buffer2[12] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\outputs.output_gen.count[5] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\outputs.signal_buffer2[11] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0934_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\outputs.signal_buffer2[17] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\outputs.divider_buffer2[7] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\outputs.signal_buffer2[13] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0937_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\outputs.signal_buffer2[1] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\inputs.random_note_generator.out[3] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0923_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\outputs.output_gen.count[4] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\outputs.signal_buffer2[0] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\outputs.signal_buffer2[15] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\outputs.divider_buffer2[4] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0518_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\outputs.divider_buffer2[1] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0515_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\outputs.signal_buffer2[10] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0933_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\inputs.keypad_synchronizer.half_sync[16] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\outputs.divider_buffer2[8] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\outputs.divider_buffer2[11] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0526_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\outputs.divider_buffer2[17] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\outputs.signal_buffer2[4] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\outputs.div.q[2] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\outputs.divider_buffer2[3] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0517_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\outputs.div.divisor[9] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\outputs.signal_buffer2[14] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\inputs.keypad_synchronizer.half_sync[5] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\inputs.random_note_generator.out[9] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\outputs.divider_buffer2[0] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\outputs.div.a[18] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\outputs.divider_buffer2[5] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0519_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\outputs.shaper.count[11] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\outputs.div.a[17] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\outputs.div.q[0] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\outputs.signal_buffer2[3] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\outputs.div.count[1] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\outputs.div.q[25] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\inputs.random_note_generator.out[1] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0073_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\outputs.divider_buffer2[16] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0531_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\outputs.output_gen.count[3] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\outputs.div.divisor[14] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0529_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\outputs.signal_buffer2[8] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\outputs.divider_buffer2[13] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\outputs.shaper.count[14] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\outputs.div.a[25] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\inputs.keypad_synchronizer.half_sync[14] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\outputs.divider_buffer2[10] ),
    .X(net275));
 sky130_fd_sc_hd__buf_1 hold221 (.A(\outputs.div.divisor[12] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\outputs.div.oscillator_out[8] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\outputs.div.divisor[11] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\outputs.div.divisor[2] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0516_),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\outputs.div.a[20] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\outputs.shaper.count[10] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\outputs.div.a[22] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\inputs.random_update_clock.count[17] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\inputs.keypad_synchronizer.half_sync[13] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_1062_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\outputs.divider_buffer2[14] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0918_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\outputs.div.a[9] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\outputs.div.q_out[4] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\outputs.sig_gen.count[4] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\outputs.divider_buffer2[2] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\outputs.div.divisor[3] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\inputs.random_update_clock.count[5] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\outputs.sig_gen.count[2] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\inputs.keypad_synchronizer.half_sync[6] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\outputs.div.a[19] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\inputs.down.ff_out ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\outputs.div.divisor[0] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\outputs.div.divisor[16] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\outputs.div.a[3] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\outputs.div.oscillator_out[1] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\outputs.sig_gen.count[17] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\outputs.div.oscillator_out[13] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\outputs.scaled_buffer[7] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\outputs.div.oscillator_out[11] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\inputs.keypad_synchronizer.half_sync[15] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\inputs.up.ff_out ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\outputs.div.divisor[13] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\inputs.random_update_clock.count[18] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\outputs.div.divisor[8] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\outputs.div.oscillator_out[10] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\outputs.div.divisor[1] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\outputs.div.divisor[4] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\outputs.div.divisor[12] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\outputs.div.divisor[15] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\outputs.output_gen.count[4] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\inputs.random_note_generator.out[6] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\outputs.div.divisor[2] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\outputs.div.divisor[6] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\outputs.div.divisor[0] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\outputs.div.divisor[3] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\inputs.random_note_generator.out[12] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\inputs.random_note_generator.out[0] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\inputs.random_note_generator.out[4] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\inputs.random_note_generator.out[2] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\inputs.keypad_synchronizer.half_sync[0] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\inputs.random_note_generator.out[12] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\inputs.keypad_synchronizer.half_sync[10] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\inputs.random_note_generator.out[13] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\inputs.key_encoder.octave_key_up ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\inputs.random_note_generator.out[10] ),
    .X(net89));
 sky130_fd_sc_hd__buf_1 hold35 (.A(\outputs.output_gen.count[0] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\outputs.output_gen.next_count[1] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\outputs.div.oscillator_out[3] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0058_),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\inputs.key_encoder.sync_keys[15] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\inputs.keypad_synchronizer.half_sync[11] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\inputs.key_encoder.mode_key ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\inputs.random_update_clock.count[22] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\inputs.random_update_clock.next_count[22] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\outputs.div.oscillator_out[4] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0059_),
    .X(net99));
 sky130_fd_sc_hd__buf_1 hold45 (.A(\outputs.sample_rate.count[0] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\outputs.div.oscillator_out[14] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0069_),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\outputs.div.oscillator_out[15] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0070_),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\inputs.keypad_synchronizer.half_sync[12] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\outputs.div.q_out[1] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0088_),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\outputs.div.oscillator_out[6] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0061_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\outputs.div.oscillator_out[16] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0071_),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\outputs.divider_buffer2[9] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\outputs.sample_rate.count[2] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_1085_),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\outputs.sample_rate.count[1] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\inputs.keypad_synchronizer.half_sync[4] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\inputs.mode_edge.ff_out ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\outputs.div.q[15] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0062_),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\outputs.div.q[19] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0066_),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\outputs.div.q[10] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0057_),
    .X(net121));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold67 (.A(\outputs.div.q[4] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0091_),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\outputs.div.q[16] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\outputs.output_gen.pwm_ff ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0063_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\outputs.div.a[14] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\outputs.div.oscillator_out[12] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0067_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\outputs.div.q_out[0] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0087_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\outputs.sample_rate.count[5] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_1087_),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\outputs.div.a[24] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\outputs.div.q[17] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\inputs.keypad_synchronizer.half_sync[9] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0064_),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\outputs.div.q[9] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0056_),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\outputs.div.q_out[6] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0093_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\outputs.div.a[0] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\outputs.sample_rate.count[4] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\outputs.sample_rate.next_count[4] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\outputs.div.q_out[5] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0092_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\inputs.keypad_synchronizer.half_sync[8] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\outputs.sample_rate.count[3] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\outputs.div.q[18] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0065_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\outputs.output_gen.count[7] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\outputs.output_gen.next_count[7] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\outputs.div.oscillator_out[5] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0060_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\outputs.div.q[21] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0068_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\outputs.div.a[4] ),
    .X(net154));
 sky130_fd_sc_hd__buf_4 input1 (.A(cs),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(gpio[1]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(gpio[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(gpio[3]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(gpio[4]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(gpio[5]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(gpio[6]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(gpio[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(gpio[8]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(gpio[9]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(nrst),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(gpio[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(gpio[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(gpio[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(gpio[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(gpio[13]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(gpio[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(gpio[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(gpio[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(pwm));
 sky130_fd_sc_hd__clkbuf_4 wire21 (.A(_1244_),
    .X(net21));
endmodule

