magic
tech sky130A
magscale 1 2
timestamp 1693970307
<< obsli1 >>
rect 1104 2159 29440 30481
<< obsm1 >>
rect 14 2128 29702 30512
<< metal2 >>
rect 2594 31925 2650 32725
rect 6458 31925 6514 32725
rect 9678 31925 9734 32725
rect 13542 31925 13598 32725
rect 17406 31925 17462 32725
rect 21270 31925 21326 32725
rect 25134 31925 25190 32725
rect 28998 31925 29054 32725
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10966 0 11022 800
rect 14830 0 14886 800
rect 18694 0 18750 800
rect 21914 0 21970 800
rect 25778 0 25834 800
rect 29642 0 29698 800
<< obsm2 >>
rect 20 31869 2538 32042
rect 2706 31869 6402 32042
rect 6570 31869 9622 32042
rect 9790 31869 13486 32042
rect 13654 31869 17350 32042
rect 17518 31869 21214 32042
rect 21382 31869 25078 32042
rect 25246 31869 28942 32042
rect 29110 31869 29696 32042
rect 20 856 29696 31869
rect 130 734 3182 856
rect 3350 734 7046 856
rect 7214 734 10910 856
rect 11078 734 14774 856
rect 14942 734 18638 856
rect 18806 734 21858 856
rect 22026 734 25722 856
rect 25890 734 29586 856
<< metal3 >>
rect 0 31288 800 31408
rect 29781 30608 30581 30728
rect 0 27208 800 27328
rect 29781 26528 30581 26648
rect 0 23128 800 23248
rect 29781 22448 30581 22568
rect 0 19728 800 19848
rect 29781 18368 30581 18488
rect 0 15648 800 15768
rect 29781 14288 30581 14408
rect 0 11568 800 11688
rect 29781 10888 30581 11008
rect 0 7488 800 7608
rect 29781 6808 30581 6928
rect 0 3408 800 3528
rect 29781 2728 30581 2848
<< obsm3 >>
rect 880 31208 29930 31378
rect 798 30808 29930 31208
rect 798 30528 29701 30808
rect 798 27408 29930 30528
rect 880 27128 29930 27408
rect 798 26728 29930 27128
rect 798 26448 29701 26728
rect 798 23328 29930 26448
rect 880 23048 29930 23328
rect 798 22648 29930 23048
rect 798 22368 29701 22648
rect 798 19928 29930 22368
rect 880 19648 29930 19928
rect 798 18568 29930 19648
rect 798 18288 29701 18568
rect 798 15848 29930 18288
rect 880 15568 29930 15848
rect 798 14488 29930 15568
rect 798 14208 29701 14488
rect 798 11768 29930 14208
rect 880 11488 29930 11768
rect 798 11088 29930 11488
rect 798 10808 29701 11088
rect 798 7688 29930 10808
rect 880 7408 29930 7688
rect 798 7008 29930 7408
rect 798 6728 29701 7008
rect 798 3608 29930 6728
rect 880 3328 29930 3608
rect 798 2928 29930 3328
rect 798 2648 29701 2928
rect 798 2143 29930 2648
<< metal4 >>
rect 4485 2128 4805 30512
rect 8026 2128 8346 30512
rect 11568 2128 11888 30512
rect 15109 2128 15429 30512
rect 18651 2128 18971 30512
rect 22192 2128 22512 30512
rect 25734 2128 26054 30512
rect 29275 2128 29595 30512
<< obsm4 >>
rect 10179 5475 11488 29069
rect 11968 5475 15029 29069
rect 15509 5475 18571 29069
rect 19051 5475 22112 29069
rect 22592 5475 25654 29069
rect 26134 5475 28829 29069
<< labels >>
rlabel metal3 s 0 7488 800 7608 6 clk
port 1 nsew signal input
rlabel metal2 s 28998 31925 29054 32725 6 nrst
port 2 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 out_0[0]
port 3 nsew signal output
rlabel metal2 s 9678 31925 9734 32725 6 out_0[1]
port 4 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 out_0[2]
port 5 nsew signal output
rlabel metal3 s 29781 10888 30581 11008 6 out_0[3]
port 6 nsew signal output
rlabel metal2 s 17406 31925 17462 32725 6 out_0[4]
port 7 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 out_0[5]
port 8 nsew signal output
rlabel metal3 s 29781 18368 30581 18488 6 out_0[6]
port 9 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 out_1[0]
port 10 nsew signal output
rlabel metal3 s 29781 22448 30581 22568 6 out_1[1]
port 11 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 out_1[2]
port 12 nsew signal output
rlabel metal2 s 18 0 74 800 6 out_1[3]
port 13 nsew signal output
rlabel metal2 s 21270 31925 21326 32725 6 out_1[4]
port 14 nsew signal output
rlabel metal2 s 25134 31925 25190 32725 6 out_1[5]
port 15 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 out_1[6]
port 16 nsew signal output
rlabel metal2 s 6458 31925 6514 32725 6 out_2[0]
port 17 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 out_2[1]
port 18 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 out_2[2]
port 19 nsew signal output
rlabel metal3 s 29781 2728 30581 2848 6 out_2[3]
port 20 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 out_2[4]
port 21 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 out_2[5]
port 22 nsew signal output
rlabel metal2 s 2594 31925 2650 32725 6 out_2[6]
port 23 nsew signal output
rlabel metal3 s 29781 6808 30581 6928 6 out_3[0]
port 24 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 out_3[1]
port 25 nsew signal output
rlabel metal3 s 29781 26528 30581 26648 6 out_3[2]
port 26 nsew signal output
rlabel metal3 s 29781 30608 30581 30728 6 out_3[3]
port 27 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 out_3[4]
port 28 nsew signal output
rlabel metal2 s 13542 31925 13598 32725 6 out_3[5]
port 29 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 out_3[6]
port 30 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 pb_0
port 31 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 pb_1
port 32 nsew signal input
rlabel metal3 s 29781 14288 30581 14408 6 time_done
port 33 nsew signal output
rlabel metal4 s 4485 2128 4805 30512 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 11568 2128 11888 30512 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 18651 2128 18971 30512 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 25734 2128 26054 30512 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 8026 2128 8346 30512 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 15109 2128 15429 30512 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 22192 2128 22512 30512 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 29275 2128 29595 30512 6 vssd1
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30581 32725
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2965024
string GDS_FILE /home/designer-25/CUP/openlane/stopwatch/runs/23_09_05_20_15/results/signoff/stopwatch.magic.gds
string GDS_START 731616
<< end >>

