VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Synthia
  CLASS BLOCK ;
  FOREIGN Synthia ;
  ORIGIN 0.000 0.000 ;
  SIZE 268.400 BY 279.120 ;
  PIN PWM_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 264.400 27.240 268.400 27.840 ;
    END
  END PWM_o
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 266.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 262.900 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 262.900 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 266.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 262.900 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 262.900 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 264.400 214.240 268.400 214.840 ;
    END
  END clk
  PIN modes
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 275.120 151.710 279.120 ;
    END
  END modes
  PIN octaves
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END octaves
  PIN pb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END pb[0]
  PIN pb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 275.120 90.530 279.120 ;
    END
  END pb[10]
  PIN pb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END pb[11]
  PIN pb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 267.350 275.120 267.630 279.120 ;
    END
  END pb[12]
  PIN pb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END pb[1]
  PIN pb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END pb[2]
  PIN pb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END pb[3]
  PIN pb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 264.400 153.040 268.400 153.640 ;
    END
  END pb[4]
  PIN pb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END pb[5]
  PIN pb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 275.120 209.670 279.120 ;
    END
  END pb[6]
  PIN pb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END pb[7]
  PIN pb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END pb[8]
  PIN pb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 275.120 32.570 279.120 ;
    END
  END pb[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 264.400 88.440 268.400 89.040 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 262.660 266.645 ;
      LAYER met1 ;
        RECT 0.070 10.640 267.650 266.800 ;
      LAYER met2 ;
        RECT 0.100 274.840 32.010 275.120 ;
        RECT 32.850 274.840 89.970 275.120 ;
        RECT 90.810 274.840 151.150 275.120 ;
        RECT 151.990 274.840 209.110 275.120 ;
        RECT 209.950 274.840 267.070 275.120 ;
        RECT 0.100 4.280 267.620 274.840 ;
        RECT 0.650 4.000 57.770 4.280 ;
        RECT 58.610 4.000 115.730 4.280 ;
        RECT 116.570 4.000 176.910 4.280 ;
        RECT 177.750 4.000 234.870 4.280 ;
        RECT 235.710 4.000 267.620 4.280 ;
      LAYER met3 ;
        RECT 4.000 249.240 264.400 266.725 ;
        RECT 4.400 247.840 264.400 249.240 ;
        RECT 4.000 215.240 264.400 247.840 ;
        RECT 4.000 213.840 264.000 215.240 ;
        RECT 4.000 188.040 264.400 213.840 ;
        RECT 4.400 186.640 264.400 188.040 ;
        RECT 4.000 154.040 264.400 186.640 ;
        RECT 4.000 152.640 264.000 154.040 ;
        RECT 4.000 123.440 264.400 152.640 ;
        RECT 4.400 122.040 264.400 123.440 ;
        RECT 4.000 89.440 264.400 122.040 ;
        RECT 4.000 88.040 264.000 89.440 ;
        RECT 4.000 62.240 264.400 88.040 ;
        RECT 4.400 60.840 264.400 62.240 ;
        RECT 4.000 28.240 264.400 60.840 ;
        RECT 4.000 26.840 264.000 28.240 ;
        RECT 4.000 10.715 264.400 26.840 ;
      LAYER met4 ;
        RECT 49.975 32.135 79.745 241.905 ;
  END
END Synthia
END LIBRARY

