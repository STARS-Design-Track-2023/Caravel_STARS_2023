VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Guitar_Villains
  CLASS BLOCK ;
  FOREIGN Guitar_Villains ;
  ORIGIN 0.000 0.000 ;
  SIZE 317.825 BY 328.545 ;
  PIN bottom_row[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END bottom_row[0]
  PIN bottom_row[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END bottom_row[1]
  PIN bottom_row[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 324.545 61.550 328.545 ;
    END
  END bottom_row[2]
  PIN bottom_row[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 267.350 324.545 267.630 328.545 ;
    END
  END bottom_row[3]
  PIN bottom_row[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END bottom_row[4]
  PIN bottom_row[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END bottom_row[5]
  PIN bottom_row[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END bottom_row[6]
  PIN button[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 324.545 232.210 328.545 ;
    END
  END button[0]
  PIN button[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END button[1]
  PIN button[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 313.825 200.640 317.825 201.240 ;
    END
  END button[2]
  PIN button[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 324.545 196.790 328.545 ;
    END
  END button[3]
  PIN chip_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END chip_select
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END clk
  PIN green_disp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 313.825 20.440 317.825 21.040 ;
    END
  END green_disp
  PIN n_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 313.825 166.640 317.825 167.240 ;
    END
  END n_rst
  PIN red_disp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 313.825 238.040 317.825 238.640 ;
    END
  END red_disp
  PIN ss0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END ss0[0]
  PIN ss0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 324.545 164.590 328.545 ;
    END
  END ss0[1]
  PIN ss0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END ss0[2]
  PIN ss0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 324.545 96.970 328.545 ;
    END
  END ss0[3]
  PIN ss0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 324.545 26.130 328.545 ;
    END
  END ss0[4]
  PIN ss0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END ss0[5]
  PIN ss0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 324.545 299.830 328.545 ;
    END
  END ss0[6]
  PIN ss1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 313.825 57.840 317.825 58.440 ;
    END
  END ss1[0]
  PIN ss1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END ss1[1]
  PIN ss1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END ss1[2]
  PIN ss1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END ss1[3]
  PIN ss1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 313.825 95.240 317.825 95.840 ;
    END
  END ss1[4]
  PIN ss1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END ss1[5]
  PIN ss1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 313.825 275.440 317.825 276.040 ;
    END
  END ss1[6]
  PIN top_row[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 313.825 309.440 317.825 310.040 ;
    END
  END top_row[0]
  PIN top_row[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END top_row[1]
  PIN top_row[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 128.890 324.545 129.170 328.545 ;
    END
  END top_row[2]
  PIN top_row[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END top_row[3]
  PIN top_row[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END top_row[4]
  PIN top_row[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END top_row[5]
  PIN top_row[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 313.825 129.240 317.825 129.840 ;
    END
  END top_row[6]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 315.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 315.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 311.880 315.605 ;
      LAYER met1 ;
        RECT 0.070 10.640 312.270 315.760 ;
      LAYER met2 ;
        RECT 0.100 324.265 25.570 324.545 ;
        RECT 26.410 324.265 60.990 324.545 ;
        RECT 61.830 324.265 96.410 324.545 ;
        RECT 97.250 324.265 128.610 324.545 ;
        RECT 129.450 324.265 164.030 324.545 ;
        RECT 164.870 324.265 196.230 324.545 ;
        RECT 197.070 324.265 231.650 324.545 ;
        RECT 232.490 324.265 267.070 324.545 ;
        RECT 267.910 324.265 299.270 324.545 ;
        RECT 300.110 324.265 312.250 324.545 ;
        RECT 0.100 4.280 312.250 324.265 ;
        RECT 0.650 3.670 32.010 4.280 ;
        RECT 32.850 3.670 67.430 4.280 ;
        RECT 68.270 3.670 99.630 4.280 ;
        RECT 100.470 3.670 135.050 4.280 ;
        RECT 135.890 3.670 167.250 4.280 ;
        RECT 168.090 3.670 202.670 4.280 ;
        RECT 203.510 3.670 238.090 4.280 ;
        RECT 238.930 3.670 270.290 4.280 ;
        RECT 271.130 3.670 305.710 4.280 ;
        RECT 306.550 3.670 312.250 4.280 ;
      LAYER met3 ;
        RECT 4.400 322.640 313.825 323.505 ;
        RECT 3.990 310.440 313.825 322.640 ;
        RECT 3.990 309.040 313.425 310.440 ;
        RECT 3.990 286.640 313.825 309.040 ;
        RECT 4.400 285.240 313.825 286.640 ;
        RECT 3.990 276.440 313.825 285.240 ;
        RECT 3.990 275.040 313.425 276.440 ;
        RECT 3.990 252.640 313.825 275.040 ;
        RECT 4.400 251.240 313.825 252.640 ;
        RECT 3.990 239.040 313.825 251.240 ;
        RECT 3.990 237.640 313.425 239.040 ;
        RECT 3.990 215.240 313.825 237.640 ;
        RECT 4.400 213.840 313.825 215.240 ;
        RECT 3.990 201.640 313.825 213.840 ;
        RECT 3.990 200.240 313.425 201.640 ;
        RECT 3.990 177.840 313.825 200.240 ;
        RECT 4.400 176.440 313.825 177.840 ;
        RECT 3.990 167.640 313.825 176.440 ;
        RECT 3.990 166.240 313.425 167.640 ;
        RECT 3.990 143.840 313.825 166.240 ;
        RECT 4.400 142.440 313.825 143.840 ;
        RECT 3.990 130.240 313.825 142.440 ;
        RECT 3.990 128.840 313.425 130.240 ;
        RECT 3.990 106.440 313.825 128.840 ;
        RECT 4.400 105.040 313.825 106.440 ;
        RECT 3.990 96.240 313.825 105.040 ;
        RECT 3.990 94.840 313.425 96.240 ;
        RECT 3.990 72.440 313.825 94.840 ;
        RECT 4.400 71.040 313.825 72.440 ;
        RECT 3.990 58.840 313.825 71.040 ;
        RECT 3.990 57.440 313.425 58.840 ;
        RECT 3.990 35.040 313.825 57.440 ;
        RECT 4.400 33.640 313.825 35.040 ;
        RECT 3.990 21.440 313.825 33.640 ;
        RECT 3.990 20.040 313.425 21.440 ;
        RECT 3.990 10.715 313.825 20.040 ;
      LAYER met4 ;
        RECT 61.015 11.735 97.440 311.265 ;
        RECT 99.840 11.735 174.240 311.265 ;
        RECT 176.640 11.735 251.040 311.265 ;
        RECT 253.440 11.735 280.305 311.265 ;
  END
END Guitar_Villains
END LIBRARY

