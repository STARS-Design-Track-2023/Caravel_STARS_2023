VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_asic
  CLASS BLOCK ;
  FOREIGN top_asic ;
  ORIGIN 0.000 0.000 ;
  SIZE 436.300 BY 447.020 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 432.300 81.640 436.300 82.240 ;
    END
  END clk
  PIN mode_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 434.790 443.020 435.070 447.020 ;
    END
  END mode_out[0]
  PIN mode_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 264.130 443.020 264.410 447.020 ;
    END
  END mode_out[1]
  PIN pb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END pb[0]
  PIN pb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 432.300 357.040 436.300 357.640 ;
    END
  END pb[10]
  PIN pb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END pb[11]
  PIN pb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END pb[12]
  PIN pb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 443.020 177.470 447.020 ;
    END
  END pb[13]
  PIN pb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END pb[14]
  PIN pb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 443.020 90.530 447.020 ;
    END
  END pb[1]
  PIN pb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END pb[2]
  PIN pb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END pb[3]
  PIN pb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END pb[4]
  PIN pb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 432.300 265.240 436.300 265.840 ;
    END
  END pb[5]
  PIN pb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END pb[6]
  PIN pb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 351.070 443.020 351.350 447.020 ;
    END
  END pb[7]
  PIN pb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END pb[8]
  PIN pb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END pb[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 3.310 443.020 3.590 447.020 ;
    END
  END reset
  PIN sigout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 432.300 173.440 436.300 174.040 ;
    END
  END sigout
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 435.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 435.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 430.560 435.285 ;
      LAYER met1 ;
        RECT 0.070 10.640 435.090 435.440 ;
      LAYER met2 ;
        RECT 0.100 442.740 3.030 443.770 ;
        RECT 3.870 442.740 89.970 443.770 ;
        RECT 90.810 442.740 176.910 443.770 ;
        RECT 177.750 442.740 263.850 443.770 ;
        RECT 264.690 442.740 350.790 443.770 ;
        RECT 351.630 442.740 434.510 443.770 ;
        RECT 0.100 4.280 435.060 442.740 ;
        RECT 0.650 4.000 83.530 4.280 ;
        RECT 84.370 4.000 170.470 4.280 ;
        RECT 171.310 4.000 257.410 4.280 ;
        RECT 258.250 4.000 344.350 4.280 ;
        RECT 345.190 4.000 431.290 4.280 ;
        RECT 432.130 4.000 435.060 4.280 ;
      LAYER met3 ;
        RECT 3.990 364.840 432.300 435.365 ;
        RECT 4.400 363.440 432.300 364.840 ;
        RECT 3.990 358.040 432.300 363.440 ;
        RECT 3.990 356.640 431.900 358.040 ;
        RECT 3.990 273.040 432.300 356.640 ;
        RECT 4.400 271.640 432.300 273.040 ;
        RECT 3.990 266.240 432.300 271.640 ;
        RECT 3.990 264.840 431.900 266.240 ;
        RECT 3.990 181.240 432.300 264.840 ;
        RECT 4.400 179.840 432.300 181.240 ;
        RECT 3.990 174.440 432.300 179.840 ;
        RECT 3.990 173.040 431.900 174.440 ;
        RECT 3.990 89.440 432.300 173.040 ;
        RECT 4.400 88.040 432.300 89.440 ;
        RECT 3.990 82.640 432.300 88.040 ;
        RECT 3.990 81.240 431.900 82.640 ;
        RECT 3.990 10.715 432.300 81.240 ;
      LAYER met4 ;
        RECT 52.735 36.895 97.440 428.225 ;
        RECT 99.840 36.895 174.240 428.225 ;
        RECT 176.640 36.895 251.040 428.225 ;
        RECT 253.440 36.895 327.840 428.225 ;
        RECT 330.240 36.895 403.585 428.225 ;
  END
END top_asic
END LIBRARY

