magic
tech sky130A
magscale 1 2
timestamp 1693969956
<< obsli1 >>
rect 1104 2159 45172 46257
<< obsm1 >>
rect 14 2128 45342 46288
<< metal2 >>
rect 6458 47681 6514 48481
rect 14830 47681 14886 48481
rect 23846 47681 23902 48481
rect 32862 47681 32918 48481
rect 41878 47681 41934 48481
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
rect 26422 0 26478 800
rect 34794 0 34850 800
rect 43810 0 43866 800
<< obsm2 >>
rect 20 47625 6402 47818
rect 6570 47625 14774 47818
rect 14942 47625 23790 47818
rect 23958 47625 32806 47818
rect 32974 47625 41822 47818
rect 41990 47625 45338 47818
rect 20 856 45338 47625
rect 130 800 8334 856
rect 8502 800 17350 856
rect 17518 800 26366 856
rect 26534 800 34738 856
rect 34906 800 43754 856
rect 43922 800 45338 856
<< metal3 >>
rect 0 46248 800 46368
rect 45537 44208 46337 44328
rect 0 36728 800 36848
rect 45537 34688 46337 34808
rect 0 27888 800 28008
rect 45537 25168 46337 25288
rect 0 18368 800 18488
rect 45537 16328 46337 16448
rect 0 8848 800 8968
rect 45537 6808 46337 6928
<< obsm3 >>
rect 880 46168 45537 46341
rect 800 44408 45537 46168
rect 800 44128 45457 44408
rect 800 36928 45537 44128
rect 880 36648 45537 36928
rect 800 34888 45537 36648
rect 800 34608 45457 34888
rect 800 28088 45537 34608
rect 880 27808 45537 28088
rect 800 25368 45537 27808
rect 800 25088 45457 25368
rect 800 18568 45537 25088
rect 880 18288 45537 18568
rect 800 16528 45537 18288
rect 800 16248 45457 16528
rect 800 9048 45537 16248
rect 880 8768 45537 9048
rect 800 7008 45537 8768
rect 800 6728 45457 7008
rect 800 2143 45537 6728
<< metal4 >>
rect 4208 2128 4528 46288
rect 19568 2128 19888 46288
rect 34928 2128 35248 46288
<< obsm4 >>
rect 12387 6835 19488 34645
rect 19968 6835 33245 34645
<< labels >>
rlabel metal2 s 34794 0 34850 800 6 clk
port 1 nsew signal input
rlabel metal3 s 45537 44208 46337 44328 6 cs
port 2 nsew signal input
rlabel metal2 s 41878 47681 41934 48481 6 gpio[0]
port 3 nsew signal input
rlabel metal2 s 23846 47681 23902 48481 6 gpio[10]
port 4 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 gpio[11]
port 5 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 gpio[12]
port 6 nsew signal input
rlabel metal3 s 45537 6808 46337 6928 6 gpio[13]
port 7 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 gpio[14]
port 8 nsew signal input
rlabel metal3 s 45537 34688 46337 34808 6 gpio[15]
port 9 nsew signal input
rlabel metal2 s 18 0 74 800 6 gpio[16]
port 10 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 gpio[1]
port 11 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 gpio[2]
port 12 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 gpio[3]
port 13 nsew signal input
rlabel metal2 s 14830 47681 14886 48481 6 gpio[4]
port 14 nsew signal input
rlabel metal3 s 45537 25168 46337 25288 6 gpio[5]
port 15 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 gpio[6]
port 16 nsew signal input
rlabel metal2 s 32862 47681 32918 48481 6 gpio[7]
port 17 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 gpio[8]
port 18 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 gpio[9]
port 19 nsew signal input
rlabel metal2 s 6458 47681 6514 48481 6 nrst
port 20 nsew signal input
rlabel metal3 s 45537 16328 46337 16448 6 pwm
port 21 nsew signal output
rlabel metal4 s 4208 2128 4528 46288 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 46288 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 46288 6 vssd1
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 46337 48481
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5263142
string GDS_FILE /home/designer-25/CUP/openlane/silly-sythensizer/runs/23_09_05_20_08/results/signoff/silly_synthesizer.magic.gds
string GDS_START 757944
<< end >>

