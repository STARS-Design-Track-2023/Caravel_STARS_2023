// This is the unpowered netlist.
module synth (clk,
    en,
    n_rst,
    pwm_o,
    keypad_i,
    sound_series);
 input clk;
 input en;
 input n_rst;
 output pwm_o;
 input [14:0] keypad_i;
 output [3:0] sound_series;

 wire \SS_FSM.count[0] ;
 wire \SS_FSM.count[1] ;
 wire \SS_FSM.count[2] ;
 wire \SS_FSM.count[3] ;
 wire \SS_FSM.count[4] ;
 wire \SS_FSM.count[5] ;
 wire \SS_FSM.count[6] ;
 wire \SS_FSM.count[7] ;
 wire \SS_FSM.count[8] ;
 wire \SS_FSM.next_sound[0] ;
 wire \SS_FSM.next_sound[1] ;
 wire \SS_FSM.sound[0] ;
 wire \SS_FSM.sound[1] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire \clk8.count[0] ;
 wire \clk8.count[10] ;
 wire \clk8.count[11] ;
 wire \clk8.count[12] ;
 wire \clk8.count[13] ;
 wire \clk8.count[14] ;
 wire \clk8.count[15] ;
 wire \clk8.count[16] ;
 wire \clk8.count[17] ;
 wire \clk8.count[18] ;
 wire \clk8.count[19] ;
 wire \clk8.count[1] ;
 wire \clk8.count[20] ;
 wire \clk8.count[2] ;
 wire \clk8.count[3] ;
 wire \clk8.count[4] ;
 wire \clk8.count[5] ;
 wire \clk8.count[6] ;
 wire \clk8.count[7] ;
 wire \clk8.count[8] ;
 wire \clk8.count[9] ;
 wire \clk8.next_count[0] ;
 wire \clk8.next_count[10] ;
 wire \clk8.next_count[11] ;
 wire \clk8.next_count[12] ;
 wire \clk8.next_count[13] ;
 wire \clk8.next_count[14] ;
 wire \clk8.next_count[15] ;
 wire \clk8.next_count[16] ;
 wire \clk8.next_count[17] ;
 wire \clk8.next_count[18] ;
 wire \clk8.next_count[19] ;
 wire \clk8.next_count[1] ;
 wire \clk8.next_count[20] ;
 wire \clk8.next_count[2] ;
 wire \clk8.next_count[3] ;
 wire \clk8.next_count[4] ;
 wire \clk8.next_count[5] ;
 wire \clk8.next_count[6] ;
 wire \clk8.next_count[7] ;
 wire \clk8.next_count[8] ;
 wire \clk8.next_count[9] ;
 wire \clk_div.count[0] ;
 wire \clk_div.count[1] ;
 wire \clk_div.count[2] ;
 wire \clk_div.count[3] ;
 wire \clk_div.count[4] ;
 wire \clk_div.count[5] ;
 wire \clk_div.count[6] ;
 wire \clk_div.count[7] ;
 wire \clk_div.next_count[0] ;
 wire \clk_div.next_count[1] ;
 wire \clk_div.next_count[2] ;
 wire \clk_div.next_count[3] ;
 wire \clk_div.next_count[4] ;
 wire \clk_div.next_count[5] ;
 wire \clk_div.next_count[6] ;
 wire \clk_div.next_count[7] ;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire \kp_encoder.last_mk ;
 wire \kp_encoder.last_sk ;
 wire \kp_encoder.q[0] ;
 wire \kp_encoder.q[10] ;
 wire \kp_encoder.q[11] ;
 wire \kp_encoder.q[12] ;
 wire \kp_encoder.q[13] ;
 wire \kp_encoder.q[14] ;
 wire \kp_encoder.q[1] ;
 wire \kp_encoder.q[2] ;
 wire \kp_encoder.q[3] ;
 wire \kp_encoder.q[4] ;
 wire \kp_encoder.q[5] ;
 wire \kp_encoder.q[6] ;
 wire \kp_encoder.q[7] ;
 wire \kp_encoder.q[8] ;
 wire \kp_encoder.q[9] ;
 wire \kp_encoder.sync_out[0] ;
 wire \kp_encoder.sync_out[10] ;
 wire \kp_encoder.sync_out[11] ;
 wire \kp_encoder.sync_out[12] ;
 wire \kp_encoder.sync_out[13] ;
 wire \kp_encoder.sync_out[14] ;
 wire \kp_encoder.sync_out[1] ;
 wire \kp_encoder.sync_out[2] ;
 wire \kp_encoder.sync_out[3] ;
 wire \kp_encoder.sync_out[4] ;
 wire \kp_encoder.sync_out[5] ;
 wire \kp_encoder.sync_out[6] ;
 wire \kp_encoder.sync_out[7] ;
 wire \kp_encoder.sync_out[8] ;
 wire \kp_encoder.sync_out[9] ;
 wire \mode_FSM.mode[0] ;
 wire \mode_FSM.mode[1] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \osc.count[0] ;
 wire \osc.count[10] ;
 wire \osc.count[11] ;
 wire \osc.count[12] ;
 wire \osc.count[13] ;
 wire \osc.count[14] ;
 wire \osc.count[15] ;
 wire \osc.count[1] ;
 wire \osc.count[2] ;
 wire \osc.count[3] ;
 wire \osc.count[4] ;
 wire \osc.count[5] ;
 wire \osc.count[6] ;
 wire \osc.count[7] ;
 wire \osc.count[8] ;
 wire \osc.count[9] ;
 wire \osc.next_count[0] ;
 wire \osc.next_count[10] ;
 wire \osc.next_count[11] ;
 wire \osc.next_count[12] ;
 wire \osc.next_count[13] ;
 wire \osc.next_count[14] ;
 wire \osc.next_count[15] ;
 wire \osc.next_count[1] ;
 wire \osc.next_count[2] ;
 wire \osc.next_count[3] ;
 wire \osc.next_count[4] ;
 wire \osc.next_count[5] ;
 wire \osc.next_count[6] ;
 wire \osc.next_count[7] ;
 wire \osc.next_count[8] ;
 wire \osc.next_count[9] ;
 wire \pwm.count[0] ;
 wire \pwm.count[1] ;
 wire \pwm.count[2] ;
 wire \pwm.count[3] ;
 wire \pwm.count[4] ;
 wire \pwm.count[5] ;
 wire \pwm.count[6] ;
 wire \pwm.count[7] ;
 wire \pwm.next_count[0] ;
 wire \pwm.next_count[1] ;
 wire \pwm.next_count[2] ;
 wire \pwm.next_count[3] ;
 wire \pwm.next_count[4] ;
 wire \pwm.next_count[5] ;
 wire \pwm.next_count[6] ;
 wire \pwm.next_count[7] ;
 wire \pwm.pwm ;
 wire \seq_div.D[0] ;
 wire \seq_div.D[10] ;
 wire \seq_div.D[11] ;
 wire \seq_div.D[12] ;
 wire \seq_div.D[13] ;
 wire \seq_div.D[14] ;
 wire \seq_div.D[15] ;
 wire \seq_div.D[1] ;
 wire \seq_div.D[2] ;
 wire \seq_div.D[3] ;
 wire \seq_div.D[4] ;
 wire \seq_div.D[5] ;
 wire \seq_div.D[6] ;
 wire \seq_div.D[7] ;
 wire \seq_div.D[8] ;
 wire \seq_div.D[9] ;
 wire \seq_div.Q[0] ;
 wire \seq_div.Q[1] ;
 wire \seq_div.Q[2] ;
 wire \seq_div.Q[3] ;
 wire \seq_div.Q[4] ;
 wire \seq_div.Q[5] ;
 wire \seq_div.Q[6] ;
 wire \seq_div.Q[7] ;
 wire \seq_div.R[10] ;
 wire \seq_div.R[11] ;
 wire \seq_div.R[12] ;
 wire \seq_div.R[13] ;
 wire \seq_div.R[14] ;
 wire \seq_div.R[15] ;
 wire \seq_div.R[16] ;
 wire \seq_div.R[17] ;
 wire \seq_div.R[18] ;
 wire \seq_div.R[19] ;
 wire \seq_div.R[20] ;
 wire \seq_div.R[21] ;
 wire \seq_div.R[22] ;
 wire \seq_div.R[23] ;
 wire \seq_div.R[8] ;
 wire \seq_div.R[9] ;
 wire \seq_div.count_div[0] ;
 wire \seq_div.count_div[1] ;
 wire \seq_div.count_div[2] ;
 wire \seq_div.dividend[0] ;
 wire \seq_div.dividend[10] ;
 wire \seq_div.dividend[11] ;
 wire \seq_div.dividend[12] ;
 wire \seq_div.dividend[13] ;
 wire \seq_div.dividend[14] ;
 wire \seq_div.dividend[15] ;
 wire \seq_div.dividend[1] ;
 wire \seq_div.dividend[2] ;
 wire \seq_div.dividend[3] ;
 wire \seq_div.dividend[4] ;
 wire \seq_div.dividend[5] ;
 wire \seq_div.dividend[6] ;
 wire \seq_div.dividend[7] ;
 wire \seq_div.dividend[8] ;
 wire \seq_div.dividend[9] ;
 wire \seq_div.q_out[0] ;
 wire \seq_div.q_out[1] ;
 wire \seq_div.q_out[2] ;
 wire \seq_div.q_out[3] ;
 wire \seq_div.q_out[4] ;
 wire \seq_div.q_out[5] ;
 wire \seq_div.q_out[6] ;
 wire \seq_div.q_out[7] ;
 wire \seq_div.state[0] ;
 wire \seq_div.state[1] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_94 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__inv_2 _0779_ (.A(\SS_FSM.count[0] ),
    .Y(_0154_));
 sky130_fd_sc_hd__buf_4 _0780_ (.A(\SS_FSM.count[1] ),
    .X(_0155_));
 sky130_fd_sc_hd__or4_4 _0781_ (.A(\SS_FSM.count[0] ),
    .B(_0155_),
    .C(\SS_FSM.count[3] ),
    .D(\SS_FSM.count[2] ),
    .X(_0156_));
 sky130_fd_sc_hd__nor3_4 _0782_ (.A(\SS_FSM.count[4] ),
    .B(\SS_FSM.count[5] ),
    .C(_0156_),
    .Y(_0157_));
 sky130_fd_sc_hd__o21a_2 _0783_ (.A1(\SS_FSM.count[4] ),
    .A2(_0156_),
    .B1(\SS_FSM.count[5] ),
    .X(_0158_));
 sky130_fd_sc_hd__nor2_8 _0784_ (.A(_0157_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__or3_2 _0785_ (.A(\SS_FSM.count[0] ),
    .B(_0155_),
    .C(\SS_FSM.count[2] ),
    .X(_0160_));
 sky130_fd_sc_hd__o21ai_2 _0786_ (.A1(\SS_FSM.count[0] ),
    .A2(_0155_),
    .B1(\SS_FSM.count[2] ),
    .Y(_0161_));
 sky130_fd_sc_hd__and2_2 _0787_ (.A(_0160_),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__nor4_4 _0788_ (.A(\SS_FSM.count[0] ),
    .B(_0155_),
    .C(\SS_FSM.count[3] ),
    .D(\SS_FSM.count[2] ),
    .Y(_0163_));
 sky130_fd_sc_hd__o31a_2 _0789_ (.A1(\SS_FSM.count[0] ),
    .A2(_0155_),
    .A3(\SS_FSM.count[2] ),
    .B1(\SS_FSM.count[3] ),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_8 _0790_ (.A(_0163_),
    .B(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__xnor2_2 _0791_ (.A(\SS_FSM.count[4] ),
    .B(net27),
    .Y(_0166_));
 sky130_fd_sc_hd__buf_4 _0792_ (.A(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__o211a_1 _0793_ (.A1(_0162_),
    .A2(_0165_),
    .B1(_0167_),
    .C1(\SS_FSM.sound[1] ),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(\SS_FSM.count[6] ),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_1 _0795_ (.A(_0169_),
    .B(net25),
    .Y(_0170_));
 sky130_fd_sc_hd__or2_1 _0796_ (.A(\SS_FSM.count[7] ),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_1 _0797_ (.A(\SS_FSM.count[6] ),
    .B(\SS_FSM.count[7] ),
    .Y(_0172_));
 sky130_fd_sc_hd__nor3_1 _0798_ (.A(\SS_FSM.count[4] ),
    .B(\SS_FSM.count[5] ),
    .C(\SS_FSM.count[8] ),
    .Y(_0173_));
 sky130_fd_sc_hd__and3_1 _0799_ (.A(net27),
    .B(_0172_),
    .C(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_4 _0800_ (.A1(\SS_FSM.count[8] ),
    .A2(_0171_),
    .B1(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__xnor2_4 _0801_ (.A(_0169_),
    .B(net25),
    .Y(_0176_));
 sky130_fd_sc_hd__or2_1 _0802_ (.A(_0157_),
    .B(_0158_),
    .X(_0177_));
 sky130_fd_sc_hd__buf_4 _0803_ (.A(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__buf_4 _0804_ (.A(\SS_FSM.count[0] ),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _0805_ (.A(\SS_FSM.count[6] ),
    .B(\SS_FSM.count[7] ),
    .X(_0180_));
 sky130_fd_sc_hd__or3_1 _0806_ (.A(\SS_FSM.count[4] ),
    .B(\SS_FSM.count[5] ),
    .C(\SS_FSM.count[8] ),
    .X(_0181_));
 sky130_fd_sc_hd__xnor2_1 _0807_ (.A(\SS_FSM.count[0] ),
    .B(_0155_),
    .Y(_0182_));
 sky130_fd_sc_hd__o31a_2 _0808_ (.A1(_0156_),
    .A2(_0180_),
    .A3(_0181_),
    .B1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(_0155_),
    .Y(_0184_));
 sky130_fd_sc_hd__and3_1 _0810_ (.A(_0184_),
    .B(_0160_),
    .C(_0161_),
    .X(_0185_));
 sky130_fd_sc_hd__o21ba_2 _0811_ (.A1(_0162_),
    .A2(_0183_),
    .B1_N(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__or3_1 _0812_ (.A(_0179_),
    .B(_0165_),
    .C(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__or2_1 _0813_ (.A(_0163_),
    .B(_0164_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_4 _0814_ (.A(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__or3_2 _0815_ (.A(_0154_),
    .B(_0155_),
    .C(\SS_FSM.count[2] ),
    .X(_0190_));
 sky130_fd_sc_hd__o21a_1 _0816_ (.A1(_0162_),
    .A2(_0183_),
    .B1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__or2_1 _0817_ (.A(_0189_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__inv_2 _0818_ (.A(\SS_FSM.count[2] ),
    .Y(_0193_));
 sky130_fd_sc_hd__and3_1 _0819_ (.A(_0154_),
    .B(\SS_FSM.count[3] ),
    .C(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__or4_4 _0820_ (.A(_0179_),
    .B(_0162_),
    .C(_0165_),
    .D(_0183_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(\SS_FSM.count[3] ),
    .Y(_0196_));
 sky130_fd_sc_hd__or4_1 _0822_ (.A(_0154_),
    .B(_0184_),
    .C(_0196_),
    .D(\SS_FSM.count[2] ),
    .X(_0197_));
 sky130_fd_sc_hd__or3_2 _0823_ (.A(\SS_FSM.count[0] ),
    .B(_0184_),
    .C(\SS_FSM.count[2] ),
    .X(_0198_));
 sky130_fd_sc_hd__a21o_1 _0824_ (.A1(_0160_),
    .A2(_0161_),
    .B1(_0155_),
    .X(_0199_));
 sky130_fd_sc_hd__a21o_1 _0825_ (.A1(_0198_),
    .A2(_0199_),
    .B1(_0189_),
    .X(_0200_));
 sky130_fd_sc_hd__a31o_1 _0826_ (.A1(_0195_),
    .A2(_0197_),
    .A3(_0200_),
    .B1(_0167_),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _0827_ (.A(_0167_),
    .B(_0194_),
    .Y(_0202_));
 sky130_fd_sc_hd__o211a_1 _0828_ (.A1(_0194_),
    .A2(_0201_),
    .B1(_0202_),
    .C1(_0159_),
    .X(_0203_));
 sky130_fd_sc_hd__a31o_1 _0829_ (.A1(_0178_),
    .A2(_0187_),
    .A3(_0192_),
    .B1(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(\SS_FSM.count[4] ),
    .Y(_0205_));
 sky130_fd_sc_hd__nand2_2 _0831_ (.A(_0205_),
    .B(_0165_),
    .Y(_0206_));
 sky130_fd_sc_hd__nor2_1 _0832_ (.A(_0206_),
    .B(_0191_),
    .Y(_0207_));
 sky130_fd_sc_hd__nor2_1 _0833_ (.A(_0178_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__or3_2 _0834_ (.A(_0156_),
    .B(_0180_),
    .C(_0181_),
    .X(_0209_));
 sky130_fd_sc_hd__or3_2 _0835_ (.A(_0179_),
    .B(_0155_),
    .C(_0193_),
    .X(_0210_));
 sky130_fd_sc_hd__or4_2 _0836_ (.A(\SS_FSM.count[4] ),
    .B(net27),
    .C(_0164_),
    .D(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__or2_1 _0837_ (.A(_0196_),
    .B(_0160_),
    .X(_0212_));
 sky130_fd_sc_hd__or2_1 _0838_ (.A(_0166_),
    .B(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__xnor2_4 _0839_ (.A(\SS_FSM.count[6] ),
    .B(net24),
    .Y(_0214_));
 sky130_fd_sc_hd__a41o_1 _0840_ (.A1(_0209_),
    .A2(_0178_),
    .A3(_0211_),
    .A4(_0213_),
    .B1(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_1 _0841_ (.A(\SS_FSM.count[7] ),
    .B(_0170_),
    .Y(_0216_));
 sky130_fd_sc_hd__and2_1 _0842_ (.A(_0171_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__o221a_1 _0843_ (.A1(_0176_),
    .A2(_0204_),
    .B1(_0208_),
    .B2(_0215_),
    .C1(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_2 _0844_ (.A(_0160_),
    .B(_0161_),
    .Y(_0219_));
 sky130_fd_sc_hd__a21o_1 _0845_ (.A1(_0219_),
    .A2(_0165_),
    .B1(_0174_),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _0846_ (.A(_0159_),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _0847_ (.A(_0179_),
    .B(_0155_),
    .Y(_0222_));
 sky130_fd_sc_hd__a31o_1 _0848_ (.A1(net27),
    .A2(_0172_),
    .A3(_0173_),
    .B1(_0179_),
    .X(_0223_));
 sky130_fd_sc_hd__nand3_1 _0849_ (.A(_0219_),
    .B(_0222_),
    .C(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__or2_1 _0850_ (.A(_0189_),
    .B(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__o22a_1 _0851_ (.A1(_0179_),
    .A2(_0221_),
    .B1(_0225_),
    .B2(_0159_),
    .X(_0226_));
 sky130_fd_sc_hd__o21a_1 _0852_ (.A1(_0167_),
    .A2(_0226_),
    .B1(_0211_),
    .X(_0227_));
 sky130_fd_sc_hd__xnor2_4 _0853_ (.A(_0205_),
    .B(net26),
    .Y(_0228_));
 sky130_fd_sc_hd__o31a_1 _0854_ (.A1(_0179_),
    .A2(_0162_),
    .A3(_0183_),
    .B1(_0190_),
    .X(_0229_));
 sky130_fd_sc_hd__a21o_1 _0855_ (.A1(_0209_),
    .A2(_0210_),
    .B1(_0167_),
    .X(_0230_));
 sky130_fd_sc_hd__o41a_1 _0856_ (.A1(_0169_),
    .A2(_0165_),
    .A3(_0228_),
    .A4(_0229_),
    .B1(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_2 _0857_ (.A(_0171_),
    .B(_0216_),
    .Y(_0232_));
 sky130_fd_sc_hd__o221a_1 _0858_ (.A1(_0176_),
    .A2(_0227_),
    .B1(_0231_),
    .B2(_0159_),
    .C1(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__or3_2 _0859_ (.A(_0180_),
    .B(_0206_),
    .C(_0178_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _0860_ (.A(_0219_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__inv_2 _0861_ (.A(\SS_FSM.sound[1] ),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_2 _0862_ (.A(\SS_FSM.sound[0] ),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__a21oi_1 _0863_ (.A1(_0175_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__o31a_1 _0864_ (.A1(_0175_),
    .A2(_0218_),
    .A3(_0233_),
    .B1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__inv_2 _0865_ (.A(\SS_FSM.sound[0] ),
    .Y(_0240_));
 sky130_fd_sc_hd__a311o_1 _0866_ (.A1(_0154_),
    .A2(_0159_),
    .A3(_0168_),
    .B1(_0239_),
    .C1(_0240_),
    .X(net19));
 sky130_fd_sc_hd__nand2_1 _0867_ (.A(_0159_),
    .B(_0213_),
    .Y(_0241_));
 sky130_fd_sc_hd__nor2_1 _0868_ (.A(_0206_),
    .B(_0186_),
    .Y(_0242_));
 sky130_fd_sc_hd__a21o_1 _0869_ (.A1(_0154_),
    .A2(_0242_),
    .B1(_0159_),
    .X(_0243_));
 sky130_fd_sc_hd__a31o_1 _0870_ (.A1(_0219_),
    .A2(_0222_),
    .A3(_0223_),
    .B1(_0185_),
    .X(_0244_));
 sky130_fd_sc_hd__a41o_1 _0871_ (.A1(_0205_),
    .A2(_0165_),
    .A3(_0159_),
    .A4(_0244_),
    .B1(_0214_),
    .X(_0245_));
 sky130_fd_sc_hd__nor2_1 _0872_ (.A(_0167_),
    .B(_0195_),
    .Y(_0246_));
 sky130_fd_sc_hd__a211oi_1 _0873_ (.A1(_0241_),
    .A2(_0243_),
    .B1(_0245_),
    .C1(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__a21boi_1 _0874_ (.A1(_0165_),
    .A2(_0244_),
    .B1_N(_0195_),
    .Y(_0248_));
 sky130_fd_sc_hd__a21oi_2 _0875_ (.A1(_0209_),
    .A2(_0210_),
    .B1(_0165_),
    .Y(_0249_));
 sky130_fd_sc_hd__and4_1 _0876_ (.A(_0154_),
    .B(_0155_),
    .C(_0196_),
    .D(\SS_FSM.count[2] ),
    .X(_0250_));
 sky130_fd_sc_hd__o21ai_1 _0877_ (.A1(_0249_),
    .A2(_0250_),
    .B1(_0228_),
    .Y(_0251_));
 sky130_fd_sc_hd__o211a_1 _0878_ (.A1(_0228_),
    .A2(_0248_),
    .B1(_0251_),
    .C1(_0178_),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _0879_ (.A(\SS_FSM.count[3] ),
    .B(_0162_),
    .Y(_0253_));
 sky130_fd_sc_hd__o311a_1 _0880_ (.A1(_0184_),
    .A2(\SS_FSM.count[5] ),
    .A3(_0253_),
    .B1(_0198_),
    .C1(_0224_),
    .X(_0254_));
 sky130_fd_sc_hd__a21oi_1 _0881_ (.A1(_0224_),
    .A2(_0198_),
    .B1(_0165_),
    .Y(_0255_));
 sky130_fd_sc_hd__a211o_1 _0882_ (.A1(_0155_),
    .A2(_0196_),
    .B1(\SS_FSM.count[2] ),
    .C1(_0179_),
    .X(_0256_));
 sky130_fd_sc_hd__o21a_1 _0883_ (.A1(_0228_),
    .A2(_0256_),
    .B1(_0159_),
    .X(_0257_));
 sky130_fd_sc_hd__o31a_1 _0884_ (.A1(_0167_),
    .A2(_0254_),
    .A3(_0255_),
    .B1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__o21a_1 _0885_ (.A1(_0252_),
    .A2(_0258_),
    .B1(_0214_),
    .X(_0259_));
 sky130_fd_sc_hd__o21a_1 _0886_ (.A1(_0247_),
    .A2(_0259_),
    .B1(_0217_),
    .X(_0260_));
 sky130_fd_sc_hd__nor2_1 _0887_ (.A(_0179_),
    .B(_0183_),
    .Y(_0261_));
 sky130_fd_sc_hd__or2_1 _0888_ (.A(_0162_),
    .B(_0183_),
    .X(_0262_));
 sky130_fd_sc_hd__a221o_1 _0889_ (.A1(_0219_),
    .A2(_0261_),
    .B1(_0262_),
    .B2(_0210_),
    .C1(_0189_),
    .X(_0263_));
 sky130_fd_sc_hd__nor2_1 _0890_ (.A(_0166_),
    .B(_0249_),
    .Y(_0264_));
 sky130_fd_sc_hd__a32o_1 _0891_ (.A1(_0167_),
    .A2(_0195_),
    .A3(_0263_),
    .B1(_0264_),
    .B2(_0225_),
    .X(_0265_));
 sky130_fd_sc_hd__o2111a_1 _0892_ (.A1(_0184_),
    .A2(\SS_FSM.count[2] ),
    .B1(_0166_),
    .C1(_0196_),
    .D1(_0154_),
    .X(_0266_));
 sky130_fd_sc_hd__a311oi_1 _0893_ (.A1(_0228_),
    .A2(_0261_),
    .A3(_0253_),
    .B1(_0266_),
    .C1(_0178_),
    .Y(_0267_));
 sky130_fd_sc_hd__a211o_1 _0894_ (.A1(_0178_),
    .A2(_0265_),
    .B1(_0267_),
    .C1(_0176_),
    .X(_0268_));
 sky130_fd_sc_hd__or2_2 _0895_ (.A(\SS_FSM.count[3] ),
    .B(_0190_),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_1 _0896_ (.A(_0154_),
    .B(\SS_FSM.count[5] ),
    .Y(_0270_));
 sky130_fd_sc_hd__a2111o_1 _0897_ (.A1(_0167_),
    .A2(_0269_),
    .B1(_0270_),
    .C1(_0264_),
    .D1(_0214_),
    .X(_0271_));
 sky130_fd_sc_hd__a31o_1 _0898_ (.A1(_0232_),
    .A2(_0268_),
    .A3(_0271_),
    .B1(_0175_),
    .X(_0272_));
 sky130_fd_sc_hd__o21a_1 _0899_ (.A1(_0260_),
    .A2(_0272_),
    .B1(_0238_),
    .X(_0273_));
 sky130_fd_sc_hd__a311o_2 _0900_ (.A1(_0155_),
    .A2(_0159_),
    .A3(_0168_),
    .B1(_0273_),
    .C1(_0240_),
    .X(net20));
 sky130_fd_sc_hd__nor2_1 _0901_ (.A(_0240_),
    .B(\SS_FSM.sound[1] ),
    .Y(_0274_));
 sky130_fd_sc_hd__or3_1 _0902_ (.A(_0179_),
    .B(_0184_),
    .C(\SS_FSM.count[3] ),
    .X(_0275_));
 sky130_fd_sc_hd__o31a_1 _0903_ (.A1(_0179_),
    .A2(_0165_),
    .A3(_0186_),
    .B1(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__o21a_1 _0904_ (.A1(_0206_),
    .A2(_0191_),
    .B1(_0156_),
    .X(_0277_));
 sky130_fd_sc_hd__nor2_1 _0905_ (.A(\SS_FSM.count[4] ),
    .B(_0156_),
    .Y(_0278_));
 sky130_fd_sc_hd__o22a_1 _0906_ (.A1(_0167_),
    .A2(_0276_),
    .B1(_0277_),
    .B2(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__o211a_1 _0907_ (.A1(_0189_),
    .A2(_0229_),
    .B1(_0228_),
    .C1(_0209_),
    .X(_0280_));
 sky130_fd_sc_hd__a311o_1 _0908_ (.A1(_0167_),
    .A2(_0187_),
    .A3(_0192_),
    .B1(_0280_),
    .C1(_0159_),
    .X(_0281_));
 sky130_fd_sc_hd__o211ai_1 _0909_ (.A1(_0178_),
    .A2(_0279_),
    .B1(_0281_),
    .C1(_0214_),
    .Y(_0282_));
 sky130_fd_sc_hd__or4_1 _0910_ (.A(_0179_),
    .B(_0165_),
    .C(_0166_),
    .D(_0186_),
    .X(_0283_));
 sky130_fd_sc_hd__a21oi_1 _0911_ (.A1(_0211_),
    .A2(_0283_),
    .B1(_0178_),
    .Y(_0284_));
 sky130_fd_sc_hd__o311a_1 _0912_ (.A1(_0179_),
    .A2(_0193_),
    .A3(_0228_),
    .B1(_0269_),
    .C1(_0209_),
    .X(_0285_));
 sky130_fd_sc_hd__nor2_1 _0913_ (.A(_0159_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__o31a_1 _0914_ (.A1(_0214_),
    .A2(_0284_),
    .A3(_0286_),
    .B1(_0232_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_1 _0915_ (.A(_0189_),
    .B(_0198_),
    .X(_0288_));
 sky130_fd_sc_hd__a31o_1 _0916_ (.A1(_0195_),
    .A2(_0197_),
    .A3(_0288_),
    .B1(_0167_),
    .X(_0289_));
 sky130_fd_sc_hd__a21oi_1 _0917_ (.A1(_0202_),
    .A2(_0289_),
    .B1(_0178_),
    .Y(_0290_));
 sky130_fd_sc_hd__o211a_1 _0918_ (.A1(_0249_),
    .A2(_0250_),
    .B1(\SS_FSM.count[5] ),
    .C1(_0167_),
    .X(_0291_));
 sky130_fd_sc_hd__a211o_1 _0919_ (.A1(_0179_),
    .A2(\SS_FSM.count[2] ),
    .B1(_0196_),
    .C1(_0155_),
    .X(_0292_));
 sky130_fd_sc_hd__a21oi_1 _0920_ (.A1(_0195_),
    .A2(_0292_),
    .B1(_0167_),
    .Y(_0293_));
 sky130_fd_sc_hd__a211o_1 _0921_ (.A1(_0178_),
    .A2(_0207_),
    .B1(_0245_),
    .C1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__o311a_1 _0922_ (.A1(_0176_),
    .A2(_0290_),
    .A3(_0291_),
    .B1(_0294_),
    .C1(_0217_),
    .X(_0295_));
 sky130_fd_sc_hd__a21oi_1 _0923_ (.A1(_0282_),
    .A2(_0287_),
    .B1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__o31ai_4 _0924_ (.A1(\SS_FSM.count[3] ),
    .A2(\SS_FSM.count[2] ),
    .A3(_0234_),
    .B1(_0175_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21ai_4 _0925_ (.A1(_0175_),
    .A2(_0296_),
    .B1(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_2 _0926_ (.A(_0240_),
    .B(_0236_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _0927_ (.A(_0179_),
    .B(_0184_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _0928_ (.A(_0185_),
    .B(_0270_),
    .Y(_0301_));
 sky130_fd_sc_hd__or2_1 _0929_ (.A(_0178_),
    .B(_0300_),
    .X(_0302_));
 sky130_fd_sc_hd__or3b_1 _0930_ (.A(\SS_FSM.count[5] ),
    .B(_0162_),
    .C_N(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__a221o_1 _0931_ (.A1(_0189_),
    .A2(_0300_),
    .B1(_0301_),
    .B2(_0303_),
    .C1(_0228_),
    .X(_0304_));
 sky130_fd_sc_hd__a22oi_4 _0932_ (.A1(_0274_),
    .A2(_0298_),
    .B1(_0299_),
    .B2(_0304_),
    .Y(net21));
 sky130_fd_sc_hd__o21ai_1 _0933_ (.A1(_0242_),
    .A2(_0246_),
    .B1(_0178_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21ai_1 _0934_ (.A1(_0165_),
    .A2(_0229_),
    .B1(_0212_),
    .Y(_0306_));
 sky130_fd_sc_hd__or4_1 _0935_ (.A(_0179_),
    .B(_0162_),
    .C(_0228_),
    .D(_0183_),
    .X(_0307_));
 sky130_fd_sc_hd__o211a_1 _0936_ (.A1(_0165_),
    .A2(_0229_),
    .B1(_0212_),
    .C1(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__a211o_1 _0937_ (.A1(_0167_),
    .A2(_0306_),
    .B1(_0308_),
    .C1(_0178_),
    .X(_0309_));
 sky130_fd_sc_hd__a21o_1 _0938_ (.A1(_0305_),
    .A2(_0309_),
    .B1(_0214_),
    .X(_0310_));
 sky130_fd_sc_hd__o21a_1 _0939_ (.A1(_0189_),
    .A2(_0186_),
    .B1(_0178_),
    .X(_0311_));
 sky130_fd_sc_hd__a221o_1 _0940_ (.A1(_0201_),
    .A2(_0257_),
    .B1(_0311_),
    .B2(_0187_),
    .C1(_0176_),
    .X(_0312_));
 sky130_fd_sc_hd__a211o_1 _0941_ (.A1(_0310_),
    .A2(_0312_),
    .B1(_0175_),
    .C1(_0232_),
    .X(_0313_));
 sky130_fd_sc_hd__nor2_1 _0942_ (.A(_0228_),
    .B(_0248_),
    .Y(_0314_));
 sky130_fd_sc_hd__a21oi_1 _0943_ (.A1(_0210_),
    .A2(_0262_),
    .B1(_0189_),
    .Y(_0315_));
 sky130_fd_sc_hd__o21a_1 _0944_ (.A1(_0249_),
    .A2(_0315_),
    .B1(_0228_),
    .X(_0316_));
 sky130_fd_sc_hd__o21a_1 _0945_ (.A1(_0189_),
    .A2(_0186_),
    .B1(_0205_),
    .X(_0317_));
 sky130_fd_sc_hd__o21a_1 _0946_ (.A1(_0205_),
    .A2(_0288_),
    .B1(_0228_),
    .X(_0318_));
 sky130_fd_sc_hd__o211a_1 _0947_ (.A1(_0167_),
    .A2(_0195_),
    .B1(_0213_),
    .C1(_0159_),
    .X(_0319_));
 sky130_fd_sc_hd__o21ai_1 _0948_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__o311a_1 _0949_ (.A1(_0159_),
    .A2(_0314_),
    .A3(_0316_),
    .B1(_0320_),
    .C1(_0214_),
    .X(_0321_));
 sky130_fd_sc_hd__inv_2 _0950_ (.A(_0190_),
    .Y(_0322_));
 sky130_fd_sc_hd__o21ai_1 _0951_ (.A1(_0322_),
    .A2(_0250_),
    .B1(_0167_),
    .Y(_0323_));
 sky130_fd_sc_hd__a21oi_1 _0952_ (.A1(_0230_),
    .A2(_0323_),
    .B1(_0159_),
    .Y(_0324_));
 sky130_fd_sc_hd__o21a_1 _0953_ (.A1(_0284_),
    .A2(_0324_),
    .B1(_0176_),
    .X(_0325_));
 sky130_fd_sc_hd__o21ai_1 _0954_ (.A1(_0321_),
    .A2(_0325_),
    .B1(_0232_),
    .Y(_0326_));
 sky130_fd_sc_hd__a31o_1 _0955_ (.A1(_0297_),
    .A2(_0313_),
    .A3(_0326_),
    .B1(_0237_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(\SS_FSM.count[5] ),
    .A1(_0302_),
    .S(_0219_),
    .X(_0328_));
 sky130_fd_sc_hd__o21ai_1 _0957_ (.A1(_0206_),
    .A2(_0328_),
    .B1(_0299_),
    .Y(_0329_));
 sky130_fd_sc_hd__and2_1 _0958_ (.A(_0327_),
    .B(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _0959_ (.A(_0330_),
    .X(net22));
 sky130_fd_sc_hd__buf_4 _0960_ (.A(net1),
    .X(_0331_));
 sky130_fd_sc_hd__or4_2 _0961_ (.A(\kp_encoder.sync_out[0] ),
    .B(\kp_encoder.sync_out[1] ),
    .C(\kp_encoder.sync_out[2] ),
    .D(\kp_encoder.sync_out[3] ),
    .X(_0332_));
 sky130_fd_sc_hd__or4_1 _0962_ (.A(\kp_encoder.sync_out[4] ),
    .B(\kp_encoder.sync_out[5] ),
    .C(\kp_encoder.sync_out[6] ),
    .D(\kp_encoder.sync_out[7] ),
    .X(_0333_));
 sky130_fd_sc_hd__or2_1 _0963_ (.A(_0332_),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__or4_1 _0964_ (.A(\kp_encoder.sync_out[8] ),
    .B(\kp_encoder.sync_out[9] ),
    .C(\kp_encoder.sync_out[10] ),
    .D(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__or3b_1 _0965_ (.A(_0335_),
    .B(\kp_encoder.sync_out[11] ),
    .C_N(\kp_encoder.sync_out[12] ),
    .X(_0336_));
 sky130_fd_sc_hd__nor2_1 _0966_ (.A(\kp_encoder.sync_out[8] ),
    .B(_0334_),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(\kp_encoder.sync_out[10] ),
    .Y(_0338_));
 sky130_fd_sc_hd__or3b_1 _0968_ (.A(\kp_encoder.sync_out[4] ),
    .B(\kp_encoder.sync_out[5] ),
    .C_N(\kp_encoder.sync_out[6] ),
    .X(_0339_));
 sky130_fd_sc_hd__o221a_1 _0969_ (.A1(\kp_encoder.sync_out[9] ),
    .A2(_0338_),
    .B1(_0332_),
    .B2(_0339_),
    .C1(_0337_),
    .X(_0340_));
 sky130_fd_sc_hd__nand2_1 _0970_ (.A(_0340_),
    .B(_0336_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(\kp_encoder.sync_out[11] ),
    .Y(_0342_));
 sky130_fd_sc_hd__nor2_1 _0972_ (.A(_0342_),
    .B(_0335_),
    .Y(_0343_));
 sky130_fd_sc_hd__a211o_2 _0973_ (.A1(\kp_encoder.sync_out[9] ),
    .A2(_0337_),
    .B1(_0341_),
    .C1(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__nand3_1 _0974_ (.A(_0297_),
    .B(_0313_),
    .C(_0326_),
    .Y(_0345_));
 sky130_fd_sc_hd__o31ai_4 _0975_ (.A1(\SS_FSM.sound[1] ),
    .A2(_0298_),
    .A3(_0345_),
    .B1(\SS_FSM.sound[0] ),
    .Y(_0346_));
 sky130_fd_sc_hd__or2b_1 _0976_ (.A(_0332_),
    .B_N(_0333_),
    .X(_0347_));
 sky130_fd_sc_hd__nand4_2 _0977_ (.A(_0336_),
    .B(_0344_),
    .C(_0346_),
    .D(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__or2_1 _0978_ (.A(net21),
    .B(_0344_),
    .X(_0349_));
 sky130_fd_sc_hd__clkinv_8 _0979_ (.A(net1),
    .Y(_0350_));
 sky130_fd_sc_hd__a21o_1 _0980_ (.A1(_0348_),
    .A2(_0349_),
    .B1(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_2 _0981_ (.A(_0344_),
    .B(_0346_),
    .Y(_0352_));
 sky130_fd_sc_hd__or3_1 _0982_ (.A(net20),
    .B(_0344_),
    .C(_0346_),
    .X(_0353_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(\kp_encoder.sync_out[9] ),
    .Y(_0354_));
 sky130_fd_sc_hd__nor2_1 _0984_ (.A(\kp_encoder.sync_out[2] ),
    .B(\kp_encoder.sync_out[3] ),
    .Y(_0355_));
 sky130_fd_sc_hd__or4b_1 _0985_ (.A(\kp_encoder.sync_out[4] ),
    .B(\kp_encoder.sync_out[5] ),
    .C(\kp_encoder.sync_out[6] ),
    .D_N(\kp_encoder.sync_out[7] ),
    .X(_0356_));
 sky130_fd_sc_hd__a311oi_1 _0986_ (.A1(_0355_),
    .A2(_0339_),
    .A3(_0356_),
    .B1(\kp_encoder.sync_out[1] ),
    .C1(\kp_encoder.sync_out[0] ),
    .Y(_0357_));
 sky130_fd_sc_hd__a311o_1 _0987_ (.A1(_0354_),
    .A2(\kp_encoder.sync_out[10] ),
    .A3(_0337_),
    .B1(_0343_),
    .C1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__a31o_1 _0988_ (.A1(_0344_),
    .A2(_0346_),
    .A3(_0358_),
    .B1(_0350_),
    .X(_0359_));
 sky130_fd_sc_hd__a21o_1 _0989_ (.A1(_0352_),
    .A2(_0353_),
    .B1(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_4 _0990_ (.A(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__or3_2 _0991_ (.A(net19),
    .B(_0344_),
    .C(_0346_),
    .X(_0362_));
 sky130_fd_sc_hd__inv_2 _0992_ (.A(\kp_encoder.sync_out[5] ),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(\kp_encoder.sync_out[2] ),
    .Y(_0364_));
 sky130_fd_sc_hd__a21oi_1 _0994_ (.A1(_0364_),
    .A2(\kp_encoder.sync_out[3] ),
    .B1(\kp_encoder.sync_out[1] ),
    .Y(_0365_));
 sky130_fd_sc_hd__o32a_1 _0995_ (.A1(\kp_encoder.sync_out[4] ),
    .A2(_0363_),
    .A3(_0332_),
    .B1(_0365_),
    .B2(\kp_encoder.sync_out[0] ),
    .X(_0366_));
 sky130_fd_sc_hd__o21ai_1 _0996_ (.A1(_0332_),
    .A2(_0356_),
    .B1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__a211o_1 _0997_ (.A1(\kp_encoder.sync_out[9] ),
    .A2(_0337_),
    .B1(_0343_),
    .C1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__a31o_1 _0998_ (.A1(_0344_),
    .A2(_0346_),
    .A3(_0368_),
    .B1(_0350_),
    .X(_0369_));
 sky130_fd_sc_hd__a21oi_4 _0999_ (.A1(_0352_),
    .A2(_0362_),
    .B1(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a21oi_1 _1000_ (.A1(_0327_),
    .A2(_0329_),
    .B1(_0344_),
    .Y(_0371_));
 sky130_fd_sc_hd__a31o_1 _1001_ (.A1(_0334_),
    .A2(_0344_),
    .A3(_0346_),
    .B1(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__and2_2 _1002_ (.A(net1),
    .B(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__o31ai_1 _1003_ (.A1(_0351_),
    .A2(_0361_),
    .A3(_0370_),
    .B1(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__a21oi_4 _1004_ (.A1(_0348_),
    .A2(_0349_),
    .B1(_0350_),
    .Y(_0375_));
 sky130_fd_sc_hd__nor2_1 _1005_ (.A(_0375_),
    .B(_0361_),
    .Y(_0376_));
 sky130_fd_sc_hd__a21o_2 _1006_ (.A1(_0352_),
    .A2(_0362_),
    .B1(_0369_),
    .X(_0377_));
 sky130_fd_sc_hd__nor2_2 _1007_ (.A(_0361_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__a21o_1 _1008_ (.A1(_0361_),
    .A2(_0377_),
    .B1(_0351_),
    .X(_0379_));
 sky130_fd_sc_hd__or3_1 _1009_ (.A(_0373_),
    .B(_0361_),
    .C(_0377_),
    .X(_0380_));
 sky130_fd_sc_hd__buf_2 _1010_ (.A(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_4 _1011_ (.A(net1),
    .B(_0372_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_2 _1012_ (.A(_0382_),
    .B(_0375_),
    .Y(_0383_));
 sky130_fd_sc_hd__a2bb2o_1 _1013_ (.A1_N(_0378_),
    .A2_N(_0379_),
    .B1(_0381_),
    .B2(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__o21a_1 _1014_ (.A1(_0374_),
    .A2(_0376_),
    .B1(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_2 _1015_ (.A(_0373_),
    .B(_0361_),
    .Y(_0386_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(_0375_),
    .A1(_0379_),
    .S(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _1017_ (.A1(\osc.count[12] ),
    .A2(_0385_),
    .B1(_0387_),
    .B2(\osc.count[13] ),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_1 _1018_ (.A(\osc.count[12] ),
    .B(_0385_),
    .Y(_0389_));
 sky130_fd_sc_hd__nor2_1 _1019_ (.A(_0375_),
    .B(_0370_),
    .Y(_0390_));
 sky130_fd_sc_hd__xnor2_2 _1020_ (.A(_0361_),
    .B(_0377_),
    .Y(_0391_));
 sky130_fd_sc_hd__a21o_1 _1021_ (.A1(_0375_),
    .A2(_0391_),
    .B1(_0382_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _1022_ (.A(_0375_),
    .B(_0381_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _1023_ (.A(_0370_),
    .B(_0383_),
    .X(_0394_));
 sky130_fd_sc_hd__o211a_1 _1024_ (.A1(_0390_),
    .A2(_0392_),
    .B1(_0393_),
    .C1(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__nor2_1 _1025_ (.A(\osc.count[11] ),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__and2_1 _1026_ (.A(_0351_),
    .B(_0361_),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _1027_ (.A(_0382_),
    .B(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_1 _1028_ (.A(\osc.count[15] ),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _1029_ (.A(\osc.count[15] ),
    .B(_0398_),
    .Y(_0400_));
 sky130_fd_sc_hd__or2_1 _1030_ (.A(\osc.count[13] ),
    .B(_0387_),
    .X(_0401_));
 sky130_fd_sc_hd__o211ai_4 _1031_ (.A1(_0375_),
    .A2(_0386_),
    .B1(_0381_),
    .C1(_0383_),
    .Y(_0402_));
 sky130_fd_sc_hd__xnor2_1 _1032_ (.A(\osc.count[14] ),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__and4b_1 _1033_ (.A_N(_0399_),
    .B(_0400_),
    .C(_0401_),
    .D(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__or4b_2 _1034_ (.A(_0388_),
    .B(_0389_),
    .C(_0396_),
    .D_N(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__nand3_2 _1035_ (.A(_0351_),
    .B(_0361_),
    .C(_0377_),
    .Y(_0406_));
 sky130_fd_sc_hd__a21o_1 _1036_ (.A1(_0379_),
    .A2(_0406_),
    .B1(_0382_),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _1037_ (.A(_0374_),
    .B(_0394_),
    .X(_0408_));
 sky130_fd_sc_hd__a32o_1 _1038_ (.A1(\osc.count[8] ),
    .A2(_0393_),
    .A3(_0407_),
    .B1(_0408_),
    .B2(\osc.count[9] ),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _1039_ (.A(_0375_),
    .B(_0361_),
    .Y(_0410_));
 sky130_fd_sc_hd__o21a_1 _1040_ (.A1(_0382_),
    .A2(_0375_),
    .B1(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__o22a_1 _1041_ (.A1(\osc.count[9] ),
    .A2(_0408_),
    .B1(_0411_),
    .B2(\osc.count[10] ),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _1042_ (.A1(\osc.count[11] ),
    .A2(_0395_),
    .B1(_0411_),
    .B2(\osc.count[10] ),
    .X(_0413_));
 sky130_fd_sc_hd__a21oi_1 _1043_ (.A1(_0409_),
    .A2(_0412_),
    .B1(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__nand2_1 _1044_ (.A(_0388_),
    .B(_0404_),
    .Y(_0415_));
 sky130_fd_sc_hd__or3b_1 _1045_ (.A(_0399_),
    .B(_0402_),
    .C_N(\osc.count[14] ),
    .X(_0416_));
 sky130_fd_sc_hd__o2111a_4 _1046_ (.A1(_0405_),
    .A2(_0414_),
    .B1(_0415_),
    .C1(_0416_),
    .D1(_0400_),
    .X(_0417_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(\osc.count[7] ),
    .Y(_0418_));
 sky130_fd_sc_hd__nand3_2 _1048_ (.A(_0383_),
    .B(_0381_),
    .C(_0386_),
    .Y(_0419_));
 sky130_fd_sc_hd__o31a_2 _1049_ (.A1(_0382_),
    .A2(_0361_),
    .A3(_0370_),
    .B1(_0351_),
    .X(_0420_));
 sky130_fd_sc_hd__a21o_1 _1050_ (.A1(_0375_),
    .A2(_0361_),
    .B1(_0382_),
    .X(_0421_));
 sky130_fd_sc_hd__a2bb2o_1 _1051_ (.A1_N(_0375_),
    .A2_N(_0391_),
    .B1(_0421_),
    .B2(_0377_),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_1 _1052_ (.A1(\osc.count[3] ),
    .A2(_0420_),
    .B1(_0422_),
    .B2(\osc.count[2] ),
    .X(_0423_));
 sky130_fd_sc_hd__o21ai_1 _1053_ (.A1(\osc.count[3] ),
    .A2(_0420_),
    .B1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__o21ai_1 _1054_ (.A1(_0361_),
    .A2(_0370_),
    .B1(_0382_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(_0361_),
    .B(_0370_),
    .Y(_0426_));
 sky130_fd_sc_hd__a31o_1 _1056_ (.A1(_0375_),
    .A2(_0425_),
    .A3(_0426_),
    .B1(_0420_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _1057_ (.A(\osc.count[1] ),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__and2_1 _1058_ (.A(_0361_),
    .B(_0377_),
    .X(_0429_));
 sky130_fd_sc_hd__o22ai_2 _1059_ (.A1(_0383_),
    .A2(_0378_),
    .B1(_0429_),
    .B2(_0382_),
    .Y(_0430_));
 sky130_fd_sc_hd__o22ai_1 _1060_ (.A1(\osc.count[1] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\osc.count[0] ),
    .Y(_0431_));
 sky130_fd_sc_hd__o22ai_1 _1061_ (.A1(\osc.count[3] ),
    .A2(_0420_),
    .B1(_0422_),
    .B2(\osc.count[2] ),
    .Y(_0432_));
 sky130_fd_sc_hd__a211o_1 _1062_ (.A1(_0428_),
    .A2(_0431_),
    .B1(_0432_),
    .C1(_0423_),
    .X(_0433_));
 sky130_fd_sc_hd__a21oi_1 _1063_ (.A1(_0381_),
    .A2(_0392_),
    .B1(\osc.count[4] ),
    .Y(_0434_));
 sky130_fd_sc_hd__o221ai_4 _1064_ (.A1(_0373_),
    .A2(_0429_),
    .B1(_0379_),
    .B2(_0378_),
    .C1(_0406_),
    .Y(_0435_));
 sky130_fd_sc_hd__a32o_1 _1065_ (.A1(\osc.count[4] ),
    .A2(_0381_),
    .A3(_0392_),
    .B1(_0435_),
    .B2(\osc.count[5] ),
    .X(_0436_));
 sky130_fd_sc_hd__nand2_1 _1066_ (.A(_0375_),
    .B(_0391_),
    .Y(_0437_));
 sky130_fd_sc_hd__o32a_1 _1067_ (.A1(\osc.count[6] ),
    .A2(_0373_),
    .A3(_0437_),
    .B1(_0435_),
    .B2(\osc.count[5] ),
    .X(_0438_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(\osc.count[6] ),
    .Y(_0439_));
 sky130_fd_sc_hd__a31o_1 _1069_ (.A1(_0382_),
    .A2(_0375_),
    .A3(_0391_),
    .B1(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__o21a_1 _1070_ (.A1(_0418_),
    .A2(_0419_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__or4bb_1 _1071_ (.A(_0434_),
    .B(_0436_),
    .C_N(_0438_),
    .D_N(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a221o_1 _1072_ (.A1(_0418_),
    .A2(_0419_),
    .B1(_0424_),
    .B2(_0433_),
    .C1(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _1073_ (.A(_0438_),
    .B(_0436_),
    .Y(_0444_));
 sky130_fd_sc_hd__a22o_1 _1074_ (.A1(_0418_),
    .A2(_0419_),
    .B1(_0441_),
    .B2(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__a21oi_1 _1075_ (.A1(_0393_),
    .A2(_0407_),
    .B1(\osc.count[8] ),
    .Y(_0446_));
 sky130_fd_sc_hd__or3b_1 _1076_ (.A(_0409_),
    .B(_0446_),
    .C_N(_0412_),
    .X(_0447_));
 sky130_fd_sc_hd__a2111o_4 _1077_ (.A1(_0443_),
    .A2(_0445_),
    .B1(_0405_),
    .C1(_0413_),
    .D1(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__nand4_1 _1078_ (.A(_0331_),
    .B(net97),
    .C(_0417_),
    .D(_0448_),
    .Y(\osc.next_count[0] ));
 sky130_fd_sc_hd__nand2_1 _1079_ (.A(\osc.count[0] ),
    .B(\osc.count[1] ),
    .Y(_0449_));
 sky130_fd_sc_hd__or2_1 _1080_ (.A(\osc.count[0] ),
    .B(\osc.count[1] ),
    .X(_0450_));
 sky130_fd_sc_hd__and4_1 _1081_ (.A(_0417_),
    .B(_0448_),
    .C(_0449_),
    .D(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _1082_ (.A(_0451_),
    .X(\osc.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1083_ (.A(\osc.count[0] ),
    .B(\osc.count[2] ),
    .C(\osc.count[1] ),
    .X(_0452_));
 sky130_fd_sc_hd__a21o_1 _1084_ (.A1(\osc.count[0] ),
    .A2(\osc.count[1] ),
    .B1(\osc.count[2] ),
    .X(_0453_));
 sky130_fd_sc_hd__and4b_1 _1085_ (.A_N(_0452_),
    .B(_0417_),
    .C(_0448_),
    .D(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _1086_ (.A(_0454_),
    .X(\osc.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1087_ (.A(\osc.count[3] ),
    .B(_0452_),
    .X(_0455_));
 sky130_fd_sc_hd__or2_1 _1088_ (.A(\osc.count[3] ),
    .B(_0452_),
    .X(_0456_));
 sky130_fd_sc_hd__and4b_1 _1089_ (.A_N(_0455_),
    .B(_0417_),
    .C(_0448_),
    .D(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _1090_ (.A(_0457_),
    .X(\osc.next_count[3] ));
 sky130_fd_sc_hd__and3_1 _1091_ (.A(\osc.count[4] ),
    .B(\osc.count[3] ),
    .C(_0452_),
    .X(_0458_));
 sky130_fd_sc_hd__or2_1 _1092_ (.A(\osc.count[4] ),
    .B(_0455_),
    .X(_0459_));
 sky130_fd_sc_hd__and4b_1 _1093_ (.A_N(_0458_),
    .B(_0417_),
    .C(_0448_),
    .D(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _1094_ (.A(_0460_),
    .X(\osc.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1095_ (.A(\osc.count[5] ),
    .B(\osc.count[4] ),
    .C(_0455_),
    .X(_0461_));
 sky130_fd_sc_hd__or2_1 _1096_ (.A(\osc.count[5] ),
    .B(_0458_),
    .X(_0462_));
 sky130_fd_sc_hd__and4b_1 _1097_ (.A_N(_0461_),
    .B(_0417_),
    .C(_0448_),
    .D(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _1098_ (.A(_0463_),
    .X(\osc.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _1099_ (.A(\osc.count[6] ),
    .B(_0461_),
    .X(_0464_));
 sky130_fd_sc_hd__or2_1 _1100_ (.A(\osc.count[6] ),
    .B(_0461_),
    .X(_0465_));
 sky130_fd_sc_hd__and4b_1 _1101_ (.A_N(_0464_),
    .B(_0417_),
    .C(_0448_),
    .D(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _1102_ (.A(_0466_),
    .X(\osc.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _1103_ (.A(\osc.count[7] ),
    .B(\osc.count[6] ),
    .C(_0461_),
    .X(_0467_));
 sky130_fd_sc_hd__or2_1 _1104_ (.A(\osc.count[7] ),
    .B(_0464_),
    .X(_0468_));
 sky130_fd_sc_hd__and4b_1 _1105_ (.A_N(_0467_),
    .B(_0417_),
    .C(_0448_),
    .D(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _1106_ (.A(_0469_),
    .X(\osc.next_count[7] ));
 sky130_fd_sc_hd__and2_1 _1107_ (.A(\osc.count[8] ),
    .B(_0467_),
    .X(_0470_));
 sky130_fd_sc_hd__or2_1 _1108_ (.A(\osc.count[8] ),
    .B(_0467_),
    .X(_0471_));
 sky130_fd_sc_hd__and4b_1 _1109_ (.A_N(_0470_),
    .B(_0417_),
    .C(_0448_),
    .D(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _1110_ (.A(_0472_),
    .X(\osc.next_count[8] ));
 sky130_fd_sc_hd__and3_1 _1111_ (.A(\osc.count[9] ),
    .B(\osc.count[8] ),
    .C(_0467_),
    .X(_0473_));
 sky130_fd_sc_hd__or2_1 _1112_ (.A(\osc.count[9] ),
    .B(_0470_),
    .X(_0474_));
 sky130_fd_sc_hd__and4b_1 _1113_ (.A_N(_0473_),
    .B(_0417_),
    .C(_0448_),
    .D(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _1114_ (.A(_0475_),
    .X(\osc.next_count[9] ));
 sky130_fd_sc_hd__and2_1 _1115_ (.A(\osc.count[10] ),
    .B(_0473_),
    .X(_0476_));
 sky130_fd_sc_hd__or2_1 _1116_ (.A(\osc.count[10] ),
    .B(_0473_),
    .X(_0477_));
 sky130_fd_sc_hd__and4b_1 _1117_ (.A_N(_0476_),
    .B(_0417_),
    .C(_0448_),
    .D(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _1118_ (.A(_0478_),
    .X(\osc.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _1119_ (.A(\osc.count[11] ),
    .B(\osc.count[10] ),
    .C(_0473_),
    .X(_0479_));
 sky130_fd_sc_hd__or2_1 _1120_ (.A(\osc.count[11] ),
    .B(_0476_),
    .X(_0480_));
 sky130_fd_sc_hd__and4b_1 _1121_ (.A_N(_0479_),
    .B(_0417_),
    .C(_0448_),
    .D(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _1122_ (.A(_0481_),
    .X(\osc.next_count[11] ));
 sky130_fd_sc_hd__and3_1 _1123_ (.A(\osc.count[12] ),
    .B(\osc.count[11] ),
    .C(_0476_),
    .X(_0482_));
 sky130_fd_sc_hd__or2_1 _1124_ (.A(\osc.count[12] ),
    .B(_0479_),
    .X(_0483_));
 sky130_fd_sc_hd__and4b_1 _1125_ (.A_N(_0482_),
    .B(_0417_),
    .C(_0448_),
    .D(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _1126_ (.A(_0484_),
    .X(\osc.next_count[12] ));
 sky130_fd_sc_hd__and2_1 _1127_ (.A(\osc.count[13] ),
    .B(_0482_),
    .X(_0485_));
 sky130_fd_sc_hd__or2_1 _1128_ (.A(\osc.count[13] ),
    .B(_0482_),
    .X(_0486_));
 sky130_fd_sc_hd__and4b_1 _1129_ (.A_N(_0485_),
    .B(_0417_),
    .C(_0448_),
    .D(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _1130_ (.A(_0487_),
    .X(\osc.next_count[13] ));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(\osc.count[14] ),
    .B(_0485_),
    .Y(_0488_));
 sky130_fd_sc_hd__or2_1 _1132_ (.A(\osc.count[14] ),
    .B(_0485_),
    .X(_0489_));
 sky130_fd_sc_hd__and4_1 _1133_ (.A(_0417_),
    .B(_0448_),
    .C(_0488_),
    .D(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _1134_ (.A(_0490_),
    .X(\osc.next_count[14] ));
 sky130_fd_sc_hd__xnor2_1 _1135_ (.A(\osc.count[15] ),
    .B(_0488_),
    .Y(_0491_));
 sky130_fd_sc_hd__and4_1 _1136_ (.A(_0331_),
    .B(_0417_),
    .C(_0448_),
    .D(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _1137_ (.A(_0492_),
    .X(\osc.next_count[15] ));
 sky130_fd_sc_hd__nor2_1 _1138_ (.A(_0350_),
    .B(net64),
    .Y(\clk_div.next_count[0] ));
 sky130_fd_sc_hd__a21oi_1 _1139_ (.A1(net94),
    .A2(\clk_div.count[0] ),
    .B1(_0350_),
    .Y(_0493_));
 sky130_fd_sc_hd__o21a_1 _1140_ (.A1(net94),
    .A2(net64),
    .B1(_0493_),
    .X(\clk_div.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1141_ (.A(\clk_div.count[1] ),
    .B(\clk_div.count[0] ),
    .C(\clk_div.count[2] ),
    .X(_0494_));
 sky130_fd_sc_hd__a21o_1 _1142_ (.A1(\clk_div.count[1] ),
    .A2(\clk_div.count[0] ),
    .B1(\clk_div.count[2] ),
    .X(_0495_));
 sky130_fd_sc_hd__and3b_1 _1143_ (.A_N(_0494_),
    .B(_0331_),
    .C(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _1144_ (.A(_0496_),
    .X(\clk_div.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1145_ (.A(\clk_div.count[3] ),
    .B(_0494_),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_1 _1146_ (.A(_0350_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__o21a_1 _1147_ (.A1(net70),
    .A2(_0494_),
    .B1(_0498_),
    .X(\clk_div.next_count[3] ));
 sky130_fd_sc_hd__a21oi_1 _1148_ (.A1(net93),
    .A2(_0497_),
    .B1(_0350_),
    .Y(_0499_));
 sky130_fd_sc_hd__o21a_1 _1149_ (.A1(net93),
    .A2(_0497_),
    .B1(_0499_),
    .X(\clk_div.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1150_ (.A(\clk_div.count[5] ),
    .B(\clk_div.count[4] ),
    .C(_0497_),
    .X(_0500_));
 sky130_fd_sc_hd__a31o_1 _1151_ (.A1(\clk_div.count[3] ),
    .A2(\clk_div.count[4] ),
    .A3(_0494_),
    .B1(\clk_div.count[5] ),
    .X(_0501_));
 sky130_fd_sc_hd__and3b_1 _1152_ (.A_N(_0500_),
    .B(_0331_),
    .C(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _1153_ (.A(_0502_),
    .X(\clk_div.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _1154_ (.A(\clk_div.count[6] ),
    .B(_0500_),
    .X(_0503_));
 sky130_fd_sc_hd__or2_1 _1155_ (.A(\clk_div.count[6] ),
    .B(_0500_),
    .X(_0504_));
 sky130_fd_sc_hd__and3b_1 _1156_ (.A_N(_0503_),
    .B(_0331_),
    .C(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _1157_ (.A(_0505_),
    .X(\clk_div.next_count[6] ));
 sky130_fd_sc_hd__or2_1 _1158_ (.A(\clk_div.count[7] ),
    .B(_0503_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_2 _1159_ (.A(\clk_div.count[7] ),
    .B(_0503_),
    .Y(_0507_));
 sky130_fd_sc_hd__and3_1 _1160_ (.A(_0331_),
    .B(_0506_),
    .C(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _1161_ (.A(_0508_),
    .X(\clk_div.next_count[7] ));
 sky130_fd_sc_hd__nor2_1 _1162_ (.A(_0350_),
    .B(net58),
    .Y(\pwm.next_count[0] ));
 sky130_fd_sc_hd__o21ai_1 _1163_ (.A1(\pwm.count[0] ),
    .A2(net71),
    .B1(_0331_),
    .Y(_0509_));
 sky130_fd_sc_hd__a21oi_1 _1164_ (.A1(net58),
    .A2(net71),
    .B1(_0509_),
    .Y(\pwm.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1165_ (.A(\pwm.count[2] ),
    .B(\pwm.count[0] ),
    .C(\pwm.count[1] ),
    .X(_0510_));
 sky130_fd_sc_hd__a21o_1 _1166_ (.A1(\pwm.count[0] ),
    .A2(\pwm.count[1] ),
    .B1(\pwm.count[2] ),
    .X(_0511_));
 sky130_fd_sc_hd__and3b_1 _1167_ (.A_N(_0510_),
    .B(_0511_),
    .C(_0331_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _1168_ (.A(_0512_),
    .X(\pwm.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1169_ (.A(\pwm.count[3] ),
    .B(_0510_),
    .X(_0513_));
 sky130_fd_sc_hd__o21ai_1 _1170_ (.A1(\pwm.count[3] ),
    .A2(_0510_),
    .B1(_0331_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _1171_ (.A(_0513_),
    .B(_0514_),
    .Y(\pwm.next_count[3] ));
 sky130_fd_sc_hd__a31o_1 _1172_ (.A1(\pwm.count[4] ),
    .A2(\pwm.count[3] ),
    .A3(_0510_),
    .B1(_0350_),
    .X(_0515_));
 sky130_fd_sc_hd__o21ba_1 _1173_ (.A1(\pwm.count[4] ),
    .A2(_0513_),
    .B1_N(_0515_),
    .X(\pwm.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1174_ (.A(\pwm.count[5] ),
    .B(\pwm.count[4] ),
    .C(_0513_),
    .X(_0516_));
 sky130_fd_sc_hd__a31o_1 _1175_ (.A1(\pwm.count[4] ),
    .A2(\pwm.count[3] ),
    .A3(_0510_),
    .B1(\pwm.count[5] ),
    .X(_0517_));
 sky130_fd_sc_hd__and3b_1 _1176_ (.A_N(_0516_),
    .B(_0331_),
    .C(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1177_ (.A(_0518_),
    .X(\pwm.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _1178_ (.A(\pwm.count[6] ),
    .B(_0516_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _1179_ (.A(\pwm.count[6] ),
    .B(_0516_),
    .X(_0520_));
 sky130_fd_sc_hd__and3b_1 _1180_ (.A_N(_0519_),
    .B(_0331_),
    .C(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _1181_ (.A(_0521_),
    .X(\pwm.next_count[6] ));
 sky130_fd_sc_hd__o21ai_1 _1182_ (.A1(net61),
    .A2(_0519_),
    .B1(_0331_),
    .Y(_0522_));
 sky130_fd_sc_hd__a21oi_1 _1183_ (.A1(net61),
    .A2(_0519_),
    .B1(_0522_),
    .Y(\pwm.next_count[7] ));
 sky130_fd_sc_hd__or4b_1 _1184_ (.A(\clk8.count[3] ),
    .B(\clk8.count[2] ),
    .C(\clk8.count[4] ),
    .D_N(\clk8.count[5] ),
    .X(_0523_));
 sky130_fd_sc_hd__or4b_1 _1185_ (.A(\clk8.count[11] ),
    .B(\clk8.count[10] ),
    .C(\clk8.count[12] ),
    .D_N(\clk8.count[13] ),
    .X(_0524_));
 sky130_fd_sc_hd__and4b_1 _1186_ (.A_N(\clk8.count[7] ),
    .B(\clk8.count[6] ),
    .C(\clk8.count[9] ),
    .D(\clk8.count[8] ),
    .X(_0525_));
 sky130_fd_sc_hd__and4b_1 _1187_ (.A_N(\clk8.count[16] ),
    .B(\clk8.count[20] ),
    .C(\clk8.count[14] ),
    .D(\clk8.count[15] ),
    .X(_0526_));
 sky130_fd_sc_hd__and3b_1 _1188_ (.A_N(\clk8.count[19] ),
    .B(\clk8.count[18] ),
    .C(\clk8.count[17] ),
    .X(_0527_));
 sky130_fd_sc_hd__and4b_1 _1189_ (.A_N(_0524_),
    .B(_0525_),
    .C(_0526_),
    .D(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__or4b_1 _1190_ (.A(\clk8.count[1] ),
    .B(\clk8.count[0] ),
    .C(_0523_),
    .D_N(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__and2_1 _1191_ (.A(_0331_),
    .B(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__buf_2 _1192_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__and2b_1 _1193_ (.A_N(\clk8.count[0] ),
    .B(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1194_ (.A(_0532_),
    .X(\clk8.next_count[0] ));
 sky130_fd_sc_hd__o21ai_1 _1195_ (.A1(net65),
    .A2(\clk8.count[0] ),
    .B1(_0331_),
    .Y(_0533_));
 sky130_fd_sc_hd__a21oi_1 _1196_ (.A1(net65),
    .A2(\clk8.count[0] ),
    .B1(_0533_),
    .Y(\clk8.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1197_ (.A(\clk8.count[1] ),
    .B(\clk8.count[0] ),
    .C(\clk8.count[2] ),
    .X(_0534_));
 sky130_fd_sc_hd__a21o_1 _1198_ (.A1(\clk8.count[1] ),
    .A2(\clk8.count[0] ),
    .B1(\clk8.count[2] ),
    .X(_0535_));
 sky130_fd_sc_hd__and3b_1 _1199_ (.A_N(_0534_),
    .B(_0331_),
    .C(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1200_ (.A(_0536_),
    .X(\clk8.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1201_ (.A(\clk8.count[3] ),
    .B(_0534_),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_1 _1202_ (.A(_0350_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__o21a_1 _1203_ (.A1(net90),
    .A2(_0534_),
    .B1(_0538_),
    .X(\clk8.next_count[3] ));
 sky130_fd_sc_hd__a21oi_1 _1204_ (.A1(\clk8.count[4] ),
    .A2(_0537_),
    .B1(_0350_),
    .Y(_0539_));
 sky130_fd_sc_hd__o21a_1 _1205_ (.A1(net103),
    .A2(_0537_),
    .B1(_0539_),
    .X(\clk8.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1206_ (.A(\clk8.count[4] ),
    .B(\clk8.count[5] ),
    .C(_0537_),
    .X(_0540_));
 sky130_fd_sc_hd__a31o_1 _1207_ (.A1(\clk8.count[3] ),
    .A2(\clk8.count[4] ),
    .A3(_0534_),
    .B1(\clk8.count[5] ),
    .X(_0541_));
 sky130_fd_sc_hd__and3b_1 _1208_ (.A_N(_0540_),
    .B(_0541_),
    .C(_0531_),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_1 _1209_ (.A(_0542_),
    .X(\clk8.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _1210_ (.A(\clk8.count[6] ),
    .B(_0540_),
    .X(_0543_));
 sky130_fd_sc_hd__o21ai_1 _1211_ (.A1(\clk8.count[6] ),
    .A2(_0540_),
    .B1(_0531_),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_1 _1212_ (.A(_0543_),
    .B(_0544_),
    .Y(\clk8.next_count[6] ));
 sky130_fd_sc_hd__a31o_1 _1213_ (.A1(\clk8.count[7] ),
    .A2(\clk8.count[6] ),
    .A3(_0540_),
    .B1(_0350_),
    .X(_0545_));
 sky130_fd_sc_hd__o21ba_1 _1214_ (.A1(net106),
    .A2(_0543_),
    .B1_N(_0545_),
    .X(\clk8.next_count[7] ));
 sky130_fd_sc_hd__and3_1 _1215_ (.A(\clk8.count[7] ),
    .B(\clk8.count[8] ),
    .C(_0543_),
    .X(_0546_));
 sky130_fd_sc_hd__a31o_1 _1216_ (.A1(\clk8.count[7] ),
    .A2(\clk8.count[6] ),
    .A3(_0540_),
    .B1(\clk8.count[8] ),
    .X(_0547_));
 sky130_fd_sc_hd__and3b_1 _1217_ (.A_N(_0546_),
    .B(_0531_),
    .C(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_1 _1218_ (.A(_0548_),
    .X(\clk8.next_count[8] ));
 sky130_fd_sc_hd__and2_1 _1219_ (.A(\clk8.count[9] ),
    .B(_0546_),
    .X(_0549_));
 sky130_fd_sc_hd__or2_1 _1220_ (.A(\clk8.count[9] ),
    .B(_0546_),
    .X(_0550_));
 sky130_fd_sc_hd__and3b_1 _1221_ (.A_N(_0549_),
    .B(_0531_),
    .C(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_1 _1222_ (.A(_0551_),
    .X(\clk8.next_count[9] ));
 sky130_fd_sc_hd__a31o_1 _1223_ (.A1(\clk8.count[9] ),
    .A2(\clk8.count[10] ),
    .A3(_0546_),
    .B1(_0350_),
    .X(_0552_));
 sky130_fd_sc_hd__o21ba_1 _1224_ (.A1(net110),
    .A2(_0549_),
    .B1_N(_0552_),
    .X(\clk8.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _1225_ (.A(\clk8.count[11] ),
    .B(\clk8.count[10] ),
    .C(_0549_),
    .X(_0553_));
 sky130_fd_sc_hd__a31o_1 _1226_ (.A1(\clk8.count[9] ),
    .A2(\clk8.count[10] ),
    .A3(_0546_),
    .B1(\clk8.count[11] ),
    .X(_0554_));
 sky130_fd_sc_hd__and3b_1 _1227_ (.A_N(_0553_),
    .B(_0331_),
    .C(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_1 _1228_ (.A(_0555_),
    .X(\clk8.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _1229_ (.A(\clk8.count[12] ),
    .B(_0553_),
    .X(_0556_));
 sky130_fd_sc_hd__or2_1 _1230_ (.A(\clk8.count[12] ),
    .B(_0553_),
    .X(_0557_));
 sky130_fd_sc_hd__and3b_1 _1231_ (.A_N(_0556_),
    .B(_0331_),
    .C(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_1 _1232_ (.A(_0558_),
    .X(\clk8.next_count[12] ));
 sky130_fd_sc_hd__a21boi_1 _1233_ (.A1(\clk8.count[13] ),
    .A2(_0556_),
    .B1_N(_0531_),
    .Y(_0559_));
 sky130_fd_sc_hd__o21a_1 _1234_ (.A1(net101),
    .A2(_0556_),
    .B1(_0559_),
    .X(\clk8.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _1235_ (.A(\clk8.count[13] ),
    .B(\clk8.count[14] ),
    .C(_0556_),
    .X(_0560_));
 sky130_fd_sc_hd__a31o_1 _1236_ (.A1(\clk8.count[12] ),
    .A2(\clk8.count[13] ),
    .A3(_0553_),
    .B1(\clk8.count[14] ),
    .X(_0561_));
 sky130_fd_sc_hd__and3b_1 _1237_ (.A_N(_0560_),
    .B(_0531_),
    .C(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_1 _1238_ (.A(_0562_),
    .X(\clk8.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _1239_ (.A(\clk8.count[15] ),
    .B(_0560_),
    .X(_0563_));
 sky130_fd_sc_hd__or2_1 _1240_ (.A(\clk8.count[15] ),
    .B(_0560_),
    .X(_0564_));
 sky130_fd_sc_hd__and3b_1 _1241_ (.A_N(_0563_),
    .B(_0531_),
    .C(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1242_ (.A(_0565_),
    .X(\clk8.next_count[15] ));
 sky130_fd_sc_hd__a31o_1 _1243_ (.A1(\clk8.count[15] ),
    .A2(\clk8.count[16] ),
    .A3(_0560_),
    .B1(_0350_),
    .X(_0566_));
 sky130_fd_sc_hd__o21ba_1 _1244_ (.A1(net105),
    .A2(_0563_),
    .B1_N(_0566_),
    .X(\clk8.next_count[16] ));
 sky130_fd_sc_hd__and3_1 _1245_ (.A(\clk8.count[16] ),
    .B(\clk8.count[17] ),
    .C(_0563_),
    .X(_0567_));
 sky130_fd_sc_hd__a31o_1 _1246_ (.A1(\clk8.count[15] ),
    .A2(\clk8.count[16] ),
    .A3(_0560_),
    .B1(\clk8.count[17] ),
    .X(_0568_));
 sky130_fd_sc_hd__and3b_1 _1247_ (.A_N(_0567_),
    .B(_0531_),
    .C(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_1 _1248_ (.A(_0569_),
    .X(\clk8.next_count[17] ));
 sky130_fd_sc_hd__and2_1 _1249_ (.A(\clk8.count[18] ),
    .B(_0567_),
    .X(_0570_));
 sky130_fd_sc_hd__or2_1 _1250_ (.A(\clk8.count[18] ),
    .B(_0567_),
    .X(_0571_));
 sky130_fd_sc_hd__and3b_1 _1251_ (.A_N(_0570_),
    .B(_0531_),
    .C(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_1 _1252_ (.A(_0572_),
    .X(\clk8.next_count[18] ));
 sky130_fd_sc_hd__and3_1 _1253_ (.A(\clk8.count[19] ),
    .B(\clk8.count[18] ),
    .C(_0567_),
    .X(_0573_));
 sky130_fd_sc_hd__or2_1 _1254_ (.A(\clk8.count[19] ),
    .B(_0570_),
    .X(_0574_));
 sky130_fd_sc_hd__and3b_1 _1255_ (.A_N(_0573_),
    .B(_0331_),
    .C(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_1 _1256_ (.A(_0575_),
    .X(\clk8.next_count[19] ));
 sky130_fd_sc_hd__o21ai_1 _1257_ (.A1(net56),
    .A2(_0573_),
    .B1(_0531_),
    .Y(_0576_));
 sky130_fd_sc_hd__a21oi_1 _1258_ (.A1(net56),
    .A2(_0573_),
    .B1(_0576_),
    .Y(\clk8.next_count[20] ));
 sky130_fd_sc_hd__and2b_1 _1259_ (.A_N(\kp_encoder.last_sk ),
    .B(\kp_encoder.sync_out[14] ),
    .X(_0577_));
 sky130_fd_sc_hd__nand2_1 _1260_ (.A(\SS_FSM.sound[0] ),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__or2_1 _1261_ (.A(\SS_FSM.sound[0] ),
    .B(_0577_),
    .X(_0579_));
 sky130_fd_sc_hd__and2_1 _1262_ (.A(_0578_),
    .B(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_1 _1263_ (.A(_0580_),
    .X(\SS_FSM.next_sound[0] ));
 sky130_fd_sc_hd__a22o_1 _1264_ (.A1(_0274_),
    .A2(_0577_),
    .B1(_0578_),
    .B2(\SS_FSM.sound[1] ),
    .X(\SS_FSM.next_sound[1] ));
 sky130_fd_sc_hd__inv_2 _1265_ (.A(\mode_FSM.mode[1] ),
    .Y(_0581_));
 sky130_fd_sc_hd__and2_2 _1266_ (.A(_0581_),
    .B(\mode_FSM.mode[0] ),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _1267_ (.A(\seq_div.q_out[6] ),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__o21a_1 _1268_ (.A1(\mode_FSM.mode[1] ),
    .A2(\seq_div.q_out[6] ),
    .B1(\mode_FSM.mode[0] ),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_4 _1269_ (.A(\seq_div.q_out[7] ),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _1270_ (.A0(_0583_),
    .A1(_0584_),
    .S(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _1271_ (.A(\mode_FSM.mode[1] ),
    .B(\mode_FSM.mode[0] ),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_2 _1272_ (.A(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__o21ai_1 _1273_ (.A1(_0585_),
    .A2(\seq_div.q_out[5] ),
    .B1(_0582_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21o_1 _1274_ (.A1(_0585_),
    .A2(\seq_div.q_out[5] ),
    .B1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__o21ba_2 _1275_ (.A1(_0581_),
    .A2(_0585_),
    .B1_N(\mode_FSM.mode[0] ),
    .X(_0591_));
 sky130_fd_sc_hd__inv_2 _1276_ (.A(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__a2bb2o_1 _1277_ (.A1_N(\seq_div.q_out[6] ),
    .A2_N(_0588_),
    .B1(_0590_),
    .B2(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__or2_1 _1278_ (.A(_0585_),
    .B(\seq_div.q_out[4] ),
    .X(_0594_));
 sky130_fd_sc_hd__nand2_1 _1279_ (.A(_0585_),
    .B(\seq_div.q_out[4] ),
    .Y(_0595_));
 sky130_fd_sc_hd__a31o_1 _1280_ (.A1(_0582_),
    .A2(_0594_),
    .A3(_0595_),
    .B1(_0591_),
    .X(_0596_));
 sky130_fd_sc_hd__o21ai_1 _1281_ (.A1(\seq_div.q_out[5] ),
    .A2(_0588_),
    .B1(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__or2_1 _1282_ (.A(_0585_),
    .B(\seq_div.q_out[3] ),
    .X(_0598_));
 sky130_fd_sc_hd__nand2_1 _1283_ (.A(_0585_),
    .B(\seq_div.q_out[3] ),
    .Y(_0599_));
 sky130_fd_sc_hd__a31o_1 _1284_ (.A1(_0582_),
    .A2(_0598_),
    .A3(_0599_),
    .B1(_0591_),
    .X(_0600_));
 sky130_fd_sc_hd__o21ai_1 _1285_ (.A1(\seq_div.q_out[4] ),
    .A2(_0588_),
    .B1(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__or2_1 _1286_ (.A(_0585_),
    .B(\seq_div.q_out[2] ),
    .X(_0602_));
 sky130_fd_sc_hd__nand2_1 _1287_ (.A(_0585_),
    .B(\seq_div.q_out[2] ),
    .Y(_0603_));
 sky130_fd_sc_hd__a31o_1 _1288_ (.A1(_0582_),
    .A2(_0602_),
    .A3(_0603_),
    .B1(_0591_),
    .X(_0604_));
 sky130_fd_sc_hd__o21ai_1 _1289_ (.A1(\seq_div.q_out[3] ),
    .A2(_0588_),
    .B1(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__or2_1 _1290_ (.A(_0585_),
    .B(\seq_div.q_out[1] ),
    .X(_0606_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(_0585_),
    .B(\seq_div.q_out[1] ),
    .Y(_0607_));
 sky130_fd_sc_hd__a31o_1 _1292_ (.A1(_0582_),
    .A2(_0606_),
    .A3(_0607_),
    .B1(_0591_),
    .X(_0608_));
 sky130_fd_sc_hd__o21ai_1 _1293_ (.A1(\seq_div.q_out[2] ),
    .A2(_0588_),
    .B1(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_1 _1294_ (.A(\mode_FSM.mode[1] ),
    .B(\seq_div.q_out[0] ),
    .Y(_0610_));
 sky130_fd_sc_hd__or2_1 _1295_ (.A(_0585_),
    .B(\seq_div.q_out[0] ),
    .X(_0611_));
 sky130_fd_sc_hd__nand2_1 _1296_ (.A(_0585_),
    .B(\seq_div.q_out[0] ),
    .Y(_0612_));
 sky130_fd_sc_hd__a31o_1 _1297_ (.A1(_0582_),
    .A2(_0611_),
    .A3(_0612_),
    .B1(_0591_),
    .X(_0613_));
 sky130_fd_sc_hd__o21ai_1 _1298_ (.A1(\seq_div.q_out[1] ),
    .A2(_0588_),
    .B1(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__or4_1 _1299_ (.A(\pwm.count[0] ),
    .B(_0592_),
    .C(_0610_),
    .D(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__o31a_1 _1300_ (.A1(\pwm.count[0] ),
    .A2(_0592_),
    .A3(_0610_),
    .B1(_0614_),
    .X(_0616_));
 sky130_fd_sc_hd__a221o_1 _1301_ (.A1(\pwm.count[1] ),
    .A2(_0615_),
    .B1(_0609_),
    .B2(\pwm.count[2] ),
    .C1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__o221a_1 _1302_ (.A1(\pwm.count[2] ),
    .A2(_0609_),
    .B1(_0605_),
    .B2(\pwm.count[3] ),
    .C1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__a221o_1 _1303_ (.A1(\pwm.count[3] ),
    .A2(_0605_),
    .B1(_0601_),
    .B2(\pwm.count[4] ),
    .C1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__o221a_1 _1304_ (.A1(\pwm.count[4] ),
    .A2(_0601_),
    .B1(_0597_),
    .B2(\pwm.count[5] ),
    .C1(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__a221o_1 _1305_ (.A1(\pwm.count[5] ),
    .A2(_0597_),
    .B1(_0593_),
    .B2(\pwm.count[6] ),
    .C1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__o221a_1 _1306_ (.A1(\pwm.count[6] ),
    .A2(_0593_),
    .B1(_0586_),
    .B2(net67),
    .C1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__a211oi_1 _1307_ (.A1(net61),
    .A2(_0586_),
    .B1(_0622_),
    .C1(_0350_),
    .Y(\pwm.pwm ));
 sky130_fd_sc_hd__inv_2 _1308_ (.A(\seq_div.state[1] ),
    .Y(_0623_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(_0623_),
    .B(\seq_div.state[0] ),
    .X(_0624_));
 sky130_fd_sc_hd__clkbuf_4 _1310_ (.A(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__xnor2_1 _1311_ (.A(net86),
    .B(_0625_),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2_1 _1312_ (.A(_0623_),
    .B(\seq_div.state[0] ),
    .Y(_0626_));
 sky130_fd_sc_hd__and3_1 _1313_ (.A(\seq_div.count_div[0] ),
    .B(\seq_div.count_div[1] ),
    .C(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_8 _1314_ (.A(_0626_),
    .X(_0628_));
 sky130_fd_sc_hd__a21oi_1 _1315_ (.A1(\seq_div.count_div[0] ),
    .A2(_0628_),
    .B1(net84),
    .Y(_0629_));
 sky130_fd_sc_hd__nor2_1 _1316_ (.A(_0627_),
    .B(net85),
    .Y(_0001_));
 sky130_fd_sc_hd__xor2_1 _1317_ (.A(net57),
    .B(_0627_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1318_ (.A(_0623_),
    .B(\seq_div.state[0] ),
    .X(_0630_));
 sky130_fd_sc_hd__clkbuf_4 _1319_ (.A(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__buf_6 _1320_ (.A(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__nor2_1 _1321_ (.A(_0626_),
    .B(_0631_),
    .Y(_0633_));
 sky130_fd_sc_hd__clkbuf_8 _1322_ (.A(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__or2b_1 _1323_ (.A(\seq_div.R[18] ),
    .B_N(\seq_div.D[11] ),
    .X(_0635_));
 sky130_fd_sc_hd__or2b_1 _1324_ (.A(\seq_div.R[17] ),
    .B_N(\seq_div.D[10] ),
    .X(_0636_));
 sky130_fd_sc_hd__or2b_1 _1325_ (.A(\seq_div.R[15] ),
    .B_N(\seq_div.D[8] ),
    .X(_0637_));
 sky130_fd_sc_hd__or2b_1 _1326_ (.A(\seq_div.R[14] ),
    .B_N(\seq_div.D[7] ),
    .X(_0638_));
 sky130_fd_sc_hd__inv_2 _1327_ (.A(\seq_div.R[16] ),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _1328_ (.A(\seq_div.D[9] ),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__and3_1 _1329_ (.A(_0637_),
    .B(_0638_),
    .C(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__and2b_1 _1330_ (.A_N(\seq_div.D[1] ),
    .B(\seq_div.R[8] ),
    .X(_0642_));
 sky130_fd_sc_hd__or2b_1 _1331_ (.A(\seq_div.R[9] ),
    .B_N(\seq_div.D[2] ),
    .X(_0643_));
 sky130_fd_sc_hd__and2b_1 _1332_ (.A_N(\seq_div.D[3] ),
    .B(\seq_div.R[10] ),
    .X(_0644_));
 sky130_fd_sc_hd__and2b_1 _1333_ (.A_N(\seq_div.D[2] ),
    .B(\seq_div.R[9] ),
    .X(_0645_));
 sky130_fd_sc_hd__a211o_1 _1334_ (.A1(_0642_),
    .A2(_0643_),
    .B1(_0644_),
    .C1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__or2b_1 _1335_ (.A(\seq_div.R[11] ),
    .B_N(\seq_div.D[4] ),
    .X(_0647_));
 sky130_fd_sc_hd__or2b_1 _1336_ (.A(\seq_div.R[10] ),
    .B_N(\seq_div.D[3] ),
    .X(_0648_));
 sky130_fd_sc_hd__and3_1 _1337_ (.A(_0646_),
    .B(_0647_),
    .C(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__and2b_1 _1338_ (.A_N(\seq_div.D[5] ),
    .B(\seq_div.R[12] ),
    .X(_0650_));
 sky130_fd_sc_hd__or2b_1 _1339_ (.A(\seq_div.D[4] ),
    .B_N(\seq_div.R[11] ),
    .X(_0651_));
 sky130_fd_sc_hd__or3b_1 _1340_ (.A(_0649_),
    .B(_0650_),
    .C_N(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or2b_1 _1341_ (.A(\seq_div.R[13] ),
    .B_N(\seq_div.D[6] ),
    .X(_0653_));
 sky130_fd_sc_hd__or2b_1 _1342_ (.A(\seq_div.R[12] ),
    .B_N(\seq_div.D[5] ),
    .X(_0654_));
 sky130_fd_sc_hd__and2b_1 _1343_ (.A_N(\seq_div.D[7] ),
    .B(\seq_div.R[14] ),
    .X(_0655_));
 sky130_fd_sc_hd__and2b_1 _1344_ (.A_N(\seq_div.D[6] ),
    .B(\seq_div.R[13] ),
    .X(_0656_));
 sky130_fd_sc_hd__a311o_1 _1345_ (.A1(_0652_),
    .A2(_0653_),
    .A3(_0654_),
    .B1(_0655_),
    .C1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__and2b_1 _1346_ (.A_N(\seq_div.D[10] ),
    .B(\seq_div.R[17] ),
    .X(_0658_));
 sky130_fd_sc_hd__or2_1 _1347_ (.A(\seq_div.D[9] ),
    .B(_0639_),
    .X(_0659_));
 sky130_fd_sc_hd__or2b_1 _1348_ (.A(\seq_div.D[8] ),
    .B_N(\seq_div.R[15] ),
    .X(_0660_));
 sky130_fd_sc_hd__a21boi_1 _1349_ (.A1(_0659_),
    .A2(_0660_),
    .B1_N(_0640_),
    .Y(_0661_));
 sky130_fd_sc_hd__a211o_1 _1350_ (.A1(_0641_),
    .A2(_0657_),
    .B1(_0658_),
    .C1(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__or2b_1 _1351_ (.A(\seq_div.D[11] ),
    .B_N(\seq_div.R[18] ),
    .X(_0663_));
 sky130_fd_sc_hd__nand2_1 _1352_ (.A(_0635_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__a21o_1 _1353_ (.A1(_0636_),
    .A2(_0662_),
    .B1(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__or2b_1 _1354_ (.A(\seq_div.R[19] ),
    .B_N(\seq_div.D[12] ),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _1355_ (.A(_0635_),
    .B(_0665_),
    .C(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__or2b_1 _1356_ (.A(\seq_div.R[20] ),
    .B_N(\seq_div.D[13] ),
    .X(_0668_));
 sky130_fd_sc_hd__and2b_1 _1357_ (.A_N(\seq_div.D[13] ),
    .B(\seq_div.R[20] ),
    .X(_0669_));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _1359_ (.A(_0668_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__or2b_1 _1360_ (.A(\seq_div.R[21] ),
    .B_N(\seq_div.D[14] ),
    .X(_0672_));
 sky130_fd_sc_hd__or2b_1 _1361_ (.A(\seq_div.D[14] ),
    .B_N(\seq_div.R[21] ),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_1 _1362_ (.A(_0672_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__or2_1 _1363_ (.A(_0671_),
    .B(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__or2b_1 _1364_ (.A(\seq_div.D[12] ),
    .B_N(\seq_div.R[19] ),
    .X(_0676_));
 sky130_fd_sc_hd__or3b_1 _1365_ (.A(_0667_),
    .B(_0675_),
    .C_N(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__inv_2 _1366_ (.A(\seq_div.D[15] ),
    .Y(_0678_));
 sky130_fd_sc_hd__and2b_1 _1367_ (.A_N(\seq_div.D[14] ),
    .B(\seq_div.R[21] ),
    .X(_0679_));
 sky130_fd_sc_hd__o221a_1 _1368_ (.A1(_0678_),
    .A2(\seq_div.R[22] ),
    .B1(_0668_),
    .B2(_0679_),
    .C1(_0672_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(_0677_),
    .B(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _1370_ (.A(_0678_),
    .B(\seq_div.R[22] ),
    .Y(_0682_));
 sky130_fd_sc_hd__or2b_1 _1371_ (.A(_0650_),
    .B_N(_0654_),
    .X(_0683_));
 sky130_fd_sc_hd__or2b_1 _1372_ (.A(_0644_),
    .B_N(_0648_),
    .X(_0684_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(_0645_),
    .Y(_0685_));
 sky130_fd_sc_hd__nand2_1 _1374_ (.A(_0643_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _1375_ (.A(_0647_),
    .B(_0651_),
    .Y(_0687_));
 sky130_fd_sc_hd__or3_1 _1376_ (.A(_0684_),
    .B(_0686_),
    .C(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__inv_2 _1377_ (.A(_0636_),
    .Y(_0689_));
 sky130_fd_sc_hd__or3_1 _1378_ (.A(_0664_),
    .B(_0689_),
    .C(_0658_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(_0640_),
    .B(_0659_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand2_1 _1380_ (.A(_0637_),
    .B(_0660_),
    .Y(_0692_));
 sky130_fd_sc_hd__or3_1 _1381_ (.A(_0690_),
    .B(_0691_),
    .C(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__or2b_1 _1382_ (.A(\seq_div.R[8] ),
    .B_N(\seq_div.D[1] ),
    .X(_0694_));
 sky130_fd_sc_hd__and2b_1 _1383_ (.A_N(_0642_),
    .B(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__or3b_1 _1384_ (.A(\seq_div.D[0] ),
    .B(_0675_),
    .C_N(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__and2b_1 _1385_ (.A_N(\seq_div.R[14] ),
    .B(\seq_div.D[7] ),
    .X(_0697_));
 sky130_fd_sc_hd__or2b_1 _1386_ (.A(\seq_div.D[6] ),
    .B_N(\seq_div.R[13] ),
    .X(_0698_));
 sky130_fd_sc_hd__nand2_1 _1387_ (.A(_0653_),
    .B(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__or3_1 _1388_ (.A(_0697_),
    .B(_0655_),
    .C(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nand2_1 _1389_ (.A(_0666_),
    .B(_0676_),
    .Y(_0701_));
 sky130_fd_sc_hd__xnor2_1 _1390_ (.A(\seq_div.D[15] ),
    .B(\seq_div.R[22] ),
    .Y(_0702_));
 sky130_fd_sc_hd__or4b_1 _1391_ (.A(_0696_),
    .B(_0700_),
    .C(_0701_),
    .D_N(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__or4_1 _1392_ (.A(_0683_),
    .B(_0688_),
    .C(_0693_),
    .D(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__and4b_1 _1393_ (.A_N(\seq_div.R[23] ),
    .B(_0681_),
    .C(_0682_),
    .D(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__clkbuf_2 _1394_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_6 _1395_ (.A(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__and3b_1 _1396_ (.A_N(_0707_),
    .B(_0628_),
    .C(\seq_div.D[0] ),
    .X(_0708_));
 sky130_fd_sc_hd__a221o_1 _1397_ (.A1(net68),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[8] ),
    .C1(_0708_),
    .X(_0003_));
 sky130_fd_sc_hd__xnor2_1 _1398_ (.A(\seq_div.D[0] ),
    .B(_0695_),
    .Y(_0709_));
 sky130_fd_sc_hd__mux2_1 _1399_ (.A0(_0709_),
    .A1(\seq_div.R[8] ),
    .S(_0707_),
    .X(_0710_));
 sky130_fd_sc_hd__a22o_1 _1400_ (.A1(net113),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[9] ),
    .X(_0711_));
 sky130_fd_sc_hd__a21o_1 _1401_ (.A1(_0628_),
    .A2(_0710_),
    .B1(_0711_),
    .X(_0004_));
 sky130_fd_sc_hd__nand2_4 _1402_ (.A(_0623_),
    .B(\seq_div.state[0] ),
    .Y(_0712_));
 sky130_fd_sc_hd__inv_2 _1403_ (.A(\seq_div.D[0] ),
    .Y(_0713_));
 sky130_fd_sc_hd__a21o_1 _1404_ (.A1(_0713_),
    .A2(_0694_),
    .B1(_0642_),
    .X(_0714_));
 sky130_fd_sc_hd__xnor2_1 _1405_ (.A(_0686_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__mux2_1 _1406_ (.A0(_0715_),
    .A1(\seq_div.R[9] ),
    .S(_0707_),
    .X(_0716_));
 sky130_fd_sc_hd__nand2_2 _1407_ (.A(_0625_),
    .B(_0712_),
    .Y(_0717_));
 sky130_fd_sc_hd__or2_1 _1408_ (.A(\seq_div.R[10] ),
    .B(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__o221a_1 _1409_ (.A1(net96),
    .A2(_0712_),
    .B1(_0716_),
    .B2(_0625_),
    .C1(_0718_),
    .X(_0005_));
 sky130_fd_sc_hd__a21o_1 _1410_ (.A1(_0643_),
    .A2(_0714_),
    .B1(_0645_),
    .X(_0719_));
 sky130_fd_sc_hd__xnor2_1 _1411_ (.A(_0684_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__mux2_1 _1412_ (.A0(_0720_),
    .A1(\seq_div.R[10] ),
    .S(_0707_),
    .X(_0721_));
 sky130_fd_sc_hd__a22o_1 _1413_ (.A1(\seq_div.dividend[3] ),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[11] ),
    .X(_0722_));
 sky130_fd_sc_hd__a21o_1 _1414_ (.A1(_0628_),
    .A2(_0721_),
    .B1(_0722_),
    .X(_0006_));
 sky130_fd_sc_hd__a21oi_1 _1415_ (.A1(_0648_),
    .A2(_0719_),
    .B1(_0644_),
    .Y(_0723_));
 sky130_fd_sc_hd__xor2_1 _1416_ (.A(_0687_),
    .B(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _1417_ (.A0(_0724_),
    .A1(\seq_div.R[11] ),
    .S(_0707_),
    .X(_0725_));
 sky130_fd_sc_hd__or2_1 _1418_ (.A(\seq_div.R[12] ),
    .B(_0717_),
    .X(_0726_));
 sky130_fd_sc_hd__o221a_1 _1419_ (.A1(net83),
    .A2(_0712_),
    .B1(_0725_),
    .B2(_0625_),
    .C1(_0726_),
    .X(_0007_));
 sky130_fd_sc_hd__o21ai_1 _1420_ (.A1(_0687_),
    .A2(_0723_),
    .B1(_0651_),
    .Y(_0727_));
 sky130_fd_sc_hd__xnor2_1 _1421_ (.A(_0683_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__mux2_1 _1422_ (.A0(_0728_),
    .A1(\seq_div.R[12] ),
    .S(_0707_),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _1423_ (.A1(net107),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[13] ),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_1 _1424_ (.A1(_0628_),
    .A2(_0729_),
    .B1(_0730_),
    .X(_0008_));
 sky130_fd_sc_hd__a21o_1 _1425_ (.A1(_0654_),
    .A2(_0727_),
    .B1(_0650_),
    .X(_0731_));
 sky130_fd_sc_hd__xnor2_1 _1426_ (.A(_0699_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__mux2_1 _1427_ (.A0(_0732_),
    .A1(\seq_div.R[13] ),
    .S(_0707_),
    .X(_0733_));
 sky130_fd_sc_hd__a22o_1 _1428_ (.A1(net78),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[14] ),
    .X(_0734_));
 sky130_fd_sc_hd__a21o_1 _1429_ (.A1(_0628_),
    .A2(_0733_),
    .B1(_0734_),
    .X(_0009_));
 sky130_fd_sc_hd__nor2_1 _1430_ (.A(_0697_),
    .B(_0655_),
    .Y(_0735_));
 sky130_fd_sc_hd__a21o_1 _1431_ (.A1(_0653_),
    .A2(_0731_),
    .B1(_0656_),
    .X(_0736_));
 sky130_fd_sc_hd__or2_1 _1432_ (.A(_0735_),
    .B(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__a21oi_1 _1433_ (.A1(_0735_),
    .A2(_0736_),
    .B1(_0706_),
    .Y(_0738_));
 sky130_fd_sc_hd__a22o_1 _1434_ (.A1(\seq_div.R[14] ),
    .A2(_0707_),
    .B1(_0737_),
    .B2(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__or2_1 _1435_ (.A(\seq_div.R[15] ),
    .B(_0717_),
    .X(_0740_));
 sky130_fd_sc_hd__o221a_1 _1436_ (.A1(net98),
    .A2(_0712_),
    .B1(_0739_),
    .B2(_0625_),
    .C1(_0740_),
    .X(_0010_));
 sky130_fd_sc_hd__a21oi_1 _1437_ (.A1(_0638_),
    .A2(_0736_),
    .B1(_0655_),
    .Y(_0741_));
 sky130_fd_sc_hd__or2_1 _1438_ (.A(_0692_),
    .B(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__a21oi_1 _1439_ (.A1(_0692_),
    .A2(_0741_),
    .B1(_0706_),
    .Y(_0743_));
 sky130_fd_sc_hd__a221o_1 _1440_ (.A1(\seq_div.R[15] ),
    .A2(_0707_),
    .B1(_0742_),
    .B2(_0743_),
    .C1(_0625_),
    .X(_0744_));
 sky130_fd_sc_hd__o221a_1 _1441_ (.A1(net99),
    .A2(_0712_),
    .B1(_0717_),
    .B2(\seq_div.R[16] ),
    .C1(_0744_),
    .X(_0011_));
 sky130_fd_sc_hd__nand2_1 _1442_ (.A(_0660_),
    .B(_0742_),
    .Y(_0745_));
 sky130_fd_sc_hd__xor2_1 _1443_ (.A(_0691_),
    .B(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__nor2_1 _1444_ (.A(_0707_),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__a211o_1 _1445_ (.A1(\seq_div.R[16] ),
    .A2(_0707_),
    .B1(_0747_),
    .C1(_0625_),
    .X(_0748_));
 sky130_fd_sc_hd__o221a_1 _1446_ (.A1(net88),
    .A2(_0712_),
    .B1(_0717_),
    .B2(\seq_div.R[17] ),
    .C1(_0748_),
    .X(_0012_));
 sky130_fd_sc_hd__nor2_1 _1447_ (.A(_0689_),
    .B(_0658_),
    .Y(_0749_));
 sky130_fd_sc_hd__o21bai_1 _1448_ (.A1(_0691_),
    .A2(_0742_),
    .B1_N(_0661_),
    .Y(_0750_));
 sky130_fd_sc_hd__or2_1 _1449_ (.A(_0749_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__a21oi_1 _1450_ (.A1(_0749_),
    .A2(_0750_),
    .B1(_0706_),
    .Y(_0752_));
 sky130_fd_sc_hd__a221o_1 _1451_ (.A1(\seq_div.R[17] ),
    .A2(_0707_),
    .B1(_0751_),
    .B2(_0752_),
    .C1(_0625_),
    .X(_0753_));
 sky130_fd_sc_hd__o221a_1 _1452_ (.A1(net91),
    .A2(_0712_),
    .B1(_0717_),
    .B2(\seq_div.R[18] ),
    .C1(_0753_),
    .X(_0013_));
 sky130_fd_sc_hd__a21o_1 _1453_ (.A1(_0749_),
    .A2(_0750_),
    .B1(_0658_),
    .X(_0754_));
 sky130_fd_sc_hd__xnor2_1 _1454_ (.A(_0664_),
    .B(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(_0755_),
    .A1(\seq_div.R[18] ),
    .S(_0707_),
    .X(_0756_));
 sky130_fd_sc_hd__a22o_1 _1456_ (.A1(net117),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[19] ),
    .X(_0757_));
 sky130_fd_sc_hd__a21o_1 _1457_ (.A1(_0628_),
    .A2(_0756_),
    .B1(_0757_),
    .X(_0014_));
 sky130_fd_sc_hd__a21boi_1 _1458_ (.A1(_0635_),
    .A2(_0658_),
    .B1_N(_0663_),
    .Y(_0758_));
 sky130_fd_sc_hd__or4b_1 _1459_ (.A(_0664_),
    .B(_0689_),
    .C(_0658_),
    .D_N(_0661_),
    .X(_0759_));
 sky130_fd_sc_hd__o211a_1 _1460_ (.A1(_0693_),
    .A2(_0741_),
    .B1(_0758_),
    .C1(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__xor2_1 _1461_ (.A(_0701_),
    .B(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _1462_ (.A0(_0761_),
    .A1(\seq_div.R[19] ),
    .S(_0707_),
    .X(_0762_));
 sky130_fd_sc_hd__a22o_1 _1463_ (.A1(\seq_div.dividend[12] ),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[20] ),
    .X(_0763_));
 sky130_fd_sc_hd__a21o_1 _1464_ (.A1(_0628_),
    .A2(_0762_),
    .B1(_0763_),
    .X(_0015_));
 sky130_fd_sc_hd__o21ai_2 _1465_ (.A1(_0701_),
    .A2(_0760_),
    .B1(_0676_),
    .Y(_0764_));
 sky130_fd_sc_hd__xnor2_1 _1466_ (.A(_0671_),
    .B(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(_0765_),
    .A1(\seq_div.R[20] ),
    .S(_0707_),
    .X(_0766_));
 sky130_fd_sc_hd__a22o_1 _1468_ (.A1(net114),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[21] ),
    .X(_0767_));
 sky130_fd_sc_hd__a21o_1 _1469_ (.A1(_0628_),
    .A2(_0766_),
    .B1(_0767_),
    .X(_0016_));
 sky130_fd_sc_hd__a21o_1 _1470_ (.A1(_0668_),
    .A2(_0764_),
    .B1(_0669_),
    .X(_0768_));
 sky130_fd_sc_hd__xnor2_1 _1471_ (.A(_0674_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(_0769_),
    .A1(\seq_div.R[21] ),
    .S(_0707_),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _1473_ (.A1(net111),
    .A2(_0632_),
    .B1(_0634_),
    .B2(\seq_div.R[22] ),
    .X(_0771_));
 sky130_fd_sc_hd__a21o_1 _1474_ (.A1(_0628_),
    .A2(_0770_),
    .B1(_0771_),
    .X(_0017_));
 sky130_fd_sc_hd__a21oi_1 _1475_ (.A1(_0672_),
    .A2(_0768_),
    .B1(_0679_),
    .Y(_0772_));
 sky130_fd_sc_hd__xnor2_1 _1476_ (.A(_0702_),
    .B(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(_0773_),
    .A1(\seq_div.R[22] ),
    .S(_0707_),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _1478_ (.A1(\seq_div.dividend[15] ),
    .A2(_0632_),
    .B1(_0633_),
    .B2(net108),
    .X(_0775_));
 sky130_fd_sc_hd__a21o_1 _1479_ (.A1(_0628_),
    .A2(_0774_),
    .B1(net109),
    .X(_0018_));
 sky130_fd_sc_hd__nand2_4 _1480_ (.A(\seq_div.state[1] ),
    .B(\seq_div.state[0] ),
    .Y(_0776_));
 sky130_fd_sc_hd__mux2_1 _1481_ (.A0(net120),
    .A1(\seq_div.q_out[0] ),
    .S(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__clkbuf_1 _1482_ (.A(_0777_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(\seq_div.Q[1] ),
    .A1(\seq_div.q_out[1] ),
    .S(_0776_),
    .X(_0778_));
 sky130_fd_sc_hd__clkbuf_1 _1484_ (.A(_0778_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(\seq_div.Q[2] ),
    .A1(\seq_div.q_out[2] ),
    .S(_0776_),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _1486_ (.A(_0080_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(net122),
    .A1(\seq_div.q_out[3] ),
    .S(_0776_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _1488_ (.A(_0081_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(net121),
    .A1(\seq_div.q_out[4] ),
    .S(_0776_),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_1 _1490_ (.A(_0082_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1491_ (.A0(net62),
    .A1(\seq_div.q_out[5] ),
    .S(_0776_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_1 _1492_ (.A(_0083_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(\seq_div.Q[6] ),
    .A1(\seq_div.q_out[6] ),
    .S(_0776_),
    .X(_0084_));
 sky130_fd_sc_hd__clkbuf_1 _1494_ (.A(_0084_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(net59),
    .A1(_0585_),
    .S(_0776_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_0085_),
    .X(_0026_));
 sky130_fd_sc_hd__a2bb2o_1 _1497_ (.A1_N(_0625_),
    .A2_N(_0707_),
    .B1(_0634_),
    .B2(net81),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_1 _1498_ (.A1(net81),
    .A2(_0628_),
    .B1(_0634_),
    .B2(\seq_div.Q[1] ),
    .X(_0028_));
 sky130_fd_sc_hd__a22o_1 _1499_ (.A1(\seq_div.Q[1] ),
    .A2(_0628_),
    .B1(_0634_),
    .B2(net79),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _1500_ (.A1(\seq_div.Q[2] ),
    .A2(_0628_),
    .B1(_0634_),
    .B2(net75),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _1501_ (.A1(net75),
    .A2(_0628_),
    .B1(_0634_),
    .B2(net77),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _1502_ (.A1(net77),
    .A2(_0628_),
    .B1(_0634_),
    .B2(net62),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _1503_ (.A1(net62),
    .A2(_0628_),
    .B1(_0634_),
    .B2(\seq_div.Q[6] ),
    .X(_0033_));
 sky130_fd_sc_hd__a22o_1 _1504_ (.A1(\seq_div.Q[6] ),
    .A2(_0628_),
    .B1(_0634_),
    .B2(net59),
    .X(_0034_));
 sky130_fd_sc_hd__nand2_1 _1505_ (.A(net104),
    .B(_0712_),
    .Y(_0086_));
 sky130_fd_sc_hd__o21ai_1 _1506_ (.A1(_0430_),
    .A2(_0712_),
    .B1(_0086_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1507_ (.A(_0427_),
    .Y(_0087_));
 sky130_fd_sc_hd__mux2_1 _1508_ (.A0(\seq_div.D[1] ),
    .A1(_0087_),
    .S(_0632_),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _1509_ (.A(_0088_),
    .X(_0036_));
 sky130_fd_sc_hd__inv_2 _1510_ (.A(_0422_),
    .Y(_0089_));
 sky130_fd_sc_hd__mux2_1 _1511_ (.A0(\seq_div.D[2] ),
    .A1(_0089_),
    .S(_0632_),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _1512_ (.A(_0090_),
    .X(_0037_));
 sky130_fd_sc_hd__inv_2 _1513_ (.A(_0420_),
    .Y(_0091_));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(\seq_div.D[3] ),
    .A1(_0091_),
    .S(_0632_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _1515_ (.A(_0092_),
    .X(_0038_));
 sky130_fd_sc_hd__nand2_1 _1516_ (.A(_0381_),
    .B(_0392_),
    .Y(_0093_));
 sky130_fd_sc_hd__mux2_1 _1517_ (.A0(\seq_div.D[4] ),
    .A1(_0093_),
    .S(_0632_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _1518_ (.A(_0094_),
    .X(_0039_));
 sky130_fd_sc_hd__inv_2 _1519_ (.A(_0435_),
    .Y(_0095_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(net118),
    .A1(_0095_),
    .S(_0632_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_1 _1521_ (.A(_0096_),
    .X(_0040_));
 sky130_fd_sc_hd__a31o_1 _1522_ (.A1(_0382_),
    .A2(_0375_),
    .A3(_0391_),
    .B1(_0712_),
    .X(_0097_));
 sky130_fd_sc_hd__o21a_1 _1523_ (.A1(net87),
    .A2(_0632_),
    .B1(_0097_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(\seq_div.D[7] ),
    .A1(_0419_),
    .S(_0632_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _1525_ (.A(_0098_),
    .X(_0042_));
 sky130_fd_sc_hd__nand2_1 _1526_ (.A(_0393_),
    .B(_0407_),
    .Y(_0099_));
 sky130_fd_sc_hd__mux2_1 _1527_ (.A0(\seq_div.D[8] ),
    .A1(_0099_),
    .S(_0632_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _1528_ (.A(_0100_),
    .X(_0043_));
 sky130_fd_sc_hd__inv_2 _1529_ (.A(_0408_),
    .Y(_0101_));
 sky130_fd_sc_hd__mux2_1 _1530_ (.A0(\seq_div.D[9] ),
    .A1(_0101_),
    .S(_0631_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _1531_ (.A(_0102_),
    .X(_0044_));
 sky130_fd_sc_hd__inv_2 _1532_ (.A(_0411_),
    .Y(_0103_));
 sky130_fd_sc_hd__mux2_1 _1533_ (.A0(net119),
    .A1(_0103_),
    .S(_0631_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _1534_ (.A(_0104_),
    .X(_0045_));
 sky130_fd_sc_hd__inv_2 _1535_ (.A(_0395_),
    .Y(_0105_));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(\seq_div.D[11] ),
    .A1(_0105_),
    .S(_0631_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _1537_ (.A(_0106_),
    .X(_0046_));
 sky130_fd_sc_hd__inv_2 _1538_ (.A(_0385_),
    .Y(_0107_));
 sky130_fd_sc_hd__mux2_1 _1539_ (.A0(net115),
    .A1(_0107_),
    .S(_0631_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _1540_ (.A(_0108_),
    .X(_0047_));
 sky130_fd_sc_hd__inv_2 _1541_ (.A(_0387_),
    .Y(_0109_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(\seq_div.D[13] ),
    .A1(_0109_),
    .S(_0631_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _1543_ (.A(_0110_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(\seq_div.D[14] ),
    .A1(_0402_),
    .S(_0631_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _1545_ (.A(_0111_),
    .X(_0049_));
 sky130_fd_sc_hd__nor2_1 _1546_ (.A(_0382_),
    .B(_0397_),
    .Y(_0112_));
 sky130_fd_sc_hd__mux2_1 _1547_ (.A0(\seq_div.D[15] ),
    .A1(_0112_),
    .S(_0631_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _1548_ (.A(_0113_),
    .X(_0050_));
 sky130_fd_sc_hd__nor2_1 _1549_ (.A(_0350_),
    .B(_0529_),
    .Y(_0114_));
 sky130_fd_sc_hd__nor2_1 _1550_ (.A(_0240_),
    .B(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__or3_1 _1551_ (.A(_0196_),
    .B(_0193_),
    .C(_0222_),
    .X(_0116_));
 sky130_fd_sc_hd__a41o_1 _1552_ (.A1(_0172_),
    .A2(_0173_),
    .A3(_0269_),
    .A4(_0116_),
    .B1(_0236_),
    .X(_0117_));
 sky130_fd_sc_hd__nand2_1 _1553_ (.A(_0179_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__and2_1 _1554_ (.A(\SS_FSM.sound[0] ),
    .B(_0114_),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _1555_ (.A1(_0179_),
    .A2(_0115_),
    .B1(_0118_),
    .B2(_0119_),
    .X(_0051_));
 sky130_fd_sc_hd__a32o_1 _1556_ (.A1(_0182_),
    .A2(_0117_),
    .A3(_0119_),
    .B1(_0115_),
    .B2(_0155_),
    .X(_0052_));
 sky130_fd_sc_hd__o41ai_1 _1557_ (.A1(\SS_FSM.sound[1] ),
    .A2(_0180_),
    .A3(_0181_),
    .A4(_0269_),
    .B1(\SS_FSM.sound[0] ),
    .Y(_0120_));
 sky130_fd_sc_hd__or3b_1 _1558_ (.A(_0219_),
    .B(net23),
    .C_N(_0117_),
    .X(_0121_));
 sky130_fd_sc_hd__or2_1 _1559_ (.A(_0240_),
    .B(_0114_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_2 _1560_ (.A(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1561_ (.A0(\SS_FSM.count[2] ),
    .A1(_0121_),
    .S(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _1562_ (.A(_0124_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _1563_ (.A(_0165_),
    .B(_0117_),
    .Y(_0125_));
 sky130_fd_sc_hd__a22o_1 _1564_ (.A1(\SS_FSM.count[3] ),
    .A2(_0115_),
    .B1(_0119_),
    .B2(_0125_),
    .X(_0054_));
 sky130_fd_sc_hd__nor2_1 _1565_ (.A(_0237_),
    .B(_0167_),
    .Y(_0126_));
 sky130_fd_sc_hd__a21o_1 _1566_ (.A1(_0174_),
    .A2(_0299_),
    .B1(_0115_),
    .X(_0127_));
 sky130_fd_sc_hd__o22a_1 _1567_ (.A1(\SS_FSM.count[4] ),
    .A2(_0123_),
    .B1(_0126_),
    .B2(_0127_),
    .X(_0055_));
 sky130_fd_sc_hd__nor2_1 _1568_ (.A(_0237_),
    .B(_0159_),
    .Y(_0128_));
 sky130_fd_sc_hd__o22a_1 _1569_ (.A1(\SS_FSM.count[5] ),
    .A2(_0123_),
    .B1(_0127_),
    .B2(_0128_),
    .X(_0056_));
 sky130_fd_sc_hd__nor2_1 _1570_ (.A(_0237_),
    .B(_0214_),
    .Y(_0129_));
 sky130_fd_sc_hd__o22a_1 _1571_ (.A1(\SS_FSM.count[6] ),
    .A2(_0123_),
    .B1(_0127_),
    .B2(_0129_),
    .X(_0057_));
 sky130_fd_sc_hd__nor2_1 _1572_ (.A(_0237_),
    .B(_0217_),
    .Y(_0130_));
 sky130_fd_sc_hd__o22a_1 _1573_ (.A1(net112),
    .A2(_0123_),
    .B1(_0127_),
    .B2(_0130_),
    .X(_0058_));
 sky130_fd_sc_hd__a211o_1 _1574_ (.A1(_0236_),
    .A2(_0175_),
    .B1(_0120_),
    .C1(_0127_),
    .X(_0131_));
 sky130_fd_sc_hd__o21a_1 _1575_ (.A1(net116),
    .A2(_0123_),
    .B1(_0131_),
    .X(_0059_));
 sky130_fd_sc_hd__nor2_8 _1576_ (.A(_0350_),
    .B(_0507_),
    .Y(_0132_));
 sky130_fd_sc_hd__mux2_1 _1577_ (.A0(net123),
    .A1(\osc.count[0] ),
    .S(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _1578_ (.A(_0133_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(net126),
    .A1(\osc.count[1] ),
    .S(_0132_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _1580_ (.A(_0134_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(net128),
    .A1(\osc.count[2] ),
    .S(_0132_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _1582_ (.A(_0135_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(\seq_div.dividend[3] ),
    .A1(\osc.count[3] ),
    .S(_0132_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _1584_ (.A(_0136_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1585_ (.A0(net124),
    .A1(\osc.count[4] ),
    .S(_0132_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _1586_ (.A(_0137_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1587_ (.A0(net127),
    .A1(\osc.count[5] ),
    .S(_0132_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _1588_ (.A(_0138_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1589_ (.A0(net78),
    .A1(\osc.count[6] ),
    .S(_0132_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _1590_ (.A(_0139_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1591_ (.A0(net98),
    .A1(\osc.count[7] ),
    .S(_0132_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _1592_ (.A(_0140_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1593_ (.A0(net99),
    .A1(\osc.count[8] ),
    .S(_0132_),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _1594_ (.A(_0141_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(net88),
    .A1(\osc.count[9] ),
    .S(_0132_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _1596_ (.A(_0142_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1597_ (.A0(net91),
    .A1(\osc.count[10] ),
    .S(_0132_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _1598_ (.A(_0143_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1599_ (.A0(net125),
    .A1(\osc.count[11] ),
    .S(_0132_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _1600_ (.A(_0144_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1601_ (.A0(\seq_div.dividend[12] ),
    .A1(\osc.count[12] ),
    .S(_0132_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _1602_ (.A(_0145_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1603_ (.A0(net129),
    .A1(\osc.count[13] ),
    .S(_0132_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _1604_ (.A(_0146_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1605_ (.A0(net130),
    .A1(\osc.count[14] ),
    .S(_0132_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _1606_ (.A(_0147_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(\seq_div.dividend[15] ),
    .A1(\osc.count[15] ),
    .S(_0132_),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _1608_ (.A(_0148_),
    .X(_0075_));
 sky130_fd_sc_hd__and2b_1 _1609_ (.A_N(\seq_div.state[0] ),
    .B(_0132_),
    .X(_0149_));
 sky130_fd_sc_hd__a31o_1 _1610_ (.A1(\seq_div.count_div[0] ),
    .A2(\seq_div.count_div[1] ),
    .A3(net57),
    .B1(_0625_),
    .X(_0150_));
 sky130_fd_sc_hd__o21a_1 _1611_ (.A1(net73),
    .A2(_0149_),
    .B1(_0150_),
    .X(_0076_));
 sky130_fd_sc_hd__o21ai_1 _1612_ (.A1(_0623_),
    .A2(_0132_),
    .B1(_0634_),
    .Y(_0077_));
 sky130_fd_sc_hd__and2b_1 _1613_ (.A_N(\kp_encoder.last_mk ),
    .B(\kp_encoder.sync_out[13] ),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(\mode_FSM.mode[1] ),
    .A1(\mode_FSM.mode[0] ),
    .S(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _1615_ (.A(_0152_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(\mode_FSM.mode[0] ),
    .A1(_0581_),
    .S(_0151_),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _1617_ (.A(_0153_),
    .X(_0079_));
 sky130_fd_sc_hd__dfrtp_1 _1618_ (.CLK(clknet_4_15_0_clk),
    .D(_0000_),
    .RESET_B(net37),
    .Q(\seq_div.count_div[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1619_ (.CLK(clknet_4_15_0_clk),
    .D(_0001_),
    .RESET_B(net37),
    .Q(\seq_div.count_div[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1620_ (.CLK(clknet_4_13_0_clk),
    .D(_0002_),
    .RESET_B(net37),
    .Q(\seq_div.count_div[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1621_ (.CLK(clknet_4_3_0_clk),
    .D(\SS_FSM.next_sound[0] ),
    .RESET_B(net30),
    .Q(\SS_FSM.sound[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1622_ (.CLK(clknet_4_3_0_clk),
    .D(\SS_FSM.next_sound[1] ),
    .RESET_B(net30),
    .Q(\SS_FSM.sound[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1623_ (.CLK(clknet_4_8_0_clk),
    .D(net69),
    .RESET_B(net34),
    .Q(\seq_div.R[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1624_ (.CLK(clknet_4_10_0_clk),
    .D(_0004_),
    .RESET_B(net34),
    .Q(\seq_div.R[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1625_ (.CLK(clknet_4_10_0_clk),
    .D(_0005_),
    .RESET_B(net34),
    .Q(\seq_div.R[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1626_ (.CLK(clknet_4_10_0_clk),
    .D(_0006_),
    .RESET_B(net34),
    .Q(\seq_div.R[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1627_ (.CLK(clknet_4_10_0_clk),
    .D(_0007_),
    .RESET_B(net34),
    .Q(\seq_div.R[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1628_ (.CLK(clknet_4_10_0_clk),
    .D(_0008_),
    .RESET_B(net34),
    .Q(\seq_div.R[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1629_ (.CLK(clknet_4_10_0_clk),
    .D(_0009_),
    .RESET_B(net34),
    .Q(\seq_div.R[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1630_ (.CLK(clknet_4_11_0_clk),
    .D(_0010_),
    .RESET_B(net34),
    .Q(\seq_div.R[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1631_ (.CLK(clknet_4_11_0_clk),
    .D(net100),
    .RESET_B(net34),
    .Q(\seq_div.R[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1632_ (.CLK(clknet_4_14_0_clk),
    .D(net89),
    .RESET_B(net34),
    .Q(\seq_div.R[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1633_ (.CLK(clknet_4_14_0_clk),
    .D(net92),
    .RESET_B(net37),
    .Q(\seq_div.R[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1634_ (.CLK(clknet_4_14_0_clk),
    .D(_0014_),
    .RESET_B(net37),
    .Q(\seq_div.R[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1635_ (.CLK(clknet_4_14_0_clk),
    .D(_0015_),
    .RESET_B(net37),
    .Q(\seq_div.R[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1636_ (.CLK(clknet_4_15_0_clk),
    .D(_0016_),
    .RESET_B(net37),
    .Q(\seq_div.R[21] ));
 sky130_fd_sc_hd__dfrtp_2 _1637_ (.CLK(clknet_4_15_0_clk),
    .D(_0017_),
    .RESET_B(net37),
    .Q(\seq_div.R[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1638_ (.CLK(clknet_4_12_0_clk),
    .D(_0018_),
    .RESET_B(net37),
    .Q(\seq_div.R[23] ));
 sky130_fd_sc_hd__dfstp_2 _1639_ (.CLK(clknet_4_3_0_clk),
    .D(\osc.next_count[0] ),
    .SET_B(net30),
    .Q(\osc.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1640_ (.CLK(clknet_4_8_0_clk),
    .D(\osc.next_count[1] ),
    .RESET_B(net33),
    .Q(\osc.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1641_ (.CLK(clknet_4_8_0_clk),
    .D(\osc.next_count[2] ),
    .RESET_B(net33),
    .Q(\osc.count[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1642_ (.CLK(clknet_4_8_0_clk),
    .D(\osc.next_count[3] ),
    .RESET_B(net33),
    .Q(\osc.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1643_ (.CLK(clknet_4_8_0_clk),
    .D(\osc.next_count[4] ),
    .RESET_B(net33),
    .Q(\osc.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1644_ (.CLK(clknet_4_8_0_clk),
    .D(\osc.next_count[5] ),
    .RESET_B(net33),
    .Q(\osc.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _1645_ (.CLK(clknet_4_2_0_clk),
    .D(\osc.next_count[6] ),
    .RESET_B(net28),
    .Q(\osc.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1646_ (.CLK(clknet_4_9_0_clk),
    .D(\osc.next_count[7] ),
    .RESET_B(net33),
    .Q(\osc.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1647_ (.CLK(clknet_4_9_0_clk),
    .D(\osc.next_count[8] ),
    .RESET_B(net33),
    .Q(\osc.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1648_ (.CLK(clknet_4_9_0_clk),
    .D(\osc.next_count[9] ),
    .RESET_B(net33),
    .Q(\osc.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1649_ (.CLK(clknet_4_12_0_clk),
    .D(\osc.next_count[10] ),
    .RESET_B(net35),
    .Q(\osc.count[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1650_ (.CLK(clknet_4_3_0_clk),
    .D(\osc.next_count[11] ),
    .RESET_B(net30),
    .Q(\osc.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1651_ (.CLK(clknet_4_3_0_clk),
    .D(\osc.next_count[12] ),
    .RESET_B(net35),
    .Q(\osc.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1652_ (.CLK(clknet_4_3_0_clk),
    .D(\osc.next_count[13] ),
    .RESET_B(net35),
    .Q(\osc.count[13] ));
 sky130_fd_sc_hd__dfrtp_2 _1653_ (.CLK(clknet_4_6_0_clk),
    .D(\osc.next_count[14] ),
    .RESET_B(net35),
    .Q(\osc.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1654_ (.CLK(clknet_4_6_0_clk),
    .D(\osc.next_count[15] ),
    .RESET_B(net35),
    .Q(\osc.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1655_ (.CLK(clknet_4_7_0_clk),
    .D(\clk_div.next_count[0] ),
    .RESET_B(net30),
    .Q(\clk_div.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1656_ (.CLK(clknet_4_6_0_clk),
    .D(net95),
    .RESET_B(net30),
    .Q(\clk_div.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1657_ (.CLK(clknet_4_4_0_clk),
    .D(\clk_div.next_count[2] ),
    .RESET_B(net30),
    .Q(\clk_div.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1658_ (.CLK(clknet_4_4_0_clk),
    .D(\clk_div.next_count[3] ),
    .RESET_B(net30),
    .Q(\clk_div.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1659_ (.CLK(clknet_4_1_0_clk),
    .D(\clk_div.next_count[4] ),
    .RESET_B(net30),
    .Q(\clk_div.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1660_ (.CLK(clknet_4_6_0_clk),
    .D(\clk_div.next_count[5] ),
    .RESET_B(net30),
    .Q(\clk_div.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1661_ (.CLK(clknet_4_6_0_clk),
    .D(\clk_div.next_count[6] ),
    .RESET_B(net30),
    .Q(\clk_div.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1662_ (.CLK(clknet_4_6_0_clk),
    .D(\clk_div.next_count[7] ),
    .RESET_B(net30),
    .Q(\clk_div.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1663_ (.CLK(clknet_4_6_0_clk),
    .D(_0019_),
    .RESET_B(net35),
    .Q(\seq_div.q_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1664_ (.CLK(clknet_4_13_0_clk),
    .D(_0020_),
    .RESET_B(net35),
    .Q(\seq_div.q_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1665_ (.CLK(clknet_4_13_0_clk),
    .D(_0021_),
    .RESET_B(net35),
    .Q(\seq_div.q_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1666_ (.CLK(clknet_4_13_0_clk),
    .D(_0022_),
    .RESET_B(net36),
    .Q(\seq_div.q_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1667_ (.CLK(clknet_4_15_0_clk),
    .D(_0023_),
    .RESET_B(net37),
    .Q(\seq_div.q_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1668_ (.CLK(clknet_4_13_0_clk),
    .D(_0024_),
    .RESET_B(net36),
    .Q(\seq_div.q_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1669_ (.CLK(clknet_4_13_0_clk),
    .D(_0025_),
    .RESET_B(net36),
    .Q(\seq_div.q_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1670_ (.CLK(clknet_4_13_0_clk),
    .D(_0026_),
    .RESET_B(net36),
    .Q(\seq_div.q_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1671_ (.CLK(clknet_4_13_0_clk),
    .D(_0027_),
    .RESET_B(net35),
    .Q(\seq_div.Q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1672_ (.CLK(clknet_4_13_0_clk),
    .D(net82),
    .RESET_B(net36),
    .Q(\seq_div.Q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1673_ (.CLK(clknet_4_13_0_clk),
    .D(net80),
    .RESET_B(net36),
    .Q(\seq_div.Q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1674_ (.CLK(clknet_4_13_0_clk),
    .D(net76),
    .RESET_B(net37),
    .Q(\seq_div.Q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1675_ (.CLK(clknet_4_15_0_clk),
    .D(_0031_),
    .RESET_B(net37),
    .Q(\seq_div.Q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1676_ (.CLK(clknet_4_15_0_clk),
    .D(_0032_),
    .RESET_B(net37),
    .Q(\seq_div.Q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1677_ (.CLK(clknet_4_13_0_clk),
    .D(net63),
    .RESET_B(net36),
    .Q(\seq_div.Q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1678_ (.CLK(clknet_4_13_0_clk),
    .D(net60),
    .RESET_B(net37),
    .Q(\seq_div.Q[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1679_ (.CLK(clknet_4_9_0_clk),
    .D(_0035_),
    .RESET_B(net33),
    .Q(\seq_div.D[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1680_ (.CLK(clknet_4_10_0_clk),
    .D(_0036_),
    .RESET_B(net34),
    .Q(\seq_div.D[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1681_ (.CLK(clknet_4_8_0_clk),
    .D(_0037_),
    .RESET_B(net33),
    .Q(\seq_div.D[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1682_ (.CLK(clknet_4_8_0_clk),
    .D(_0038_),
    .RESET_B(net33),
    .Q(\seq_div.D[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1683_ (.CLK(clknet_4_10_0_clk),
    .D(_0039_),
    .RESET_B(net34),
    .Q(\seq_div.D[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1684_ (.CLK(clknet_4_10_0_clk),
    .D(_0040_),
    .RESET_B(net34),
    .Q(\seq_div.D[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1685_ (.CLK(clknet_4_11_0_clk),
    .D(_0041_),
    .RESET_B(net34),
    .Q(\seq_div.D[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1686_ (.CLK(clknet_4_11_0_clk),
    .D(_0042_),
    .RESET_B(net34),
    .Q(\seq_div.D[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1687_ (.CLK(clknet_4_9_0_clk),
    .D(_0043_),
    .RESET_B(net34),
    .Q(\seq_div.D[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1688_ (.CLK(clknet_4_11_0_clk),
    .D(_0044_),
    .RESET_B(net38),
    .Q(\seq_div.D[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1689_ (.CLK(clknet_4_14_0_clk),
    .D(_0045_),
    .RESET_B(net38),
    .Q(\seq_div.D[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1690_ (.CLK(clknet_4_12_0_clk),
    .D(_0046_),
    .RESET_B(net37),
    .Q(\seq_div.D[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1691_ (.CLK(clknet_4_14_0_clk),
    .D(_0047_),
    .RESET_B(net37),
    .Q(\seq_div.D[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1692_ (.CLK(clknet_4_12_0_clk),
    .D(_0048_),
    .RESET_B(net35),
    .Q(\seq_div.D[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1693_ (.CLK(clknet_4_12_0_clk),
    .D(_0049_),
    .RESET_B(net35),
    .Q(\seq_div.D[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1694_ (.CLK(clknet_4_12_0_clk),
    .D(_0050_),
    .RESET_B(net35),
    .Q(\seq_div.D[15] ));
 sky130_fd_sc_hd__dfrtp_4 _1695_ (.CLK(clknet_4_0_0_clk),
    .D(_0051_),
    .RESET_B(net28),
    .Q(\SS_FSM.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1696_ (.CLK(clknet_4_0_0_clk),
    .D(_0052_),
    .RESET_B(net28),
    .Q(\SS_FSM.count[1] ));
 sky130_fd_sc_hd__dfstp_4 _1697_ (.CLK(clknet_4_1_0_clk),
    .D(_0053_),
    .SET_B(net29),
    .Q(\SS_FSM.count[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1698_ (.CLK(clknet_4_1_0_clk),
    .D(_0054_),
    .RESET_B(net28),
    .Q(\SS_FSM.count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1699_ (.CLK(clknet_4_1_0_clk),
    .D(_0055_),
    .RESET_B(net29),
    .Q(\SS_FSM.count[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1700_ (.CLK(clknet_4_1_0_clk),
    .D(_0056_),
    .RESET_B(net29),
    .Q(\SS_FSM.count[5] ));
 sky130_fd_sc_hd__dfrtp_4 _1701_ (.CLK(clknet_4_1_0_clk),
    .D(_0057_),
    .RESET_B(net30),
    .Q(\SS_FSM.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1702_ (.CLK(clknet_4_4_0_clk),
    .D(_0058_),
    .RESET_B(net29),
    .Q(\SS_FSM.count[7] ));
 sky130_fd_sc_hd__dfstp_1 _1703_ (.CLK(clknet_4_1_0_clk),
    .D(_0059_),
    .SET_B(net29),
    .Q(\SS_FSM.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1704_ (.CLK(clknet_4_8_0_clk),
    .D(_0060_),
    .RESET_B(net33),
    .Q(\seq_div.dividend[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1705_ (.CLK(clknet_4_8_0_clk),
    .D(_0061_),
    .RESET_B(net33),
    .Q(\seq_div.dividend[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1706_ (.CLK(clknet_4_8_0_clk),
    .D(_0062_),
    .RESET_B(net33),
    .Q(\seq_div.dividend[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1707_ (.CLK(clknet_4_8_0_clk),
    .D(_0063_),
    .RESET_B(net33),
    .Q(\seq_div.dividend[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1708_ (.CLK(clknet_4_9_0_clk),
    .D(_0064_),
    .RESET_B(net33),
    .Q(\seq_div.dividend[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1709_ (.CLK(clknet_4_9_0_clk),
    .D(_0065_),
    .RESET_B(net33),
    .Q(\seq_div.dividend[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1710_ (.CLK(clknet_4_11_0_clk),
    .D(_0066_),
    .RESET_B(net38),
    .Q(\seq_div.dividend[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1711_ (.CLK(clknet_4_9_0_clk),
    .D(_0067_),
    .RESET_B(net38),
    .Q(\seq_div.dividend[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1712_ (.CLK(clknet_4_9_0_clk),
    .D(_0068_),
    .RESET_B(net38),
    .Q(\seq_div.dividend[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1713_ (.CLK(clknet_4_9_0_clk),
    .D(_0069_),
    .RESET_B(net38),
    .Q(\seq_div.dividend[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1714_ (.CLK(clknet_4_9_0_clk),
    .D(_0070_),
    .RESET_B(net35),
    .Q(\seq_div.dividend[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1715_ (.CLK(clknet_4_12_0_clk),
    .D(_0071_),
    .RESET_B(net35),
    .Q(\seq_div.dividend[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1716_ (.CLK(clknet_4_12_0_clk),
    .D(_0072_),
    .RESET_B(net35),
    .Q(\seq_div.dividend[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1717_ (.CLK(clknet_4_6_0_clk),
    .D(_0073_),
    .RESET_B(net35),
    .Q(\seq_div.dividend[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1718_ (.CLK(clknet_4_6_0_clk),
    .D(_0074_),
    .RESET_B(net35),
    .Q(\seq_div.dividend[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1719_ (.CLK(clknet_4_12_0_clk),
    .D(_0075_),
    .RESET_B(net35),
    .Q(\seq_div.dividend[15] ));
 sky130_fd_sc_hd__dfrtp_4 _1720_ (.CLK(clknet_4_13_0_clk),
    .D(net74),
    .RESET_B(net38),
    .Q(\seq_div.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1721_ (.CLK(clknet_4_12_0_clk),
    .D(_0077_),
    .RESET_B(net37),
    .Q(\seq_div.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1722_ (.CLK(clknet_4_13_0_clk),
    .D(\pwm.pwm ),
    .RESET_B(net36),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_2 _1723_ (.CLK(clknet_4_6_0_clk),
    .D(\pwm.next_count[0] ),
    .RESET_B(net36),
    .Q(\pwm.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1724_ (.CLK(clknet_4_6_0_clk),
    .D(net72),
    .RESET_B(net31),
    .Q(\pwm.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1725_ (.CLK(clknet_4_7_0_clk),
    .D(\pwm.next_count[2] ),
    .RESET_B(net31),
    .Q(\pwm.count[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1726_ (.CLK(clknet_4_7_0_clk),
    .D(\pwm.next_count[3] ),
    .RESET_B(net31),
    .Q(\pwm.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1727_ (.CLK(clknet_4_7_0_clk),
    .D(\pwm.next_count[4] ),
    .RESET_B(net31),
    .Q(\pwm.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1728_ (.CLK(clknet_4_7_0_clk),
    .D(\pwm.next_count[5] ),
    .RESET_B(net31),
    .Q(\pwm.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1729_ (.CLK(clknet_4_7_0_clk),
    .D(\pwm.next_count[6] ),
    .RESET_B(net31),
    .Q(\pwm.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1730_ (.CLK(clknet_4_7_0_clk),
    .D(\pwm.next_count[7] ),
    .RESET_B(net31),
    .Q(\pwm.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1731_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[0] ),
    .RESET_B(net29),
    .Q(\clk8.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1732_ (.CLK(clknet_4_4_0_clk),
    .D(net66),
    .RESET_B(net29),
    .Q(\clk8.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1733_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[2] ),
    .RESET_B(net29),
    .Q(\clk8.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1734_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[3] ),
    .RESET_B(net29),
    .Q(\clk8.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1735_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[4] ),
    .RESET_B(net29),
    .Q(\clk8.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1736_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[5] ),
    .RESET_B(net29),
    .Q(\clk8.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1737_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[6] ),
    .RESET_B(net29),
    .Q(\clk8.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1738_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[7] ),
    .RESET_B(net29),
    .Q(\clk8.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1739_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[8] ),
    .RESET_B(net29),
    .Q(\clk8.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1740_ (.CLK(clknet_4_4_0_clk),
    .D(\clk8.next_count[9] ),
    .RESET_B(net29),
    .Q(\clk8.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1741_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[10] ),
    .RESET_B(net29),
    .Q(\clk8.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1742_ (.CLK(clknet_4_7_0_clk),
    .D(\clk8.next_count[11] ),
    .RESET_B(net31),
    .Q(\clk8.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1743_ (.CLK(clknet_4_7_0_clk),
    .D(\clk8.next_count[12] ),
    .RESET_B(net31),
    .Q(\clk8.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1744_ (.CLK(clknet_4_5_0_clk),
    .D(net102),
    .RESET_B(net29),
    .Q(\clk8.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1745_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[14] ),
    .RESET_B(net32),
    .Q(\clk8.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1746_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[15] ),
    .RESET_B(net32),
    .Q(\clk8.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1747_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[16] ),
    .RESET_B(net32),
    .Q(\clk8.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1748_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[17] ),
    .RESET_B(net32),
    .Q(\clk8.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1749_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[18] ),
    .RESET_B(net32),
    .Q(\clk8.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1750_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[19] ),
    .RESET_B(net32),
    .Q(\clk8.count[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1751_ (.CLK(clknet_4_5_0_clk),
    .D(\clk8.next_count[20] ),
    .RESET_B(net32),
    .Q(\clk8.count[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1752_ (.CLK(clknet_4_8_0_clk),
    .D(net49),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1753_ (.CLK(clknet_4_2_0_clk),
    .D(net53),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1754_ (.CLK(clknet_4_8_0_clk),
    .D(net48),
    .RESET_B(net33),
    .Q(\kp_encoder.sync_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1755_ (.CLK(clknet_4_2_0_clk),
    .D(net40),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1756_ (.CLK(clknet_4_2_0_clk),
    .D(net39),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1757_ (.CLK(clknet_4_0_0_clk),
    .D(net41),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1758_ (.CLK(clknet_4_2_0_clk),
    .D(net45),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1759_ (.CLK(clknet_4_2_0_clk),
    .D(net44),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1760_ (.CLK(clknet_4_3_0_clk),
    .D(net52),
    .RESET_B(net30),
    .Q(\kp_encoder.sync_out[8] ));
 sky130_fd_sc_hd__dfrtp_2 _1761_ (.CLK(clknet_4_3_0_clk),
    .D(net54),
    .RESET_B(net30),
    .Q(\kp_encoder.sync_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1762_ (.CLK(clknet_4_2_0_clk),
    .D(net42),
    .RESET_B(net28),
    .Q(\kp_encoder.sync_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1763_ (.CLK(clknet_4_3_0_clk),
    .D(net47),
    .RESET_B(net30),
    .Q(\kp_encoder.sync_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1764_ (.CLK(clknet_4_6_0_clk),
    .D(net51),
    .RESET_B(net30),
    .Q(\kp_encoder.sync_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1765_ (.CLK(clknet_4_7_0_clk),
    .D(net43),
    .RESET_B(net31),
    .Q(\kp_encoder.sync_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1766_ (.CLK(clknet_4_15_0_clk),
    .D(net46),
    .RESET_B(net38),
    .Q(\kp_encoder.sync_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1767_ (.CLK(clknet_4_10_0_clk),
    .D(net2),
    .RESET_B(net34),
    .Q(\kp_encoder.q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1768_ (.CLK(clknet_4_10_0_clk),
    .D(net8),
    .RESET_B(net34),
    .Q(\kp_encoder.q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1769_ (.CLK(clknet_4_8_0_clk),
    .D(net9),
    .RESET_B(net28),
    .Q(\kp_encoder.q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1770_ (.CLK(clknet_4_2_0_clk),
    .D(net10),
    .RESET_B(net28),
    .Q(\kp_encoder.q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1771_ (.CLK(clknet_4_0_0_clk),
    .D(net11),
    .RESET_B(net28),
    .Q(\kp_encoder.q[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1772_ (.CLK(clknet_4_7_0_clk),
    .D(_0078_),
    .RESET_B(net36),
    .Q(\mode_FSM.mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1773_ (.CLK(clknet_4_7_0_clk),
    .D(_0079_),
    .RESET_B(net36),
    .Q(\mode_FSM.mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1774_ (.CLK(clknet_4_0_0_clk),
    .D(net12),
    .RESET_B(net28),
    .Q(\kp_encoder.q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1775_ (.CLK(clknet_4_2_0_clk),
    .D(net13),
    .RESET_B(net28),
    .Q(\kp_encoder.q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1776_ (.CLK(clknet_4_2_0_clk),
    .D(net14),
    .RESET_B(net17),
    .Q(\kp_encoder.q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1777_ (.CLK(clknet_4_14_0_clk),
    .D(net15),
    .RESET_B(net37),
    .Q(\kp_encoder.q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1778_ (.CLK(clknet_4_15_0_clk),
    .D(net16),
    .RESET_B(net38),
    .Q(\kp_encoder.q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1779_ (.CLK(clknet_4_0_0_clk),
    .D(net3),
    .RESET_B(net28),
    .Q(\kp_encoder.q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1780_ (.CLK(clknet_4_1_0_clk),
    .D(net4),
    .RESET_B(net29),
    .Q(\kp_encoder.q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1781_ (.CLK(clknet_4_5_0_clk),
    .D(net5),
    .RESET_B(net31),
    .Q(\kp_encoder.q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1782_ (.CLK(clknet_4_7_0_clk),
    .D(net6),
    .RESET_B(net31),
    .Q(\kp_encoder.q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1783_ (.CLK(clknet_4_15_0_clk),
    .D(net7),
    .RESET_B(net38),
    .Q(\kp_encoder.q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1784_ (.CLK(clknet_4_7_0_clk),
    .D(net50),
    .RESET_B(net31),
    .Q(\kp_encoder.last_mk ));
 sky130_fd_sc_hd__dfrtp_1 _1785_ (.CLK(clknet_4_3_0_clk),
    .D(net55),
    .RESET_B(net30),
    .Q(\kp_encoder.last_sk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_6 fanout28 (.A(net17),
    .X(net28));
 sky130_fd_sc_hd__buf_6 fanout29 (.A(net32),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(net32),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__buf_4 fanout32 (.A(net17),
    .X(net32));
 sky130_fd_sc_hd__buf_6 fanout33 (.A(net38),
    .X(net33));
 sky130_fd_sc_hd__buf_6 fanout34 (.A(net38),
    .X(net34));
 sky130_fd_sc_hd__buf_6 fanout35 (.A(net38),
    .X(net35));
 sky130_fd_sc_hd__buf_4 fanout36 (.A(net38),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_8 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net17),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\kp_encoder.q[4] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\kp_encoder.q[2] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\kp_encoder.q[0] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\kp_encoder.sync_out[13] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\kp_encoder.q[12] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\kp_encoder.q[8] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\kp_encoder.q[1] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\kp_encoder.q[9] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\kp_encoder.sync_out[14] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\clk8.count[20] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\seq_div.count_div[2] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\kp_encoder.q[3] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\pwm.count[0] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\seq_div.Q[7] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0034_),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\pwm.count[7] ),
    .X(net61));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold24 (.A(\seq_div.Q[5] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0033_),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\clk_div.count[0] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\clk8.count[1] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\clk8.next_count[1] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\pwm.count[7] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\kp_encoder.q[5] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\seq_div.dividend[0] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0003_),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\clk_div.count[3] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\pwm.count[1] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\pwm.next_count[1] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\seq_div.state[1] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0076_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\seq_div.Q[3] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0030_),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\seq_div.Q[4] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\kp_encoder.q[10] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\seq_div.dividend[6] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\seq_div.Q[2] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0029_),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\seq_div.Q[0] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0028_),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\seq_div.dividend[4] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\seq_div.count_div[1] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0629_),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\seq_div.count_div[0] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\seq_div.D[6] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\kp_encoder.q[13] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\seq_div.dividend[9] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0012_),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\clk8.count[3] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\seq_div.dividend[10] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0013_),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\clk_div.count[4] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\clk_div.count[1] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\clk_div.next_count[1] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\seq_div.dividend[2] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\osc.count[0] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\kp_encoder.q[7] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\seq_div.dividend[7] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\seq_div.dividend[8] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0011_),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\clk8.count[13] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\clk8.next_count[13] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\clk8.count[4] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\seq_div.D[0] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\clk8.count[16] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\clk8.count[7] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\seq_div.dividend[5] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\kp_encoder.q[6] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\seq_div.R[23] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0775_),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\clk8.count[10] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\seq_div.dividend[14] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\SS_FSM.count[7] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\seq_div.dividend[1] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\seq_div.dividend[13] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\seq_div.D[12] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\SS_FSM.count[8] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\seq_div.dividend[11] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\kp_encoder.q[14] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\seq_div.D[5] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\seq_div.D[10] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\seq_div.Q[0] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\seq_div.Q[4] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\seq_div.Q[3] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\seq_div.dividend[0] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\seq_div.dividend[4] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\seq_div.dividend[11] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\seq_div.dividend[1] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\seq_div.dividend[5] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\kp_encoder.q[11] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\seq_div.dividend[2] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\seq_div.dividend[13] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\seq_div.dividend[14] ),
    .X(net130));
 sky130_fd_sc_hd__buf_4 input1 (.A(en),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(keypad_i[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(keypad_i[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(keypad_i[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(keypad_i[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(keypad_i[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(keypad_i[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(keypad_i[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(n_rst),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(keypad_i[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(keypad_i[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(keypad_i[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(keypad_i[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(keypad_i[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(keypad_i[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(keypad_i[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(keypad_i[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap23 (.A(_0120_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 max_cap24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 max_cap25 (.A(_0157_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 max_cap26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 max_cap27 (.A(_0163_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(pwm_o));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(sound_series[0]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(sound_series[1]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(sound_series[2]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(sound_series[3]));
endmodule

