magic
tech sky130A
magscale 1 2
timestamp 1694100622
<< obsli1 >>
rect 1104 2159 274160 274737
<< obsm1 >>
rect 14 2128 275066 274768
<< metal2 >>
rect 5814 276622 5870 277422
rect 39946 276622 40002 277422
rect 73434 276622 73490 277422
rect 106922 276622 106978 277422
rect 140410 276622 140466 277422
rect 174542 276622 174598 277422
rect 208030 276622 208086 277422
rect 241518 276622 241574 277422
rect 275006 276622 275062 277422
rect 18 0 74 800
rect 33506 0 33562 800
rect 66994 0 67050 800
rect 100482 0 100538 800
rect 134614 0 134670 800
rect 168102 0 168158 800
rect 201590 0 201646 800
rect 235078 0 235134 800
rect 269210 0 269266 800
<< obsm2 >>
rect 20 276566 5758 276622
rect 5926 276566 39890 276622
rect 40058 276566 73378 276622
rect 73546 276566 106866 276622
rect 107034 276566 140354 276622
rect 140522 276566 174486 276622
rect 174654 276566 207974 276622
rect 208142 276566 241462 276622
rect 241630 276566 274950 276622
rect 20 856 275060 276566
rect 130 734 33450 856
rect 33618 734 66938 856
rect 67106 734 100426 856
rect 100594 734 134558 856
rect 134726 734 168046 856
rect 168214 734 201534 856
rect 201702 734 235022 856
rect 235190 734 269154 856
rect 269322 734 275060 856
<< metal3 >>
rect 0 248208 800 248328
rect 274478 241408 275278 241528
rect 0 212848 800 212968
rect 274478 206048 275278 206168
rect 0 177488 800 177608
rect 274478 170688 275278 170808
rect 0 141448 800 141568
rect 274478 135328 275278 135448
rect 0 106088 800 106208
rect 274478 99288 275278 99408
rect 0 70728 800 70848
rect 274478 63928 275278 64048
rect 0 35368 800 35488
rect 274478 28568 275278 28688
<< obsm3 >>
rect 800 248408 274478 274753
rect 880 248128 274478 248408
rect 800 241608 274478 248128
rect 800 241328 274398 241608
rect 800 213048 274478 241328
rect 880 212768 274478 213048
rect 800 206248 274478 212768
rect 800 205968 274398 206248
rect 800 177688 274478 205968
rect 880 177408 274478 177688
rect 800 170888 274478 177408
rect 800 170608 274398 170888
rect 800 141648 274478 170608
rect 880 141368 274478 141648
rect 800 135528 274478 141368
rect 800 135248 274398 135528
rect 800 106288 274478 135248
rect 880 106008 274478 106288
rect 800 99488 274478 106008
rect 800 99208 274398 99488
rect 800 70928 274478 99208
rect 880 70648 274478 70928
rect 800 64128 274478 70648
rect 800 63848 274398 64128
rect 800 35568 274478 63848
rect 880 35288 274478 35568
rect 800 28768 274478 35288
rect 800 28488 274398 28768
rect 800 2143 274478 28488
<< metal4 >>
rect 4208 2128 4528 274768
rect 19568 2128 19888 274768
rect 34928 2128 35248 274768
rect 50288 2128 50608 274768
rect 65648 2128 65968 274768
rect 81008 2128 81328 274768
rect 96368 2128 96688 274768
rect 111728 2128 112048 274768
rect 127088 2128 127408 274768
rect 142448 2128 142768 274768
rect 157808 2128 158128 274768
rect 173168 2128 173488 274768
rect 188528 2128 188848 274768
rect 203888 2128 204208 274768
rect 219248 2128 219568 274768
rect 234608 2128 234928 274768
rect 249968 2128 250288 274768
rect 265328 2128 265648 274768
<< obsm4 >>
rect 62619 2347 65568 273325
rect 66048 2347 80928 273325
rect 81408 2347 96288 273325
rect 96768 2347 111648 273325
rect 112128 2347 127008 273325
rect 127488 2347 142368 273325
rect 142848 2347 157728 273325
rect 158208 2347 173088 273325
rect 173568 2347 188448 273325
rect 188928 2347 203808 273325
rect 204288 2347 205837 273325
<< labels >>
rlabel metal2 s 275006 276622 275062 277422 6 clk
port 1 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 color[0]
port 2 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 color[10]
port 3 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 color[11]
port 4 nsew signal output
rlabel metal2 s 73434 276622 73490 277422 6 color[12]
port 5 nsew signal output
rlabel metal2 s 174542 276622 174598 277422 6 color[13]
port 6 nsew signal output
rlabel metal2 s 235078 0 235134 800 6 color[14]
port 7 nsew signal output
rlabel metal3 s 274478 135328 275278 135448 6 color[15]
port 8 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 color[16]
port 9 nsew signal output
rlabel metal3 s 274478 170688 275278 170808 6 color[17]
port 10 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 color[18]
port 11 nsew signal output
rlabel metal2 s 18 0 74 800 6 color[19]
port 12 nsew signal output
rlabel metal2 s 208030 276622 208086 277422 6 color[1]
port 13 nsew signal output
rlabel metal2 s 241518 276622 241574 277422 6 color[20]
port 14 nsew signal output
rlabel metal3 s 0 177488 800 177608 6 color[21]
port 15 nsew signal output
rlabel metal3 s 274478 28568 275278 28688 6 color[22]
port 16 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 color[23]
port 17 nsew signal output
rlabel metal3 s 0 248208 800 248328 6 color[2]
port 18 nsew signal output
rlabel metal2 s 269210 0 269266 800 6 color[3]
port 19 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 color[4]
port 20 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 color[5]
port 21 nsew signal output
rlabel metal2 s 39946 276622 40002 277422 6 color[6]
port 22 nsew signal output
rlabel metal3 s 274478 63928 275278 64048 6 color[7]
port 23 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 color[8]
port 24 nsew signal output
rlabel metal3 s 274478 206048 275278 206168 6 color[9]
port 25 nsew signal output
rlabel metal3 s 274478 241408 275278 241528 6 cs
port 26 nsew signal input
rlabel metal2 s 106922 276622 106978 277422 6 is_mandelbrot
port 27 nsew signal output
rlabel metal2 s 140410 276622 140466 277422 6 nrst
port 28 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 spi_clk
port 29 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 spi_data
port 30 nsew signal input
rlabel metal2 s 5814 276622 5870 277422 6 spi_en
port 31 nsew signal input
rlabel metal3 s 274478 99288 275278 99408 6 valid_out
port 32 nsew signal output
rlabel metal4 s 4208 2128 4528 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 274768 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 274768 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 274768 6 vssd1
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 275278 277422
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 80376776
string GDS_FILE /home/designer-05/Caravel_STARS_2023/openlane/DigiDoggs/runs/23_09_07_07_52/results/signoff/pushing_pixels.magic.gds
string GDS_START 1573262
<< end >>

