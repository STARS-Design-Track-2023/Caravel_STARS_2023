// This is the unpowered netlist.
module Synthia (PWM_o,
    clk,
    modes,
    octaves,
    reset,
    pb);
 output PWM_o;
 input clk;
 input modes;
 input octaves;
 input reset;
 input [12:0] pb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \d1.count[0] ;
 wire \d1.count[1] ;
 wire \d1.count[2] ;
 wire \d1.count[3] ;
 wire \d1.count[4] ;
 wire \d1.count[5] ;
 wire \d1.count[6] ;
 wire \d1.count[7] ;
 wire \d1.count[8] ;
 wire \d1.count[9] ;
 wire \d1.nxt_count[0] ;
 wire \d1.nxt_count[1] ;
 wire \d1.nxt_count[2] ;
 wire \d1.nxt_count[3] ;
 wire \d1.nxt_count[4] ;
 wire \d1.nxt_count[5] ;
 wire \d1.nxt_count[6] ;
 wire \d1.nxt_count[7] ;
 wire \d1.nxt_count[8] ;
 wire \d1.nxt_count[9] ;
 wire \d1.oct_dwn[0] ;
 wire \d1.oct_dwn[1] ;
 wire \d1.saw_temp[0] ;
 wire \d1.saw_temp[1] ;
 wire \d1.saw_temp[2] ;
 wire \d1.saw_temp[3] ;
 wire \d1.saw_temp[4] ;
 wire \d1.saw_temp[5] ;
 wire \d1.saw_temp[6] ;
 wire \d1.saw_temp[7] ;
 wire \d10.count[0] ;
 wire \d10.count[1] ;
 wire \d10.count[2] ;
 wire \d10.count[3] ;
 wire \d10.count[4] ;
 wire \d10.count[5] ;
 wire \d10.count[6] ;
 wire \d10.count[7] ;
 wire \d10.count[8] ;
 wire \d10.count[9] ;
 wire \d10.nxt_count[0] ;
 wire \d10.nxt_count[1] ;
 wire \d10.nxt_count[2] ;
 wire \d10.nxt_count[3] ;
 wire \d10.nxt_count[4] ;
 wire \d10.nxt_count[5] ;
 wire \d10.nxt_count[6] ;
 wire \d10.nxt_count[7] ;
 wire \d10.nxt_count[8] ;
 wire \d10.saw_temp[0] ;
 wire \d10.saw_temp[1] ;
 wire \d10.saw_temp[2] ;
 wire \d10.saw_temp[3] ;
 wire \d10.saw_temp[4] ;
 wire \d10.saw_temp[5] ;
 wire \d10.saw_temp[6] ;
 wire \d10.saw_temp[7] ;
 wire \d11.count[0] ;
 wire \d11.count[1] ;
 wire \d11.count[2] ;
 wire \d11.count[3] ;
 wire \d11.count[4] ;
 wire \d11.count[5] ;
 wire \d11.count[6] ;
 wire \d11.count[7] ;
 wire \d11.count[8] ;
 wire \d11.count[9] ;
 wire \d11.nxt_count[0] ;
 wire \d11.nxt_count[1] ;
 wire \d11.nxt_count[2] ;
 wire \d11.nxt_count[3] ;
 wire \d11.nxt_count[4] ;
 wire \d11.nxt_count[5] ;
 wire \d11.nxt_count[6] ;
 wire \d11.nxt_count[7] ;
 wire \d11.nxt_count[8] ;
 wire \d11.saw_temp[0] ;
 wire \d11.saw_temp[1] ;
 wire \d11.saw_temp[2] ;
 wire \d11.saw_temp[3] ;
 wire \d11.saw_temp[4] ;
 wire \d11.saw_temp[5] ;
 wire \d11.saw_temp[6] ;
 wire \d11.saw_temp[7] ;
 wire \d12.count[0] ;
 wire \d12.count[1] ;
 wire \d12.count[2] ;
 wire \d12.count[3] ;
 wire \d12.count[4] ;
 wire \d12.count[5] ;
 wire \d12.count[6] ;
 wire \d12.count[7] ;
 wire \d12.count[8] ;
 wire \d12.count[9] ;
 wire \d12.nxt_count[0] ;
 wire \d12.nxt_count[1] ;
 wire \d12.nxt_count[2] ;
 wire \d12.nxt_count[3] ;
 wire \d12.nxt_count[4] ;
 wire \d12.nxt_count[5] ;
 wire \d12.nxt_count[6] ;
 wire \d12.nxt_count[7] ;
 wire \d12.nxt_count[8] ;
 wire \d12.saw_temp[0] ;
 wire \d12.saw_temp[1] ;
 wire \d12.saw_temp[2] ;
 wire \d12.saw_temp[3] ;
 wire \d12.saw_temp[4] ;
 wire \d12.saw_temp[5] ;
 wire \d12.saw_temp[6] ;
 wire \d12.saw_temp[7] ;
 wire \d13.count[0] ;
 wire \d13.count[1] ;
 wire \d13.count[2] ;
 wire \d13.count[3] ;
 wire \d13.count[4] ;
 wire \d13.count[5] ;
 wire \d13.count[6] ;
 wire \d13.count[7] ;
 wire \d13.count[8] ;
 wire \d13.count[9] ;
 wire \d13.nxt_count[0] ;
 wire \d13.nxt_count[1] ;
 wire \d13.nxt_count[2] ;
 wire \d13.nxt_count[3] ;
 wire \d13.nxt_count[4] ;
 wire \d13.nxt_count[5] ;
 wire \d13.nxt_count[6] ;
 wire \d13.nxt_count[7] ;
 wire \d13.nxt_count[8] ;
 wire \d13.saw_temp[0] ;
 wire \d13.saw_temp[1] ;
 wire \d13.saw_temp[2] ;
 wire \d13.saw_temp[3] ;
 wire \d13.saw_temp[4] ;
 wire \d13.saw_temp[5] ;
 wire \d13.saw_temp[6] ;
 wire \d13.saw_temp[7] ;
 wire \d2.count[0] ;
 wire \d2.count[1] ;
 wire \d2.count[2] ;
 wire \d2.count[3] ;
 wire \d2.count[4] ;
 wire \d2.count[5] ;
 wire \d2.count[6] ;
 wire \d2.count[7] ;
 wire \d2.count[8] ;
 wire \d2.count[9] ;
 wire \d2.nxt_count[0] ;
 wire \d2.nxt_count[1] ;
 wire \d2.nxt_count[2] ;
 wire \d2.nxt_count[3] ;
 wire \d2.nxt_count[4] ;
 wire \d2.nxt_count[5] ;
 wire \d2.nxt_count[6] ;
 wire \d2.nxt_count[7] ;
 wire \d2.nxt_count[8] ;
 wire \d2.nxt_count[9] ;
 wire \d2.saw_temp[0] ;
 wire \d2.saw_temp[1] ;
 wire \d2.saw_temp[2] ;
 wire \d2.saw_temp[3] ;
 wire \d2.saw_temp[4] ;
 wire \d2.saw_temp[5] ;
 wire \d2.saw_temp[6] ;
 wire \d2.saw_temp[7] ;
 wire \d3.count[0] ;
 wire \d3.count[1] ;
 wire \d3.count[2] ;
 wire \d3.count[3] ;
 wire \d3.count[4] ;
 wire \d3.count[5] ;
 wire \d3.count[6] ;
 wire \d3.count[7] ;
 wire \d3.count[8] ;
 wire \d3.count[9] ;
 wire \d3.nxt_count[0] ;
 wire \d3.nxt_count[1] ;
 wire \d3.nxt_count[2] ;
 wire \d3.nxt_count[3] ;
 wire \d3.nxt_count[4] ;
 wire \d3.nxt_count[5] ;
 wire \d3.nxt_count[6] ;
 wire \d3.nxt_count[7] ;
 wire \d3.nxt_count[8] ;
 wire \d3.nxt_count[9] ;
 wire \d3.saw_temp[0] ;
 wire \d3.saw_temp[1] ;
 wire \d3.saw_temp[2] ;
 wire \d3.saw_temp[3] ;
 wire \d3.saw_temp[4] ;
 wire \d3.saw_temp[5] ;
 wire \d3.saw_temp[6] ;
 wire \d3.saw_temp[7] ;
 wire \d4.count[0] ;
 wire \d4.count[1] ;
 wire \d4.count[2] ;
 wire \d4.count[3] ;
 wire \d4.count[4] ;
 wire \d4.count[5] ;
 wire \d4.count[6] ;
 wire \d4.count[7] ;
 wire \d4.count[8] ;
 wire \d4.count[9] ;
 wire \d4.nxt_count[0] ;
 wire \d4.nxt_count[1] ;
 wire \d4.nxt_count[2] ;
 wire \d4.nxt_count[3] ;
 wire \d4.nxt_count[4] ;
 wire \d4.nxt_count[5] ;
 wire \d4.nxt_count[6] ;
 wire \d4.nxt_count[7] ;
 wire \d4.nxt_count[8] ;
 wire \d4.saw_temp[0] ;
 wire \d4.saw_temp[1] ;
 wire \d4.saw_temp[2] ;
 wire \d4.saw_temp[3] ;
 wire \d4.saw_temp[4] ;
 wire \d4.saw_temp[5] ;
 wire \d4.saw_temp[6] ;
 wire \d4.saw_temp[7] ;
 wire \d5.count[0] ;
 wire \d5.count[1] ;
 wire \d5.count[2] ;
 wire \d5.count[3] ;
 wire \d5.count[4] ;
 wire \d5.count[5] ;
 wire \d5.count[6] ;
 wire \d5.count[7] ;
 wire \d5.count[8] ;
 wire \d5.count[9] ;
 wire \d5.nxt_count[0] ;
 wire \d5.nxt_count[1] ;
 wire \d5.nxt_count[2] ;
 wire \d5.nxt_count[3] ;
 wire \d5.nxt_count[4] ;
 wire \d5.nxt_count[5] ;
 wire \d5.nxt_count[6] ;
 wire \d5.nxt_count[7] ;
 wire \d5.nxt_count[8] ;
 wire \d5.saw_temp[0] ;
 wire \d5.saw_temp[1] ;
 wire \d5.saw_temp[2] ;
 wire \d5.saw_temp[3] ;
 wire \d5.saw_temp[4] ;
 wire \d5.saw_temp[5] ;
 wire \d5.saw_temp[6] ;
 wire \d5.saw_temp[7] ;
 wire \d6.count[0] ;
 wire \d6.count[1] ;
 wire \d6.count[2] ;
 wire \d6.count[3] ;
 wire \d6.count[4] ;
 wire \d6.count[5] ;
 wire \d6.count[6] ;
 wire \d6.count[7] ;
 wire \d6.count[8] ;
 wire \d6.count[9] ;
 wire \d6.nxt_count[0] ;
 wire \d6.nxt_count[1] ;
 wire \d6.nxt_count[2] ;
 wire \d6.nxt_count[3] ;
 wire \d6.nxt_count[4] ;
 wire \d6.nxt_count[5] ;
 wire \d6.nxt_count[6] ;
 wire \d6.nxt_count[7] ;
 wire \d6.nxt_count[8] ;
 wire \d6.saw_temp[0] ;
 wire \d6.saw_temp[1] ;
 wire \d6.saw_temp[2] ;
 wire \d6.saw_temp[3] ;
 wire \d6.saw_temp[4] ;
 wire \d6.saw_temp[5] ;
 wire \d6.saw_temp[6] ;
 wire \d6.saw_temp[7] ;
 wire \d7.count[0] ;
 wire \d7.count[1] ;
 wire \d7.count[2] ;
 wire \d7.count[3] ;
 wire \d7.count[4] ;
 wire \d7.count[5] ;
 wire \d7.count[6] ;
 wire \d7.count[7] ;
 wire \d7.count[8] ;
 wire \d7.count[9] ;
 wire \d7.nxt_count[0] ;
 wire \d7.nxt_count[1] ;
 wire \d7.nxt_count[2] ;
 wire \d7.nxt_count[3] ;
 wire \d7.nxt_count[4] ;
 wire \d7.nxt_count[5] ;
 wire \d7.nxt_count[6] ;
 wire \d7.nxt_count[7] ;
 wire \d7.nxt_count[8] ;
 wire \d7.saw_temp[0] ;
 wire \d7.saw_temp[1] ;
 wire \d7.saw_temp[2] ;
 wire \d7.saw_temp[3] ;
 wire \d7.saw_temp[4] ;
 wire \d7.saw_temp[5] ;
 wire \d7.saw_temp[6] ;
 wire \d7.saw_temp[7] ;
 wire \d8.count[0] ;
 wire \d8.count[1] ;
 wire \d8.count[2] ;
 wire \d8.count[3] ;
 wire \d8.count[4] ;
 wire \d8.count[5] ;
 wire \d8.count[6] ;
 wire \d8.count[7] ;
 wire \d8.count[8] ;
 wire \d8.count[9] ;
 wire \d8.nxt_count[0] ;
 wire \d8.nxt_count[1] ;
 wire \d8.nxt_count[2] ;
 wire \d8.nxt_count[3] ;
 wire \d8.nxt_count[4] ;
 wire \d8.nxt_count[5] ;
 wire \d8.nxt_count[6] ;
 wire \d8.nxt_count[7] ;
 wire \d8.nxt_count[8] ;
 wire \d8.saw_temp[0] ;
 wire \d8.saw_temp[1] ;
 wire \d8.saw_temp[2] ;
 wire \d8.saw_temp[3] ;
 wire \d8.saw_temp[4] ;
 wire \d8.saw_temp[5] ;
 wire \d8.saw_temp[6] ;
 wire \d8.saw_temp[7] ;
 wire \d9.count[0] ;
 wire \d9.count[1] ;
 wire \d9.count[2] ;
 wire \d9.count[3] ;
 wire \d9.count[4] ;
 wire \d9.count[5] ;
 wire \d9.count[6] ;
 wire \d9.count[7] ;
 wire \d9.count[8] ;
 wire \d9.count[9] ;
 wire \d9.nxt_count[0] ;
 wire \d9.nxt_count[1] ;
 wire \d9.nxt_count[2] ;
 wire \d9.nxt_count[3] ;
 wire \d9.nxt_count[4] ;
 wire \d9.nxt_count[5] ;
 wire \d9.nxt_count[6] ;
 wire \d9.nxt_count[7] ;
 wire \d9.nxt_count[8] ;
 wire \d9.saw_temp[0] ;
 wire \d9.saw_temp[1] ;
 wire \d9.saw_temp[2] ;
 wire \d9.saw_temp[3] ;
 wire \d9.saw_temp[4] ;
 wire \d9.saw_temp[5] ;
 wire \d9.saw_temp[6] ;
 wire \d9.saw_temp[7] ;
 wire \e0.next_q[0] ;
 wire \e0.next_q[1] ;
 wire \em0.mixed_sample[0] ;
 wire \em0.mixed_sample[1] ;
 wire \em0.mixed_sample[2] ;
 wire \em0.mixed_sample[3] ;
 wire \em0.mixed_sample[4] ;
 wire \em0.mixed_sample[5] ;
 wire \em0.mixed_sample[6] ;
 wire \em0.mixed_sample[7] ;
 wire \em0.u1.D[10] ;
 wire \em0.u1.D[11] ;
 wire \em0.u1.D[12] ;
 wire \em0.u1.D[8] ;
 wire \em0.u1.D[9] ;
 wire \em0.u1.Q[0] ;
 wire \em0.u1.Q[1] ;
 wire \em0.u1.Q[2] ;
 wire \em0.u1.Q[3] ;
 wire \em0.u1.Q[4] ;
 wire \em0.u1.Q[5] ;
 wire \em0.u1.Q[6] ;
 wire \em0.u1.Q[7] ;
 wire \em0.u1.R[10] ;
 wire \em0.u1.R[11] ;
 wire \em0.u1.R[12] ;
 wire \em0.u1.R[13] ;
 wire \em0.u1.R[14] ;
 wire \em0.u1.R[15] ;
 wire \em0.u1.R[16] ;
 wire \em0.u1.R[17] ;
 wire \em0.u1.R[18] ;
 wire \em0.u1.R[19] ;
 wire \em0.u1.R[20] ;
 wire \em0.u1.R[21] ;
 wire \em0.u1.R[22] ;
 wire \em0.u1.R[8] ;
 wire \em0.u1.R[9] ;
 wire \em0.u1.count[0] ;
 wire \em0.u1.count[1] ;
 wire \em0.u1.count[2] ;
 wire \em0.u1.state[0] ;
 wire \em0.u1.state[1] ;
 wire \em0.u1.state[2] ;
 wire \em0.u1.state[3] ;
 wire \m0.edgo.delay ;
 wire \m0.edgo.in ;
 wire \m0.edgy.delay ;
 wire \m0.edgy.in ;
 wire \m0.synco.delay ;
 wire \m0.syncy.delay ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \p0.count[0] ;
 wire \p0.count[1] ;
 wire \p0.count[2] ;
 wire \p0.count[3] ;
 wire \p0.count[4] ;
 wire \p0.count[5] ;
 wire \p0.count[6] ;
 wire \p0.count[7] ;
 wire \p0.nxt_count[0] ;
 wire \p0.nxt_count[1] ;
 wire \p0.nxt_count[2] ;
 wire \p0.nxt_count[3] ;
 wire \p0.nxt_count[4] ;
 wire \p0.nxt_count[5] ;
 wire \p0.nxt_count[6] ;
 wire \p0.nxt_count[7] ;
 wire \p0.pwm ;
 wire \s0.next_q[0] ;
 wire \s0.next_q[1] ;
 wire \s0.type_switch[0] ;
 wire \s0.type_switch[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0738_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_92 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__or2_1 _2030_ (.A(\em0.u1.state[3] ),
    .B(\em0.u1.state[0] ),
    .X(_1709_));
 sky130_fd_sc_hd__clkbuf_1 _2031_ (.A(_1709_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_8 _2032_ (.A(\em0.u1.state[1] ),
    .X(_1710_));
 sky130_fd_sc_hd__nand3_1 _2033_ (.A(net102),
    .B(\em0.u1.count[1] ),
    .C(net60),
    .Y(_1711_));
 sky130_fd_sc_hd__a21o_1 _2034_ (.A1(_1710_),
    .A2(_1711_),
    .B1(net245),
    .X(_0001_));
 sky130_fd_sc_hd__clkbuf_8 _2035_ (.A(\d1.oct_dwn[1] ),
    .X(_1712_));
 sky130_fd_sc_hd__buf_6 _2036_ (.A(\d1.oct_dwn[0] ),
    .X(_1713_));
 sky130_fd_sc_hd__nand2_4 _2037_ (.A(_1712_),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__buf_6 _2038_ (.A(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__inv_2 _2039_ (.A(_1713_),
    .Y(_1716_));
 sky130_fd_sc_hd__nand2_1 _2040_ (.A(_1712_),
    .B(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hd__buf_6 _2041_ (.A(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__a22o_1 _2042_ (.A1(\d1.count[9] ),
    .A2(_1715_),
    .B1(_1718_),
    .B2(\d1.count[8] ),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_8 _2043_ (.A(_1718_),
    .X(_1720_));
 sky130_fd_sc_hd__inv_6 _2044_ (.A(_1712_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_2 _2045_ (.A(_1721_),
    .B(_1713_),
    .Y(_1722_));
 sky130_fd_sc_hd__buf_6 _2046_ (.A(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__nor2_8 _2047_ (.A(_1721_),
    .B(_1716_),
    .Y(_1724_));
 sky130_fd_sc_hd__nor2_4 _2048_ (.A(_1712_),
    .B(_1713_),
    .Y(_1725_));
 sky130_fd_sc_hd__nor2_4 _2049_ (.A(_1724_),
    .B(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__buf_6 _2050_ (.A(_1716_),
    .X(_1727_));
 sky130_fd_sc_hd__a22o_1 _2051_ (.A1(_1727_),
    .A2(\d1.count[4] ),
    .B1(_1718_),
    .B2(\d1.count[5] ),
    .X(_1728_));
 sky130_fd_sc_hd__nor2_2 _2052_ (.A(_1712_),
    .B(_1727_),
    .Y(_1729_));
 sky130_fd_sc_hd__o21ai_1 _2053_ (.A1(\d1.count[2] ),
    .A2(_1729_),
    .B1(\d1.count[3] ),
    .Y(_1730_));
 sky130_fd_sc_hd__or2_1 _2054_ (.A(_1712_),
    .B(_1713_),
    .X(_1731_));
 sky130_fd_sc_hd__buf_4 _2055_ (.A(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2_8 _2056_ (.A(_1714_),
    .B(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__o21a_1 _2057_ (.A1(_1713_),
    .A2(\d1.count[0] ),
    .B1(\d1.count[1] ),
    .X(_1734_));
 sky130_fd_sc_hd__buf_6 _2058_ (.A(_1712_),
    .X(_1735_));
 sky130_fd_sc_hd__o22a_1 _2059_ (.A1(\d1.count[3] ),
    .A2(_1729_),
    .B1(_1734_),
    .B2(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__o21ai_1 _2060_ (.A1(\d1.count[2] ),
    .A2(_1733_),
    .B1(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__nor2_1 _2061_ (.A(_1727_),
    .B(\d1.count[4] ),
    .Y(_1738_));
 sky130_fd_sc_hd__a21oi_1 _2062_ (.A1(_1730_),
    .A2(_1737_),
    .B1(_1738_),
    .Y(_1739_));
 sky130_fd_sc_hd__or2_1 _2063_ (.A(\d1.count[6] ),
    .B(_1726_),
    .X(_1740_));
 sky130_fd_sc_hd__o221a_1 _2064_ (.A1(\d1.count[5] ),
    .A2(_1720_),
    .B1(_1728_),
    .B2(_1739_),
    .C1(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__a221o_1 _2065_ (.A1(\d1.count[7] ),
    .A2(_1723_),
    .B1(_1726_),
    .B2(\d1.count[6] ),
    .C1(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__o221a_1 _2066_ (.A1(\d1.count[8] ),
    .A2(_1720_),
    .B1(_1723_),
    .B2(\d1.count[7] ),
    .C1(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__inv_2 _2067_ (.A(\d1.count[9] ),
    .Y(_1744_));
 sky130_fd_sc_hd__a2bb2o_2 _2068_ (.A1_N(_1719_),
    .A2_N(_1743_),
    .B1(_1744_),
    .B2(_1724_),
    .X(_1745_));
 sky130_fd_sc_hd__nand2_1 _2069_ (.A(net80),
    .B(_1745_),
    .Y(\d1.nxt_count[0] ));
 sky130_fd_sc_hd__nand2_1 _2070_ (.A(\d1.count[0] ),
    .B(\d1.count[1] ),
    .Y(_1746_));
 sky130_fd_sc_hd__or2_1 _2071_ (.A(\d1.count[0] ),
    .B(\d1.count[1] ),
    .X(_1747_));
 sky130_fd_sc_hd__and3_1 _2072_ (.A(_1745_),
    .B(_1746_),
    .C(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__clkbuf_1 _2073_ (.A(_1748_),
    .X(\d1.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2074_ (.A(\d1.count[0] ),
    .B(\d1.count[1] ),
    .C(\d1.count[2] ),
    .X(_1749_));
 sky130_fd_sc_hd__inv_2 _2075_ (.A(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__a21o_1 _2076_ (.A1(\d1.count[0] ),
    .A2(\d1.count[1] ),
    .B1(\d1.count[2] ),
    .X(_1751_));
 sky130_fd_sc_hd__and3_1 _2077_ (.A(_1745_),
    .B(_1750_),
    .C(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__clkbuf_1 _2078_ (.A(_1752_),
    .X(\d1.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2079_ (.A(\d1.count[3] ),
    .B(_1749_),
    .X(_1753_));
 sky130_fd_sc_hd__o21ai_1 _2080_ (.A1(net213),
    .A2(_1749_),
    .B1(_1745_),
    .Y(_1754_));
 sky130_fd_sc_hd__nor2_1 _2081_ (.A(_1753_),
    .B(_1754_),
    .Y(\d1.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2082_ (.A(\d1.count[3] ),
    .B(\d1.count[4] ),
    .C(_1749_),
    .X(_1755_));
 sky130_fd_sc_hd__o21ai_1 _2083_ (.A1(net250),
    .A2(_1753_),
    .B1(_1745_),
    .Y(_1756_));
 sky130_fd_sc_hd__nor2_1 _2084_ (.A(_1755_),
    .B(_1756_),
    .Y(\d1.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2085_ (.A(\d1.count[5] ),
    .B(\d1.count[4] ),
    .C(_1753_),
    .X(_1757_));
 sky130_fd_sc_hd__o21ai_1 _2086_ (.A1(net230),
    .A2(_1755_),
    .B1(_1745_),
    .Y(_1758_));
 sky130_fd_sc_hd__nor2_1 _2087_ (.A(_1757_),
    .B(_1758_),
    .Y(\d1.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2088_ (.A(\d1.count[6] ),
    .B(_1757_),
    .X(_1759_));
 sky130_fd_sc_hd__o21ai_1 _2089_ (.A1(net238),
    .A2(_1757_),
    .B1(_1745_),
    .Y(_1760_));
 sky130_fd_sc_hd__nor2_1 _2090_ (.A(_1759_),
    .B(_1760_),
    .Y(\d1.nxt_count[6] ));
 sky130_fd_sc_hd__and3_1 _2091_ (.A(\d1.count[7] ),
    .B(\d1.count[6] ),
    .C(_1757_),
    .X(_1761_));
 sky130_fd_sc_hd__o21ai_1 _2092_ (.A1(\d1.count[7] ),
    .A2(_1759_),
    .B1(_1745_),
    .Y(_1762_));
 sky130_fd_sc_hd__nor2_1 _2093_ (.A(_1761_),
    .B(_1762_),
    .Y(\d1.nxt_count[7] ));
 sky130_fd_sc_hd__o21ai_1 _2094_ (.A1(\d1.count[8] ),
    .A2(_1761_),
    .B1(_1745_),
    .Y(_1763_));
 sky130_fd_sc_hd__a21oi_1 _2095_ (.A1(net109),
    .A2(_1761_),
    .B1(_1763_),
    .Y(\d1.nxt_count[8] ));
 sky130_fd_sc_hd__a21o_1 _2096_ (.A1(\d1.count[8] ),
    .A2(_1761_),
    .B1(\d1.count[9] ),
    .X(_1764_));
 sky130_fd_sc_hd__nand3_1 _2097_ (.A(\d1.count[9] ),
    .B(\d1.count[8] ),
    .C(_1761_),
    .Y(_1765_));
 sky130_fd_sc_hd__and3_1 _2098_ (.A(_1745_),
    .B(_1764_),
    .C(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__clkbuf_1 _2099_ (.A(_1766_),
    .X(\d1.nxt_count[9] ));
 sky130_fd_sc_hd__a22o_1 _2100_ (.A1(\d2.count[9] ),
    .A2(_1714_),
    .B1(_1718_),
    .B2(\d2.count[8] ),
    .X(_1767_));
 sky130_fd_sc_hd__nand2_1 _2101_ (.A(\d2.count[7] ),
    .B(_1722_),
    .Y(_1768_));
 sky130_fd_sc_hd__o21a_1 _2102_ (.A1(_1713_),
    .A2(\d2.count[1] ),
    .B1(\d2.count[2] ),
    .X(_1769_));
 sky130_fd_sc_hd__nor2_1 _2103_ (.A(_1735_),
    .B(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__nand2_1 _2104_ (.A(\d2.count[3] ),
    .B(_1733_),
    .Y(_1771_));
 sky130_fd_sc_hd__o21ai_1 _2105_ (.A1(_1727_),
    .A2(\d2.count[5] ),
    .B1(\d2.count[4] ),
    .Y(_1772_));
 sky130_fd_sc_hd__a2bb2o_1 _2106_ (.A1_N(\d2.count[3] ),
    .A2_N(_1733_),
    .B1(_1772_),
    .B2(_1712_),
    .X(_1773_));
 sky130_fd_sc_hd__a21o_1 _2107_ (.A1(_1770_),
    .A2(_1771_),
    .B1(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__a21o_1 _2108_ (.A1(_1721_),
    .A2(\d2.count[4] ),
    .B1(\d2.count[5] ),
    .X(_1775_));
 sky130_fd_sc_hd__nand2_1 _2109_ (.A(_1715_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__buf_6 _2110_ (.A(_1732_),
    .X(_1777_));
 sky130_fd_sc_hd__nand2_1 _2111_ (.A(\d2.count[6] ),
    .B(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__o22ai_1 _2112_ (.A1(\d2.count[7] ),
    .A2(_1723_),
    .B1(_1777_),
    .B2(\d2.count[6] ),
    .Y(_1779_));
 sky130_fd_sc_hd__a31o_1 _2113_ (.A1(_1774_),
    .A2(_1776_),
    .A3(_1778_),
    .B1(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__o2bb2a_1 _2114_ (.A1_N(_1768_),
    .A2_N(_1780_),
    .B1(\d2.count[8] ),
    .B2(_1720_),
    .X(_1781_));
 sky130_fd_sc_hd__nor2_1 _2115_ (.A(\d2.count[9] ),
    .B(_1714_),
    .Y(_1782_));
 sky130_fd_sc_hd__o21bai_4 _2116_ (.A1(_1767_),
    .A2(_1781_),
    .B1_N(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__nand2_1 _2117_ (.A(net111),
    .B(_1783_),
    .Y(\d2.nxt_count[0] ));
 sky130_fd_sc_hd__nand2_1 _2118_ (.A(\d2.count[1] ),
    .B(\d2.count[0] ),
    .Y(_1784_));
 sky130_fd_sc_hd__or2_1 _2119_ (.A(\d2.count[1] ),
    .B(\d2.count[0] ),
    .X(_1785_));
 sky130_fd_sc_hd__and3_1 _2120_ (.A(_1783_),
    .B(_1784_),
    .C(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__clkbuf_1 _2121_ (.A(_1786_),
    .X(\d2.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2122_ (.A(\d2.count[1] ),
    .B(\d2.count[0] ),
    .C(\d2.count[2] ),
    .X(_1787_));
 sky130_fd_sc_hd__inv_2 _2123_ (.A(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__a21o_1 _2124_ (.A1(\d2.count[1] ),
    .A2(\d2.count[0] ),
    .B1(\d2.count[2] ),
    .X(_1789_));
 sky130_fd_sc_hd__and3_1 _2125_ (.A(_1783_),
    .B(_1788_),
    .C(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__clkbuf_1 _2126_ (.A(_1790_),
    .X(\d2.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2127_ (.A(\d2.count[3] ),
    .B(_1787_),
    .X(_1791_));
 sky130_fd_sc_hd__o21ai_1 _2128_ (.A1(net248),
    .A2(_1787_),
    .B1(_1783_),
    .Y(_1792_));
 sky130_fd_sc_hd__nor2_1 _2129_ (.A(_1791_),
    .B(_1792_),
    .Y(\d2.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2130_ (.A(\d2.count[3] ),
    .B(\d2.count[4] ),
    .C(_1787_),
    .X(_1793_));
 sky130_fd_sc_hd__o21ai_1 _2131_ (.A1(net200),
    .A2(_1791_),
    .B1(_1783_),
    .Y(_1794_));
 sky130_fd_sc_hd__nor2_1 _2132_ (.A(_1793_),
    .B(_1794_),
    .Y(\d2.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2133_ (.A(\d2.count[5] ),
    .B(\d2.count[4] ),
    .C(_1791_),
    .X(_1795_));
 sky130_fd_sc_hd__o21ai_1 _2134_ (.A1(net197),
    .A2(_1793_),
    .B1(_1783_),
    .Y(_1796_));
 sky130_fd_sc_hd__nor2_1 _2135_ (.A(_1795_),
    .B(_1796_),
    .Y(\d2.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2136_ (.A(\d2.count[6] ),
    .B(_1795_),
    .X(_1797_));
 sky130_fd_sc_hd__o21ai_1 _2137_ (.A1(\d2.count[6] ),
    .A2(_1795_),
    .B1(_1783_),
    .Y(_1798_));
 sky130_fd_sc_hd__nor2_1 _2138_ (.A(_1797_),
    .B(_1798_),
    .Y(\d2.nxt_count[6] ));
 sky130_fd_sc_hd__and3_1 _2139_ (.A(\d2.count[7] ),
    .B(\d2.count[6] ),
    .C(_1795_),
    .X(_1799_));
 sky130_fd_sc_hd__o21ai_1 _2140_ (.A1(net186),
    .A2(_1797_),
    .B1(_1783_),
    .Y(_1800_));
 sky130_fd_sc_hd__nor2_1 _2141_ (.A(_1799_),
    .B(_1800_),
    .Y(\d2.nxt_count[7] ));
 sky130_fd_sc_hd__o21ai_1 _2142_ (.A1(net98),
    .A2(_1799_),
    .B1(_1783_),
    .Y(_1801_));
 sky130_fd_sc_hd__a21oi_1 _2143_ (.A1(net98),
    .A2(_1799_),
    .B1(_1801_),
    .Y(\d2.nxt_count[8] ));
 sky130_fd_sc_hd__a21o_1 _2144_ (.A1(\d2.count[8] ),
    .A2(_1799_),
    .B1(\d2.count[9] ),
    .X(_1802_));
 sky130_fd_sc_hd__nand3_1 _2145_ (.A(\d2.count[9] ),
    .B(\d2.count[8] ),
    .C(_1799_),
    .Y(_1803_));
 sky130_fd_sc_hd__and3_1 _2146_ (.A(_1783_),
    .B(_1802_),
    .C(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__clkbuf_1 _2147_ (.A(_1804_),
    .X(\d2.nxt_count[9] ));
 sky130_fd_sc_hd__clkbuf_16 _2148_ (.A(_1715_),
    .X(_1805_));
 sky130_fd_sc_hd__a22o_1 _2149_ (.A1(\d3.count[9] ),
    .A2(_1715_),
    .B1(_1718_),
    .B2(\d3.count[8] ),
    .X(_1806_));
 sky130_fd_sc_hd__a22o_1 _2150_ (.A1(\d3.count[7] ),
    .A2(_1723_),
    .B1(_1732_),
    .B2(\d3.count[6] ),
    .X(_1807_));
 sky130_fd_sc_hd__o21ai_1 _2151_ (.A1(_1713_),
    .A2(\d3.count[0] ),
    .B1(\d3.count[1] ),
    .Y(_1808_));
 sky130_fd_sc_hd__a2bb2o_1 _2152_ (.A1_N(\d3.count[2] ),
    .A2_N(_1733_),
    .B1(_1808_),
    .B2(_1721_),
    .X(_1809_));
 sky130_fd_sc_hd__and2_1 _2153_ (.A(_1721_),
    .B(\d3.count[3] ),
    .X(_1810_));
 sky130_fd_sc_hd__a21oi_1 _2154_ (.A1(\d3.count[2] ),
    .A2(_1733_),
    .B1(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__nor2_1 _2155_ (.A(\d3.count[4] ),
    .B(_1714_),
    .Y(_1812_));
 sky130_fd_sc_hd__nor2_1 _2156_ (.A(_1721_),
    .B(\d3.count[3] ),
    .Y(_1813_));
 sky130_fd_sc_hd__a211oi_1 _2157_ (.A1(_1809_),
    .A2(_1811_),
    .B1(_1812_),
    .C1(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__and2_1 _2158_ (.A(\d3.count[4] ),
    .B(_1714_),
    .X(_1815_));
 sky130_fd_sc_hd__o32a_1 _2159_ (.A1(\d3.count[5] ),
    .A2(_1814_),
    .A3(_1815_),
    .B1(_1777_),
    .B2(\d3.count[6] ),
    .X(_1816_));
 sky130_fd_sc_hd__o22ai_1 _2160_ (.A1(\d3.count[8] ),
    .A2(_1718_),
    .B1(_1722_),
    .B2(\d3.count[7] ),
    .Y(_1817_));
 sky130_fd_sc_hd__o21ba_1 _2161_ (.A1(_1807_),
    .A2(_1816_),
    .B1_N(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__o22ai_4 _2162_ (.A1(\d3.count[9] ),
    .A2(_1805_),
    .B1(_1806_),
    .B2(_1818_),
    .Y(_1819_));
 sky130_fd_sc_hd__nand2_1 _2163_ (.A(net73),
    .B(_1819_),
    .Y(\d3.nxt_count[0] ));
 sky130_fd_sc_hd__nand2_1 _2164_ (.A(\d3.count[0] ),
    .B(\d3.count[1] ),
    .Y(_1820_));
 sky130_fd_sc_hd__or2_1 _2165_ (.A(\d3.count[0] ),
    .B(\d3.count[1] ),
    .X(_1821_));
 sky130_fd_sc_hd__and3_1 _2166_ (.A(_1819_),
    .B(_1820_),
    .C(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _2167_ (.A(_1822_),
    .X(\d3.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2168_ (.A(\d3.count[0] ),
    .B(\d3.count[1] ),
    .C(\d3.count[2] ),
    .X(_1823_));
 sky130_fd_sc_hd__inv_2 _2169_ (.A(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__a21o_1 _2170_ (.A1(\d3.count[0] ),
    .A2(\d3.count[1] ),
    .B1(\d3.count[2] ),
    .X(_1825_));
 sky130_fd_sc_hd__and3_1 _2171_ (.A(_1819_),
    .B(_1824_),
    .C(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__clkbuf_1 _2172_ (.A(_1826_),
    .X(\d3.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2173_ (.A(\d3.count[3] ),
    .B(_1823_),
    .X(_1827_));
 sky130_fd_sc_hd__o21ai_1 _2174_ (.A1(net203),
    .A2(_1823_),
    .B1(_1819_),
    .Y(_1828_));
 sky130_fd_sc_hd__nor2_1 _2175_ (.A(_1827_),
    .B(_1828_),
    .Y(\d3.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2176_ (.A(\d3.count[3] ),
    .B(\d3.count[4] ),
    .C(_1823_),
    .X(_1829_));
 sky130_fd_sc_hd__o21ai_1 _2177_ (.A1(net232),
    .A2(_1827_),
    .B1(_1819_),
    .Y(_1830_));
 sky130_fd_sc_hd__nor2_1 _2178_ (.A(_1829_),
    .B(_1830_),
    .Y(\d3.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2179_ (.A(\d3.count[4] ),
    .B(\d3.count[5] ),
    .C(_1827_),
    .X(_1831_));
 sky130_fd_sc_hd__o21ai_1 _2180_ (.A1(net184),
    .A2(_1829_),
    .B1(_1819_),
    .Y(_1832_));
 sky130_fd_sc_hd__nor2_1 _2181_ (.A(_1831_),
    .B(_1832_),
    .Y(\d3.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2182_ (.A(\d3.count[6] ),
    .B(_1831_),
    .X(_1833_));
 sky130_fd_sc_hd__o21ai_1 _2183_ (.A1(net249),
    .A2(_1831_),
    .B1(_1819_),
    .Y(_1834_));
 sky130_fd_sc_hd__nor2_1 _2184_ (.A(_1833_),
    .B(_1834_),
    .Y(\d3.nxt_count[6] ));
 sky130_fd_sc_hd__and3_1 _2185_ (.A(\d3.count[7] ),
    .B(\d3.count[6] ),
    .C(_1831_),
    .X(_1835_));
 sky130_fd_sc_hd__o21ai_1 _2186_ (.A1(net209),
    .A2(_1833_),
    .B1(_1819_),
    .Y(_1836_));
 sky130_fd_sc_hd__nor2_1 _2187_ (.A(_1835_),
    .B(_1836_),
    .Y(\d3.nxt_count[7] ));
 sky130_fd_sc_hd__o21ai_1 _2188_ (.A1(net87),
    .A2(_1835_),
    .B1(_1819_),
    .Y(_1837_));
 sky130_fd_sc_hd__a21oi_1 _2189_ (.A1(net87),
    .A2(_1835_),
    .B1(_1837_),
    .Y(\d3.nxt_count[8] ));
 sky130_fd_sc_hd__a21o_1 _2190_ (.A1(\d3.count[8] ),
    .A2(_1835_),
    .B1(\d3.count[9] ),
    .X(_1838_));
 sky130_fd_sc_hd__nand3_1 _2191_ (.A(\d3.count[9] ),
    .B(\d3.count[8] ),
    .C(_1835_),
    .Y(_1839_));
 sky130_fd_sc_hd__and3_1 _2192_ (.A(_1819_),
    .B(_1838_),
    .C(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__clkbuf_1 _2193_ (.A(_1840_),
    .X(\d3.nxt_count[9] ));
 sky130_fd_sc_hd__nand2_1 _2194_ (.A(\d4.count[6] ),
    .B(_1725_),
    .Y(_1841_));
 sky130_fd_sc_hd__or2_1 _2195_ (.A(\d4.count[6] ),
    .B(_1725_),
    .X(_1842_));
 sky130_fd_sc_hd__o211a_1 _2196_ (.A1(_1713_),
    .A2(\d4.count[0] ),
    .B1(\d4.count[1] ),
    .C1(_1721_),
    .X(_1843_));
 sky130_fd_sc_hd__inv_2 _2197_ (.A(\d4.count[7] ),
    .Y(_1844_));
 sky130_fd_sc_hd__o2111a_1 _2198_ (.A1(_1712_),
    .A2(_1844_),
    .B1(\d4.count[4] ),
    .C1(\d4.count[5] ),
    .D1(\d4.count[3] ),
    .X(_1845_));
 sky130_fd_sc_hd__o221a_1 _2199_ (.A1(\d4.count[2] ),
    .A2(_1724_),
    .B1(_1843_),
    .B2(\d4.count[7] ),
    .C1(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__and3_1 _2200_ (.A(_1841_),
    .B(_1842_),
    .C(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__a22o_1 _2201_ (.A1(_1721_),
    .A2(\d4.count[7] ),
    .B1(\d4.count[6] ),
    .B2(_1725_),
    .X(_1848_));
 sky130_fd_sc_hd__o22a_1 _2202_ (.A1(\d4.count[8] ),
    .A2(_1805_),
    .B1(_1847_),
    .B2(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__a211oi_4 _2203_ (.A1(\d4.count[8] ),
    .A2(_1805_),
    .B1(_1849_),
    .C1(\d4.count[9] ),
    .Y(_1850_));
 sky130_fd_sc_hd__nand2_1 _2204_ (.A(net74),
    .B(_1850_),
    .Y(\d4.nxt_count[0] ));
 sky130_fd_sc_hd__nand2_1 _2205_ (.A(\d4.count[0] ),
    .B(\d4.count[1] ),
    .Y(_1851_));
 sky130_fd_sc_hd__or2_1 _2206_ (.A(\d4.count[0] ),
    .B(\d4.count[1] ),
    .X(_1852_));
 sky130_fd_sc_hd__and3_1 _2207_ (.A(_1850_),
    .B(_1851_),
    .C(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__clkbuf_1 _2208_ (.A(_1853_),
    .X(\d4.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2209_ (.A(\d4.count[0] ),
    .B(\d4.count[1] ),
    .C(\d4.count[2] ),
    .X(_1854_));
 sky130_fd_sc_hd__a21o_1 _2210_ (.A1(\d4.count[0] ),
    .A2(\d4.count[1] ),
    .B1(\d4.count[2] ),
    .X(_1855_));
 sky130_fd_sc_hd__and3b_1 _2211_ (.A_N(_1854_),
    .B(_1855_),
    .C(_1850_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _2212_ (.A(_1856_),
    .X(\d4.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2213_ (.A(\d4.count[3] ),
    .B(_1854_),
    .X(_1857_));
 sky130_fd_sc_hd__or2_1 _2214_ (.A(\d4.count[3] ),
    .B(_1854_),
    .X(_1858_));
 sky130_fd_sc_hd__and3b_1 _2215_ (.A_N(_1857_),
    .B(_1858_),
    .C(_1850_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _2216_ (.A(_1859_),
    .X(\d4.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2217_ (.A(\d4.count[3] ),
    .B(\d4.count[4] ),
    .C(_1854_),
    .X(_1860_));
 sky130_fd_sc_hd__o21ai_1 _2218_ (.A1(net157),
    .A2(_1857_),
    .B1(_1850_),
    .Y(_1861_));
 sky130_fd_sc_hd__nor2_1 _2219_ (.A(_1860_),
    .B(_1861_),
    .Y(\d4.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2220_ (.A(\d4.count[4] ),
    .B(\d4.count[5] ),
    .C(_1857_),
    .X(_1862_));
 sky130_fd_sc_hd__o21ai_1 _2221_ (.A1(net141),
    .A2(_1860_),
    .B1(_1850_),
    .Y(_1863_));
 sky130_fd_sc_hd__nor2_1 _2222_ (.A(_1862_),
    .B(_1863_),
    .Y(\d4.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2223_ (.A(\d4.count[6] ),
    .B(_1862_),
    .X(_1864_));
 sky130_fd_sc_hd__o21ai_1 _2224_ (.A1(net212),
    .A2(_1862_),
    .B1(_1850_),
    .Y(_1865_));
 sky130_fd_sc_hd__nor2_1 _2225_ (.A(_1864_),
    .B(_1865_),
    .Y(\d4.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2226_ (.A(net246),
    .B(_1864_),
    .Y(_1866_));
 sky130_fd_sc_hd__or2_1 _2227_ (.A(\d4.count[7] ),
    .B(_1864_),
    .X(_1867_));
 sky130_fd_sc_hd__and3_1 _2228_ (.A(_1850_),
    .B(_1866_),
    .C(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__clkbuf_1 _2229_ (.A(_1868_),
    .X(\d4.nxt_count[7] ));
 sky130_fd_sc_hd__inv_2 _2230_ (.A(\d4.count[8] ),
    .Y(_1869_));
 sky130_fd_sc_hd__a21boi_1 _2231_ (.A1(_1869_),
    .A2(_1866_),
    .B1_N(_1850_),
    .Y(\d4.nxt_count[8] ));
 sky130_fd_sc_hd__a21oi_1 _2232_ (.A1(_1727_),
    .A2(\d5.count[6] ),
    .B1(\d5.count[7] ),
    .Y(_1870_));
 sky130_fd_sc_hd__nor2_1 _2233_ (.A(_1735_),
    .B(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__buf_6 _2234_ (.A(_1713_),
    .X(_1872_));
 sky130_fd_sc_hd__o211a_1 _2235_ (.A1(_1872_),
    .A2(\d5.count[4] ),
    .B1(\d5.count[5] ),
    .C1(_1735_),
    .X(_1873_));
 sky130_fd_sc_hd__o21a_1 _2236_ (.A1(_1713_),
    .A2(\d5.count[0] ),
    .B1(\d5.count[1] ),
    .X(_1874_));
 sky130_fd_sc_hd__o22a_1 _2237_ (.A1(\d5.count[3] ),
    .A2(_1729_),
    .B1(_1874_),
    .B2(_1712_),
    .X(_1875_));
 sky130_fd_sc_hd__o21ai_1 _2238_ (.A1(\d5.count[2] ),
    .A2(_1733_),
    .B1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__o21ai_1 _2239_ (.A1(\d5.count[2] ),
    .A2(_1729_),
    .B1(\d5.count[3] ),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _2240_ (.A(\d5.count[5] ),
    .B(_1715_),
    .Y(_1878_));
 sky130_fd_sc_hd__or2_1 _2241_ (.A(\d5.count[5] ),
    .B(_1715_),
    .X(_1879_));
 sky130_fd_sc_hd__xor2_1 _2242_ (.A(\d5.count[4] ),
    .B(_1718_),
    .X(_1880_));
 sky130_fd_sc_hd__a21oi_1 _2243_ (.A1(_1878_),
    .A2(_1879_),
    .B1(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hd__inv_2 _2244_ (.A(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__a21oi_1 _2245_ (.A1(_1876_),
    .A2(_1877_),
    .B1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__o21a_1 _2246_ (.A1(_1721_),
    .A2(\d5.count[7] ),
    .B1(\d5.count[6] ),
    .X(_1884_));
 sky130_fd_sc_hd__nor2_1 _2247_ (.A(_1725_),
    .B(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__o21ba_1 _2248_ (.A1(_1873_),
    .A2(_1883_),
    .B1_N(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__o22a_1 _2249_ (.A1(\d5.count[8] ),
    .A2(_1805_),
    .B1(_1871_),
    .B2(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__a211oi_4 _2250_ (.A1(\d5.count[8] ),
    .A2(_1805_),
    .B1(_1887_),
    .C1(net228),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_1 _2251_ (.A(net82),
    .B(_1888_),
    .Y(\d5.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2252_ (.A(\d5.count[0] ),
    .B(\d5.count[1] ),
    .X(_1889_));
 sky130_fd_sc_hd__nand2_1 _2253_ (.A(\d5.count[0] ),
    .B(\d5.count[1] ),
    .Y(_1890_));
 sky130_fd_sc_hd__and3_1 _2254_ (.A(_1888_),
    .B(_1889_),
    .C(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__clkbuf_1 _2255_ (.A(_1891_),
    .X(\d5.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2256_ (.A(\d5.count[0] ),
    .B(\d5.count[1] ),
    .C(\d5.count[2] ),
    .X(_1892_));
 sky130_fd_sc_hd__a21o_1 _2257_ (.A1(\d5.count[0] ),
    .A2(\d5.count[1] ),
    .B1(\d5.count[2] ),
    .X(_1893_));
 sky130_fd_sc_hd__and3b_1 _2258_ (.A_N(_1892_),
    .B(_1893_),
    .C(_1888_),
    .X(_1894_));
 sky130_fd_sc_hd__clkbuf_1 _2259_ (.A(_1894_),
    .X(\d5.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2260_ (.A(\d5.count[3] ),
    .B(_1892_),
    .X(_1895_));
 sky130_fd_sc_hd__or2_1 _2261_ (.A(\d5.count[3] ),
    .B(_1892_),
    .X(_1896_));
 sky130_fd_sc_hd__and3b_1 _2262_ (.A_N(_1895_),
    .B(_1896_),
    .C(_1888_),
    .X(_1897_));
 sky130_fd_sc_hd__clkbuf_1 _2263_ (.A(_1897_),
    .X(\d5.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2264_ (.A(\d5.count[3] ),
    .B(\d5.count[4] ),
    .C(_1892_),
    .X(_1898_));
 sky130_fd_sc_hd__o21ai_1 _2265_ (.A1(\d5.count[4] ),
    .A2(_1895_),
    .B1(_1888_),
    .Y(_1899_));
 sky130_fd_sc_hd__nor2_1 _2266_ (.A(_1898_),
    .B(_1899_),
    .Y(\d5.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2267_ (.A(\d5.count[5] ),
    .B(\d5.count[4] ),
    .C(_1895_),
    .X(_1900_));
 sky130_fd_sc_hd__o21ai_1 _2268_ (.A1(net194),
    .A2(_1898_),
    .B1(_1888_),
    .Y(_1901_));
 sky130_fd_sc_hd__nor2_1 _2269_ (.A(_1900_),
    .B(net195),
    .Y(\d5.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2270_ (.A(\d5.count[6] ),
    .B(_1900_),
    .X(_1902_));
 sky130_fd_sc_hd__o21ai_1 _2271_ (.A1(net162),
    .A2(_1900_),
    .B1(_1888_),
    .Y(_1903_));
 sky130_fd_sc_hd__nor2_1 _2272_ (.A(_1902_),
    .B(net163),
    .Y(\d5.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2273_ (.A(\d5.count[7] ),
    .B(_1902_),
    .Y(_1904_));
 sky130_fd_sc_hd__or2_1 _2274_ (.A(\d5.count[7] ),
    .B(_1902_),
    .X(_1905_));
 sky130_fd_sc_hd__and3_1 _2275_ (.A(_1888_),
    .B(_1904_),
    .C(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_1 _2276_ (.A(_1906_),
    .X(\d5.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2277_ (.A(\d5.count[8] ),
    .B(_1904_),
    .Y(_1907_));
 sky130_fd_sc_hd__and2_1 _2278_ (.A(_1888_),
    .B(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__clkbuf_1 _2279_ (.A(_1908_),
    .X(\d5.nxt_count[8] ));
 sky130_fd_sc_hd__a21o_1 _2280_ (.A1(_1727_),
    .A2(\d6.count[6] ),
    .B1(\d6.count[7] ),
    .X(_1909_));
 sky130_fd_sc_hd__nand2_1 _2281_ (.A(_1721_),
    .B(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hd__o21ai_1 _2282_ (.A1(_1721_),
    .A2(\d6.count[7] ),
    .B1(\d6.count[6] ),
    .Y(_1911_));
 sky130_fd_sc_hd__a21o_1 _2283_ (.A1(_1872_),
    .A2(\d6.count[5] ),
    .B1(\d6.count[4] ),
    .X(_1912_));
 sky130_fd_sc_hd__nand2_1 _2284_ (.A(_1735_),
    .B(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__a21oi_1 _2285_ (.A1(\d6.count[5] ),
    .A2(_1910_),
    .B1(_1724_),
    .Y(_1914_));
 sky130_fd_sc_hd__a211o_1 _2286_ (.A1(_1777_),
    .A2(_1911_),
    .B1(_1913_),
    .C1(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__o21a_1 _2287_ (.A1(_1872_),
    .A2(\d6.count[3] ),
    .B1(\d6.count[4] ),
    .X(_1916_));
 sky130_fd_sc_hd__a21oi_1 _2288_ (.A1(_1777_),
    .A2(_1911_),
    .B1(_1914_),
    .Y(_1917_));
 sky130_fd_sc_hd__o211ai_1 _2289_ (.A1(_1735_),
    .A2(_1916_),
    .B1(_1913_),
    .C1(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__nor2_1 _2290_ (.A(\d6.count[8] ),
    .B(_1715_),
    .Y(_1919_));
 sky130_fd_sc_hd__a31o_1 _2291_ (.A1(_1910_),
    .A2(_1915_),
    .A3(_1918_),
    .B1(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__a21oi_1 _2292_ (.A1(\d6.count[8] ),
    .A2(_1715_),
    .B1(\d6.count[9] ),
    .Y(_1921_));
 sky130_fd_sc_hd__and2_2 _2293_ (.A(_1920_),
    .B(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__nand2_1 _2294_ (.A(net70),
    .B(_1922_),
    .Y(\d6.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2295_ (.A(\d6.count[1] ),
    .B(\d6.count[0] ),
    .X(_1923_));
 sky130_fd_sc_hd__nand2_1 _2296_ (.A(\d6.count[1] ),
    .B(\d6.count[0] ),
    .Y(_1924_));
 sky130_fd_sc_hd__and3_1 _2297_ (.A(_1922_),
    .B(_1923_),
    .C(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__clkbuf_1 _2298_ (.A(_1925_),
    .X(\d6.nxt_count[1] ));
 sky130_fd_sc_hd__nand3_1 _2299_ (.A(\d6.count[1] ),
    .B(\d6.count[0] ),
    .C(\d6.count[2] ),
    .Y(_1926_));
 sky130_fd_sc_hd__a21o_1 _2300_ (.A1(\d6.count[1] ),
    .A2(\d6.count[0] ),
    .B1(\d6.count[2] ),
    .X(_1927_));
 sky130_fd_sc_hd__and3_1 _2301_ (.A(_1922_),
    .B(_1926_),
    .C(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__clkbuf_1 _2302_ (.A(_1928_),
    .X(\d6.nxt_count[2] ));
 sky130_fd_sc_hd__and4_1 _2303_ (.A(\d6.count[1] ),
    .B(\d6.count[0] ),
    .C(\d6.count[3] ),
    .D(\d6.count[2] ),
    .X(_1929_));
 sky130_fd_sc_hd__a31o_1 _2304_ (.A1(\d6.count[1] ),
    .A2(\d6.count[0] ),
    .A3(\d6.count[2] ),
    .B1(\d6.count[3] ),
    .X(_1930_));
 sky130_fd_sc_hd__and3b_1 _2305_ (.A_N(_1929_),
    .B(_1930_),
    .C(_1922_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _2306_ (.A(_1931_),
    .X(\d6.nxt_count[3] ));
 sky130_fd_sc_hd__o21ai_1 _2307_ (.A1(\d6.count[4] ),
    .A2(_1929_),
    .B1(_1922_),
    .Y(_1932_));
 sky130_fd_sc_hd__a21oi_1 _2308_ (.A1(net138),
    .A2(_1929_),
    .B1(_1932_),
    .Y(\d6.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2309_ (.A(\d6.count[4] ),
    .B(\d6.count[5] ),
    .C(_1929_),
    .X(_1933_));
 sky130_fd_sc_hd__a21o_1 _2310_ (.A1(\d6.count[4] ),
    .A2(_1929_),
    .B1(\d6.count[5] ),
    .X(_1934_));
 sky130_fd_sc_hd__and3b_1 _2311_ (.A_N(_1933_),
    .B(_1934_),
    .C(_1922_),
    .X(_1935_));
 sky130_fd_sc_hd__clkbuf_1 _2312_ (.A(_1935_),
    .X(\d6.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2313_ (.A(\d6.count[6] ),
    .B(_1933_),
    .X(_1936_));
 sky130_fd_sc_hd__o21ai_1 _2314_ (.A1(net148),
    .A2(_1933_),
    .B1(_1922_),
    .Y(_1937_));
 sky130_fd_sc_hd__nor2_1 _2315_ (.A(_1936_),
    .B(_1937_),
    .Y(\d6.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2316_ (.A(\d6.count[7] ),
    .B(_1936_),
    .Y(_1938_));
 sky130_fd_sc_hd__or2_1 _2317_ (.A(\d6.count[7] ),
    .B(_1936_),
    .X(_1939_));
 sky130_fd_sc_hd__and3_1 _2318_ (.A(_1922_),
    .B(_1938_),
    .C(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__clkbuf_1 _2319_ (.A(_1940_),
    .X(\d6.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2320_ (.A(\d6.count[8] ),
    .B(_1938_),
    .Y(_1941_));
 sky130_fd_sc_hd__and3_1 _2321_ (.A(_1920_),
    .B(_1921_),
    .C(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__clkbuf_1 _2322_ (.A(_1942_),
    .X(\d6.nxt_count[8] ));
 sky130_fd_sc_hd__nand2_1 _2323_ (.A(_1872_),
    .B(\d7.count[4] ),
    .Y(_1943_));
 sky130_fd_sc_hd__nand2_1 _2324_ (.A(_1720_),
    .B(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__inv_2 _2325_ (.A(_1718_),
    .Y(_1945_));
 sky130_fd_sc_hd__a21boi_1 _2326_ (.A1(_1735_),
    .A2(\d7.count[5] ),
    .B1_N(\d7.count[4] ),
    .Y(_1946_));
 sky130_fd_sc_hd__o221a_1 _2327_ (.A1(\d7.count[5] ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(_1872_),
    .C1(_1943_),
    .X(_1947_));
 sky130_fd_sc_hd__o21ai_1 _2328_ (.A1(_1727_),
    .A2(\d7.count[2] ),
    .B1(\d7.count[3] ),
    .Y(_1948_));
 sky130_fd_sc_hd__o22a_1 _2329_ (.A1(\d7.count[1] ),
    .A2(_1723_),
    .B1(_1777_),
    .B2(\d7.count[0] ),
    .X(_1949_));
 sky130_fd_sc_hd__and2_1 _2330_ (.A(_1727_),
    .B(\d7.count[2] ),
    .X(_1950_));
 sky130_fd_sc_hd__o221ai_1 _2331_ (.A1(\d7.count[1] ),
    .A2(_1949_),
    .B1(_1950_),
    .B2(\d7.count[3] ),
    .C1(_1948_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand2_1 _2332_ (.A(_1948_),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__a22o_1 _2333_ (.A1(\d7.count[5] ),
    .A2(_1944_),
    .B1(_1947_),
    .B2(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__o21a_1 _2334_ (.A1(\d7.count[6] ),
    .A2(_1733_),
    .B1(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__and2_1 _2335_ (.A(_1721_),
    .B(\d7.count[7] ),
    .X(_1955_));
 sky130_fd_sc_hd__a211oi_1 _2336_ (.A1(\d7.count[6] ),
    .A2(_1733_),
    .B1(_1954_),
    .C1(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__o22ai_2 _2337_ (.A1(_1721_),
    .A2(\d7.count[7] ),
    .B1(\d7.count[8] ),
    .B2(_1805_),
    .Y(_1957_));
 sky130_fd_sc_hd__a21oi_1 _2338_ (.A1(\d7.count[8] ),
    .A2(_1805_),
    .B1(\d7.count[9] ),
    .Y(_1958_));
 sky130_fd_sc_hd__o21a_2 _2339_ (.A1(_1956_),
    .A2(_1957_),
    .B1(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__nand2_1 _2340_ (.A(net85),
    .B(_1959_),
    .Y(\d7.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2341_ (.A(\d7.count[0] ),
    .B(\d7.count[1] ),
    .X(_1960_));
 sky130_fd_sc_hd__nand2_1 _2342_ (.A(\d7.count[0] ),
    .B(\d7.count[1] ),
    .Y(_1961_));
 sky130_fd_sc_hd__and3_1 _2343_ (.A(_1959_),
    .B(_1960_),
    .C(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__clkbuf_1 _2344_ (.A(_1962_),
    .X(\d7.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2345_ (.A(\d7.count[0] ),
    .B(\d7.count[1] ),
    .C(\d7.count[2] ),
    .X(_1963_));
 sky130_fd_sc_hd__a21o_1 _2346_ (.A1(\d7.count[0] ),
    .A2(\d7.count[1] ),
    .B1(\d7.count[2] ),
    .X(_1964_));
 sky130_fd_sc_hd__and3b_1 _2347_ (.A_N(_1963_),
    .B(_1964_),
    .C(_1959_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_1 _2348_ (.A(_1965_),
    .X(\d7.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2349_ (.A(\d7.count[3] ),
    .B(_1963_),
    .X(_1966_));
 sky130_fd_sc_hd__or2_1 _2350_ (.A(\d7.count[3] ),
    .B(_1963_),
    .X(_1967_));
 sky130_fd_sc_hd__and3b_1 _2351_ (.A_N(_1966_),
    .B(_1967_),
    .C(_1959_),
    .X(_1968_));
 sky130_fd_sc_hd__clkbuf_1 _2352_ (.A(_1968_),
    .X(\d7.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2353_ (.A(\d7.count[3] ),
    .B(\d7.count[4] ),
    .C(_1963_),
    .X(_1969_));
 sky130_fd_sc_hd__o21ai_1 _2354_ (.A1(net181),
    .A2(_1966_),
    .B1(_1959_),
    .Y(_1970_));
 sky130_fd_sc_hd__nor2_1 _2355_ (.A(_1969_),
    .B(_1970_),
    .Y(\d7.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2356_ (.A(\d7.count[5] ),
    .B(\d7.count[4] ),
    .C(_1966_),
    .X(_1971_));
 sky130_fd_sc_hd__o21ai_1 _2357_ (.A1(net237),
    .A2(_1969_),
    .B1(_1959_),
    .Y(_1972_));
 sky130_fd_sc_hd__nor2_1 _2358_ (.A(_1971_),
    .B(_1972_),
    .Y(\d7.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2359_ (.A(\d7.count[6] ),
    .B(_1971_),
    .X(_1973_));
 sky130_fd_sc_hd__o21ai_1 _2360_ (.A1(\d7.count[6] ),
    .A2(_1971_),
    .B1(_1959_),
    .Y(_1974_));
 sky130_fd_sc_hd__nor2_1 _2361_ (.A(_1973_),
    .B(_1974_),
    .Y(\d7.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2362_ (.A(\d7.count[7] ),
    .B(_1973_),
    .Y(_1975_));
 sky130_fd_sc_hd__or2_1 _2363_ (.A(\d7.count[7] ),
    .B(_1973_),
    .X(_1976_));
 sky130_fd_sc_hd__and3_1 _2364_ (.A(_1959_),
    .B(_1975_),
    .C(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__clkbuf_1 _2365_ (.A(_1977_),
    .X(\d7.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2366_ (.A(\d7.count[8] ),
    .B(_1975_),
    .Y(_1978_));
 sky130_fd_sc_hd__and2_1 _2367_ (.A(_1959_),
    .B(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__clkbuf_1 _2368_ (.A(_1979_),
    .X(\d7.nxt_count[8] ));
 sky130_fd_sc_hd__nor2_1 _2369_ (.A(\d8.count[4] ),
    .B(_1726_),
    .Y(_1980_));
 sky130_fd_sc_hd__a211o_1 _2370_ (.A1(_1727_),
    .A2(\d8.count[1] ),
    .B1(\d8.count[2] ),
    .C1(_1735_),
    .X(_1981_));
 sky130_fd_sc_hd__a21oi_1 _2371_ (.A1(_1720_),
    .A2(_1981_),
    .B1(\d8.count[3] ),
    .Y(_1982_));
 sky130_fd_sc_hd__a22oi_1 _2372_ (.A1(_1735_),
    .A2(\d8.count[5] ),
    .B1(\d8.count[4] ),
    .B2(_1726_),
    .Y(_1983_));
 sky130_fd_sc_hd__o21ai_1 _2373_ (.A1(_1980_),
    .A2(_1982_),
    .B1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__o221a_1 _2374_ (.A1(_1735_),
    .A2(\d8.count[5] ),
    .B1(_1733_),
    .B2(\d8.count[6] ),
    .C1(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__nand2_1 _2375_ (.A(_1721_),
    .B(\d8.count[7] ),
    .Y(_1986_));
 sky130_fd_sc_hd__a21bo_1 _2376_ (.A1(\d8.count[6] ),
    .A2(_1733_),
    .B1_N(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__or2_1 _2377_ (.A(_1721_),
    .B(\d8.count[7] ),
    .X(_1988_));
 sky130_fd_sc_hd__o221a_1 _2378_ (.A1(\d8.count[8] ),
    .A2(_1805_),
    .B1(_1985_),
    .B2(_1987_),
    .C1(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__a211oi_4 _2379_ (.A1(\d8.count[8] ),
    .A2(_1805_),
    .B1(_1989_),
    .C1(\d8.count[9] ),
    .Y(_1990_));
 sky130_fd_sc_hd__nand2_1 _2380_ (.A(net68),
    .B(_1990_),
    .Y(\d8.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2381_ (.A(\d8.count[1] ),
    .B(\d8.count[0] ),
    .X(_1991_));
 sky130_fd_sc_hd__nand2_1 _2382_ (.A(\d8.count[1] ),
    .B(\d8.count[0] ),
    .Y(_1992_));
 sky130_fd_sc_hd__and3_1 _2383_ (.A(_1990_),
    .B(_1991_),
    .C(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__clkbuf_1 _2384_ (.A(_1993_),
    .X(\d8.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2385_ (.A(\d8.count[1] ),
    .B(\d8.count[0] ),
    .C(\d8.count[2] ),
    .X(_1994_));
 sky130_fd_sc_hd__a21o_1 _2386_ (.A1(\d8.count[1] ),
    .A2(\d8.count[0] ),
    .B1(\d8.count[2] ),
    .X(_1995_));
 sky130_fd_sc_hd__and3b_1 _2387_ (.A_N(_1994_),
    .B(_1995_),
    .C(_1990_),
    .X(_1996_));
 sky130_fd_sc_hd__clkbuf_1 _2388_ (.A(_1996_),
    .X(\d8.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2389_ (.A(\d8.count[3] ),
    .B(_1994_),
    .X(_1997_));
 sky130_fd_sc_hd__or2_1 _2390_ (.A(\d8.count[3] ),
    .B(_1994_),
    .X(_1998_));
 sky130_fd_sc_hd__and3b_1 _2391_ (.A_N(_1997_),
    .B(_1998_),
    .C(_1990_),
    .X(_1999_));
 sky130_fd_sc_hd__clkbuf_1 _2392_ (.A(_1999_),
    .X(\d8.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2393_ (.A(\d8.count[3] ),
    .B(\d8.count[4] ),
    .C(_1994_),
    .X(_2000_));
 sky130_fd_sc_hd__o21ai_1 _2394_ (.A1(net236),
    .A2(_1997_),
    .B1(_1990_),
    .Y(_2001_));
 sky130_fd_sc_hd__nor2_1 _2395_ (.A(_2000_),
    .B(_2001_),
    .Y(\d8.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2396_ (.A(\d8.count[5] ),
    .B(\d8.count[4] ),
    .C(_1997_),
    .X(_2002_));
 sky130_fd_sc_hd__o21ai_1 _2397_ (.A1(\d8.count[5] ),
    .A2(_2000_),
    .B1(_1990_),
    .Y(_2003_));
 sky130_fd_sc_hd__nor2_1 _2398_ (.A(_2002_),
    .B(_2003_),
    .Y(\d8.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2399_ (.A(\d8.count[6] ),
    .B(_2002_),
    .X(_2004_));
 sky130_fd_sc_hd__o21ai_1 _2400_ (.A1(net227),
    .A2(_2002_),
    .B1(_1990_),
    .Y(_2005_));
 sky130_fd_sc_hd__nor2_1 _2401_ (.A(_2004_),
    .B(_2005_),
    .Y(\d8.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2402_ (.A(\d8.count[7] ),
    .B(_2004_),
    .Y(_2006_));
 sky130_fd_sc_hd__or2_1 _2403_ (.A(\d8.count[7] ),
    .B(_2004_),
    .X(_2007_));
 sky130_fd_sc_hd__and3_1 _2404_ (.A(_1990_),
    .B(_2006_),
    .C(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__clkbuf_1 _2405_ (.A(_2008_),
    .X(\d8.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2406_ (.A(\d8.count[8] ),
    .B(_2006_),
    .Y(_2009_));
 sky130_fd_sc_hd__and2_1 _2407_ (.A(_1990_),
    .B(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__clkbuf_1 _2408_ (.A(_2010_),
    .X(\d8.nxt_count[8] ));
 sky130_fd_sc_hd__or2_1 _2409_ (.A(_1727_),
    .B(\d9.count[6] ),
    .X(_2011_));
 sky130_fd_sc_hd__xnor2_1 _2410_ (.A(\d9.count[5] ),
    .B(_1723_),
    .Y(_2012_));
 sky130_fd_sc_hd__nand2_1 _2411_ (.A(\d9.count[4] ),
    .B(_1725_),
    .Y(_2013_));
 sky130_fd_sc_hd__or2_1 _2412_ (.A(\d9.count[4] ),
    .B(_1725_),
    .X(_2014_));
 sky130_fd_sc_hd__and3_1 _2413_ (.A(_2012_),
    .B(_2013_),
    .C(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__o21ai_1 _2414_ (.A1(_1713_),
    .A2(\d9.count[0] ),
    .B1(\d9.count[1] ),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _2415_ (.A(_1721_),
    .B(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hd__o2111a_1 _2416_ (.A1(\d9.count[2] ),
    .A2(_1724_),
    .B1(_2015_),
    .C1(_2017_),
    .D1(\d9.count[3] ),
    .X(_2018_));
 sky130_fd_sc_hd__o211a_1 _2417_ (.A1(_1872_),
    .A2(\d9.count[4] ),
    .B1(\d9.count[5] ),
    .C1(_1721_),
    .X(_2019_));
 sky130_fd_sc_hd__a211o_1 _2418_ (.A1(_1727_),
    .A2(\d9.count[6] ),
    .B1(_2018_),
    .C1(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__a22o_1 _2419_ (.A1(\d9.count[7] ),
    .A2(_1720_),
    .B1(_2011_),
    .B2(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__o221a_1 _2420_ (.A1(\d9.count[8] ),
    .A2(_1805_),
    .B1(_1720_),
    .B2(\d9.count[7] ),
    .C1(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__a211oi_4 _2421_ (.A1(\d9.count[8] ),
    .A2(_1805_),
    .B1(_2022_),
    .C1(\d9.count[9] ),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2_1 _2422_ (.A(net76),
    .B(_2023_),
    .Y(\d9.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2423_ (.A(\d9.count[0] ),
    .B(\d9.count[1] ),
    .X(_2024_));
 sky130_fd_sc_hd__nand2_1 _2424_ (.A(\d9.count[0] ),
    .B(\d9.count[1] ),
    .Y(_2025_));
 sky130_fd_sc_hd__and3_1 _2425_ (.A(_2023_),
    .B(_2024_),
    .C(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__clkbuf_1 _2426_ (.A(_2026_),
    .X(\d9.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2427_ (.A(\d9.count[0] ),
    .B(\d9.count[1] ),
    .C(\d9.count[2] ),
    .X(_2027_));
 sky130_fd_sc_hd__a21o_1 _2428_ (.A1(\d9.count[0] ),
    .A2(\d9.count[1] ),
    .B1(\d9.count[2] ),
    .X(_2028_));
 sky130_fd_sc_hd__and3b_1 _2429_ (.A_N(_2027_),
    .B(_2028_),
    .C(_2023_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _2430_ (.A(_0146_),
    .X(\d9.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2431_ (.A(\d9.count[3] ),
    .B(_2027_),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _2432_ (.A(\d9.count[3] ),
    .B(_2027_),
    .X(_0148_));
 sky130_fd_sc_hd__and3b_1 _2433_ (.A_N(_0147_),
    .B(_0148_),
    .C(_2023_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _2434_ (.A(_0149_),
    .X(\d9.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2435_ (.A(\d9.count[3] ),
    .B(\d9.count[4] ),
    .C(_2027_),
    .X(_0150_));
 sky130_fd_sc_hd__o21ai_1 _2436_ (.A1(\d9.count[4] ),
    .A2(_0147_),
    .B1(_2023_),
    .Y(_0151_));
 sky130_fd_sc_hd__nor2_1 _2437_ (.A(_0150_),
    .B(_0151_),
    .Y(\d9.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2438_ (.A(\d9.count[5] ),
    .B(\d9.count[4] ),
    .C(_0147_),
    .X(_0152_));
 sky130_fd_sc_hd__o21ai_1 _2439_ (.A1(net205),
    .A2(_0150_),
    .B1(_2023_),
    .Y(_0153_));
 sky130_fd_sc_hd__nor2_1 _2440_ (.A(_0152_),
    .B(_0153_),
    .Y(\d9.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2441_ (.A(\d9.count[6] ),
    .B(_0152_),
    .X(_0154_));
 sky130_fd_sc_hd__o21ai_1 _2442_ (.A1(net240),
    .A2(_0152_),
    .B1(_2023_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor2_1 _2443_ (.A(_0154_),
    .B(_0155_),
    .Y(\d9.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2444_ (.A(\d9.count[7] ),
    .B(_0154_),
    .Y(_0156_));
 sky130_fd_sc_hd__or2_1 _2445_ (.A(\d9.count[7] ),
    .B(_0154_),
    .X(_0157_));
 sky130_fd_sc_hd__and3_1 _2446_ (.A(_2023_),
    .B(_0156_),
    .C(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _2447_ (.A(_0158_),
    .X(\d9.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2448_ (.A(\d9.count[8] ),
    .B(_0156_),
    .Y(_0159_));
 sky130_fd_sc_hd__and2_1 _2449_ (.A(_2023_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _2450_ (.A(_0160_),
    .X(\d9.nxt_count[8] ));
 sky130_fd_sc_hd__o22a_1 _2451_ (.A1(\d10.count[8] ),
    .A2(_1715_),
    .B1(_1718_),
    .B2(\d10.count[7] ),
    .X(_0161_));
 sky130_fd_sc_hd__nor2_1 _2452_ (.A(_1727_),
    .B(\d10.count[6] ),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _2453_ (.A(\d10.count[6] ),
    .Y(_0163_));
 sky130_fd_sc_hd__nand2_1 _2454_ (.A(\d10.count[4] ),
    .B(_1733_),
    .Y(_0164_));
 sky130_fd_sc_hd__a21bo_1 _2455_ (.A1(_1723_),
    .A2(_0164_),
    .B1_N(\d10.count[5] ),
    .X(_0165_));
 sky130_fd_sc_hd__o21a_1 _2456_ (.A1(_1872_),
    .A2(\d10.count[2] ),
    .B1(\d10.count[3] ),
    .X(_0166_));
 sky130_fd_sc_hd__o22a_1 _2457_ (.A1(\d10.count[4] ),
    .A2(_1733_),
    .B1(_0166_),
    .B2(_1735_),
    .X(_0167_));
 sky130_fd_sc_hd__o211ai_1 _2458_ (.A1(\d10.count[5] ),
    .A2(_1729_),
    .B1(_0164_),
    .C1(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__o211a_1 _2459_ (.A1(_1872_),
    .A2(_0163_),
    .B1(_0165_),
    .C1(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__a2bb2o_1 _2460_ (.A1_N(_0162_),
    .A2_N(_0169_),
    .B1(\d10.count[7] ),
    .B2(_1720_),
    .X(_0170_));
 sky130_fd_sc_hd__a21o_1 _2461_ (.A1(\d10.count[8] ),
    .A2(_1715_),
    .B1(\d10.count[9] ),
    .X(_0171_));
 sky130_fd_sc_hd__a21oi_4 _2462_ (.A1(_0161_),
    .A2(_0170_),
    .B1(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _2463_ (.A(net86),
    .B(_0172_),
    .Y(\d10.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2464_ (.A(\d10.count[1] ),
    .B(\d10.count[0] ),
    .X(_0173_));
 sky130_fd_sc_hd__nand2_1 _2465_ (.A(\d10.count[1] ),
    .B(\d10.count[0] ),
    .Y(_0174_));
 sky130_fd_sc_hd__and3_1 _2466_ (.A(_0172_),
    .B(_0173_),
    .C(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_1 _2467_ (.A(_0175_),
    .X(\d10.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2468_ (.A(\d10.count[1] ),
    .B(\d10.count[0] ),
    .C(\d10.count[2] ),
    .X(_0176_));
 sky130_fd_sc_hd__a21o_1 _2469_ (.A1(\d10.count[1] ),
    .A2(\d10.count[0] ),
    .B1(\d10.count[2] ),
    .X(_0177_));
 sky130_fd_sc_hd__and3b_1 _2470_ (.A_N(_0176_),
    .B(_0177_),
    .C(_0172_),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_1 _2471_ (.A(_0178_),
    .X(\d10.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2472_ (.A(\d10.count[3] ),
    .B(_0176_),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _2473_ (.A(\d10.count[3] ),
    .B(_0176_),
    .X(_0180_));
 sky130_fd_sc_hd__and3b_1 _2474_ (.A_N(_0179_),
    .B(_0180_),
    .C(_0172_),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _2475_ (.A(_0181_),
    .X(\d10.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2476_ (.A(\d10.count[3] ),
    .B(\d10.count[4] ),
    .C(_0176_),
    .X(_0182_));
 sky130_fd_sc_hd__o21ai_1 _2477_ (.A1(net223),
    .A2(_0179_),
    .B1(_0172_),
    .Y(_0183_));
 sky130_fd_sc_hd__nor2_1 _2478_ (.A(_0182_),
    .B(_0183_),
    .Y(\d10.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2479_ (.A(\d10.count[5] ),
    .B(\d10.count[4] ),
    .C(_0179_),
    .X(_0184_));
 sky130_fd_sc_hd__o21ai_1 _2480_ (.A1(net214),
    .A2(_0182_),
    .B1(_0172_),
    .Y(_0185_));
 sky130_fd_sc_hd__nor2_1 _2481_ (.A(_0184_),
    .B(_0185_),
    .Y(\d10.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2482_ (.A(\d10.count[6] ),
    .B(_0184_),
    .X(_0186_));
 sky130_fd_sc_hd__o21ai_1 _2483_ (.A1(net193),
    .A2(_0184_),
    .B1(_0172_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _2484_ (.A(_0186_),
    .B(_0187_),
    .Y(\d10.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2485_ (.A(\d10.count[7] ),
    .B(_0186_),
    .Y(_0188_));
 sky130_fd_sc_hd__or2_1 _2486_ (.A(\d10.count[7] ),
    .B(_0186_),
    .X(_0189_));
 sky130_fd_sc_hd__and3_1 _2487_ (.A(_0172_),
    .B(_0188_),
    .C(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _2488_ (.A(_0190_),
    .X(\d10.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2489_ (.A(\d10.count[8] ),
    .B(_0188_),
    .Y(_0191_));
 sky130_fd_sc_hd__and2_1 _2490_ (.A(_0172_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _2491_ (.A(_0192_),
    .X(\d10.nxt_count[8] ));
 sky130_fd_sc_hd__o22a_1 _2492_ (.A1(_1727_),
    .A2(\d11.count[6] ),
    .B1(_1718_),
    .B2(\d11.count[7] ),
    .X(_0193_));
 sky130_fd_sc_hd__a21o_1 _2493_ (.A1(_1713_),
    .A2(\d11.count[4] ),
    .B1(\d11.count[5] ),
    .X(_0194_));
 sky130_fd_sc_hd__inv_2 _2494_ (.A(\d11.count[2] ),
    .Y(_0195_));
 sky130_fd_sc_hd__xor2_1 _2495_ (.A(_1872_),
    .B(\d11.count[3] ),
    .X(_0196_));
 sky130_fd_sc_hd__o22a_1 _2496_ (.A1(\d11.count[2] ),
    .A2(_1723_),
    .B1(_1777_),
    .B2(\d11.count[1] ),
    .X(_0197_));
 sky130_fd_sc_hd__o211a_1 _2497_ (.A1(_0195_),
    .A2(_1729_),
    .B1(_0196_),
    .C1(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__o21a_1 _2498_ (.A1(_1872_),
    .A2(\d11.count[3] ),
    .B1(\d11.count[2] ),
    .X(_0199_));
 sky130_fd_sc_hd__a211o_1 _2499_ (.A1(_1872_),
    .A2(\d11.count[3] ),
    .B1(_0198_),
    .C1(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _2500_ (.A(_1727_),
    .B(\d11.count[6] ),
    .X(_0201_));
 sky130_fd_sc_hd__o21a_1 _2501_ (.A1(_1872_),
    .A2(\d11.count[4] ),
    .B1(\d11.count[5] ),
    .X(_0202_));
 sky130_fd_sc_hd__a211o_1 _2502_ (.A1(_0194_),
    .A2(_0200_),
    .B1(_0201_),
    .C1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_1 _2503_ (.A1(\d11.count[7] ),
    .A2(_1720_),
    .B1(_0193_),
    .B2(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__o21ai_1 _2504_ (.A1(\d11.count[8] ),
    .A2(_1805_),
    .B1(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__a21oi_1 _2505_ (.A1(\d11.count[8] ),
    .A2(_1715_),
    .B1(\d11.count[9] ),
    .Y(_0206_));
 sky130_fd_sc_hd__and2_1 _2506_ (.A(_0205_),
    .B(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_2 _2507_ (.A(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _2508_ (.A(net65),
    .B(_0208_),
    .Y(\d11.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2509_ (.A(\d11.count[1] ),
    .B(\d11.count[0] ),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _2510_ (.A(\d11.count[1] ),
    .B(\d11.count[0] ),
    .Y(_0210_));
 sky130_fd_sc_hd__and3_1 _2511_ (.A(_0208_),
    .B(_0209_),
    .C(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _2512_ (.A(_0211_),
    .X(\d11.nxt_count[1] ));
 sky130_fd_sc_hd__nor2_1 _2513_ (.A(_0195_),
    .B(_0210_),
    .Y(_0212_));
 sky130_fd_sc_hd__nand2_1 _2514_ (.A(_0195_),
    .B(_0210_),
    .Y(_0213_));
 sky130_fd_sc_hd__and3b_1 _2515_ (.A_N(_0212_),
    .B(_0213_),
    .C(_0208_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _2516_ (.A(_0214_),
    .X(\d11.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2517_ (.A(\d11.count[3] ),
    .B(_0212_),
    .X(_0215_));
 sky130_fd_sc_hd__or2_1 _2518_ (.A(\d11.count[3] ),
    .B(_0212_),
    .X(_0216_));
 sky130_fd_sc_hd__and3b_1 _2519_ (.A_N(_0215_),
    .B(_0216_),
    .C(_0208_),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_1 _2520_ (.A(_0217_),
    .X(\d11.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2521_ (.A(\d11.count[3] ),
    .B(\d11.count[4] ),
    .C(_0212_),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _2522_ (.A1(net234),
    .A2(_0215_),
    .B1(_0208_),
    .Y(_0219_));
 sky130_fd_sc_hd__nor2_1 _2523_ (.A(_0218_),
    .B(_0219_),
    .Y(\d11.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2524_ (.A(\d11.count[5] ),
    .B(\d11.count[4] ),
    .C(_0215_),
    .X(_0220_));
 sky130_fd_sc_hd__o21ai_1 _2525_ (.A1(net175),
    .A2(_0218_),
    .B1(_0208_),
    .Y(_0221_));
 sky130_fd_sc_hd__nor2_1 _2526_ (.A(_0220_),
    .B(_0221_),
    .Y(\d11.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2527_ (.A(\d11.count[6] ),
    .B(_0220_),
    .X(_0222_));
 sky130_fd_sc_hd__o21ai_1 _2528_ (.A1(net159),
    .A2(_0220_),
    .B1(_0208_),
    .Y(_0223_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(_0222_),
    .B(_0223_),
    .Y(\d11.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2530_ (.A(\d11.count[7] ),
    .B(_0222_),
    .Y(_0224_));
 sky130_fd_sc_hd__or2_1 _2531_ (.A(\d11.count[7] ),
    .B(_0222_),
    .X(_0225_));
 sky130_fd_sc_hd__and3_1 _2532_ (.A(_0208_),
    .B(_0224_),
    .C(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _2533_ (.A(_0226_),
    .X(\d11.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2534_ (.A(\d11.count[8] ),
    .B(_0224_),
    .Y(_0227_));
 sky130_fd_sc_hd__and2_1 _2535_ (.A(_0208_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_1 _2536_ (.A(_0228_),
    .X(\d11.nxt_count[8] ));
 sky130_fd_sc_hd__a21o_1 _2537_ (.A1(\d12.count[8] ),
    .A2(_1715_),
    .B1(\d12.count[9] ),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\d12.count[5] ),
    .A1(\d12.count[6] ),
    .S(_1872_),
    .X(_0230_));
 sky130_fd_sc_hd__o22a_1 _2539_ (.A1(\d12.count[4] ),
    .A2(_1723_),
    .B1(_1777_),
    .B2(\d12.count[3] ),
    .X(_0231_));
 sky130_fd_sc_hd__a221o_1 _2540_ (.A1(_1872_),
    .A2(\d12.count[5] ),
    .B1(\d12.count[4] ),
    .B2(_1723_),
    .C1(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__and2_1 _2541_ (.A(_1727_),
    .B(\d12.count[6] ),
    .X(_0233_));
 sky130_fd_sc_hd__a221o_1 _2542_ (.A1(\d12.count[7] ),
    .A2(_1720_),
    .B1(_0230_),
    .B2(_0232_),
    .C1(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__o221a_1 _2543_ (.A1(\d12.count[8] ),
    .A2(_1805_),
    .B1(_1720_),
    .B2(\d12.count[7] ),
    .C1(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__nor2_2 _2544_ (.A(_0229_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _2545_ (.A(net84),
    .B(_0236_),
    .Y(\d12.nxt_count[0] ));
 sky130_fd_sc_hd__nand2_1 _2546_ (.A(\d12.count[1] ),
    .B(\d12.count[0] ),
    .Y(_0237_));
 sky130_fd_sc_hd__or2_1 _2547_ (.A(\d12.count[1] ),
    .B(\d12.count[0] ),
    .X(_0238_));
 sky130_fd_sc_hd__and3_1 _2548_ (.A(_0236_),
    .B(_0237_),
    .C(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_0239_),
    .X(\d12.nxt_count[1] ));
 sky130_fd_sc_hd__nand3_1 _2550_ (.A(\d12.count[1] ),
    .B(\d12.count[0] ),
    .C(\d12.count[2] ),
    .Y(_0240_));
 sky130_fd_sc_hd__a21o_1 _2551_ (.A1(\d12.count[1] ),
    .A2(\d12.count[0] ),
    .B1(\d12.count[2] ),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _2552_ (.A(_0236_),
    .B(_0240_),
    .C(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__clkbuf_1 _2553_ (.A(_0242_),
    .X(\d12.nxt_count[2] ));
 sky130_fd_sc_hd__and4_1 _2554_ (.A(\d12.count[1] ),
    .B(\d12.count[0] ),
    .C(\d12.count[3] ),
    .D(\d12.count[2] ),
    .X(_0243_));
 sky130_fd_sc_hd__a31o_1 _2555_ (.A1(\d12.count[1] ),
    .A2(\d12.count[0] ),
    .A3(\d12.count[2] ),
    .B1(\d12.count[3] ),
    .X(_0244_));
 sky130_fd_sc_hd__and3b_1 _2556_ (.A_N(_0243_),
    .B(_0244_),
    .C(_0236_),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_1 _2557_ (.A(_0245_),
    .X(\d12.nxt_count[3] ));
 sky130_fd_sc_hd__o21ai_1 _2558_ (.A1(net100),
    .A2(_0243_),
    .B1(_0236_),
    .Y(_0246_));
 sky130_fd_sc_hd__a21oi_1 _2559_ (.A1(net100),
    .A2(_0243_),
    .B1(_0246_),
    .Y(\d12.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2560_ (.A(\d12.count[5] ),
    .B(\d12.count[4] ),
    .C(_0243_),
    .X(_0247_));
 sky130_fd_sc_hd__a21o_1 _2561_ (.A1(\d12.count[4] ),
    .A2(_0243_),
    .B1(\d12.count[5] ),
    .X(_0248_));
 sky130_fd_sc_hd__and3b_1 _2562_ (.A_N(_0247_),
    .B(_0248_),
    .C(_0236_),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_1 _2563_ (.A(_0249_),
    .X(\d12.nxt_count[5] ));
 sky130_fd_sc_hd__o21ai_1 _2564_ (.A1(\d12.count[6] ),
    .A2(_0247_),
    .B1(_0236_),
    .Y(_0250_));
 sky130_fd_sc_hd__a21oi_1 _2565_ (.A1(net137),
    .A2(_0247_),
    .B1(_0250_),
    .Y(\d12.nxt_count[6] ));
 sky130_fd_sc_hd__nand3_1 _2566_ (.A(\d12.count[7] ),
    .B(\d12.count[6] ),
    .C(_0247_),
    .Y(_0251_));
 sky130_fd_sc_hd__a21o_1 _2567_ (.A1(\d12.count[6] ),
    .A2(_0247_),
    .B1(\d12.count[7] ),
    .X(_0252_));
 sky130_fd_sc_hd__and3_1 _2568_ (.A(_0236_),
    .B(_0251_),
    .C(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_1 _2569_ (.A(_0253_),
    .X(\d12.nxt_count[7] ));
 sky130_fd_sc_hd__inv_2 _2570_ (.A(net185),
    .Y(_0254_));
 sky130_fd_sc_hd__a21boi_1 _2571_ (.A1(_0254_),
    .A2(_0251_),
    .B1_N(_0236_),
    .Y(\d12.nxt_count[8] ));
 sky130_fd_sc_hd__o22a_1 _2572_ (.A1(\d13.count[8] ),
    .A2(_1714_),
    .B1(_1718_),
    .B2(\d13.count[7] ),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_1 _2573_ (.A1(\d13.count[7] ),
    .A2(_1717_),
    .B1(_1722_),
    .B2(\d13.count[6] ),
    .X(_0256_));
 sky130_fd_sc_hd__o22a_1 _2574_ (.A1(\d13.count[1] ),
    .A2(_1723_),
    .B1(_1777_),
    .B2(\d13.count[0] ),
    .X(_0257_));
 sky130_fd_sc_hd__or2_1 _2575_ (.A(\d13.count[1] ),
    .B(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__a21o_1 _2576_ (.A1(_1727_),
    .A2(\d13.count[2] ),
    .B1(\d13.count[3] ),
    .X(_0259_));
 sky130_fd_sc_hd__o21ai_1 _2577_ (.A1(_1727_),
    .A2(\d13.count[2] ),
    .B1(\d13.count[3] ),
    .Y(_0260_));
 sky130_fd_sc_hd__a21bo_1 _2578_ (.A1(_0258_),
    .A2(_0259_),
    .B1_N(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__o21a_1 _2579_ (.A1(\d13.count[4] ),
    .A2(_1720_),
    .B1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__a221o_1 _2580_ (.A1(\d13.count[4] ),
    .A2(_1720_),
    .B1(_1726_),
    .B2(\d13.count[5] ),
    .C1(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__o221a_1 _2581_ (.A1(\d13.count[6] ),
    .A2(_1723_),
    .B1(_1726_),
    .B2(\d13.count[5] ),
    .C1(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _2582_ (.A(_0256_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__a221oi_4 _2583_ (.A1(\d13.count[8] ),
    .A2(_1805_),
    .B1(_0255_),
    .B2(_0265_),
    .C1(\d13.count[9] ),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _2584_ (.A(net71),
    .B(_0266_),
    .Y(\d13.nxt_count[0] ));
 sky130_fd_sc_hd__or2_1 _2585_ (.A(\d13.count[0] ),
    .B(\d13.count[1] ),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _2586_ (.A(\d13.count[0] ),
    .B(\d13.count[1] ),
    .Y(_0268_));
 sky130_fd_sc_hd__and3_1 _2587_ (.A(_0266_),
    .B(_0267_),
    .C(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_1 _2588_ (.A(_0269_),
    .X(\d13.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2589_ (.A(\d13.count[0] ),
    .B(\d13.count[1] ),
    .C(\d13.count[2] ),
    .X(_0270_));
 sky130_fd_sc_hd__a21o_1 _2590_ (.A1(\d13.count[0] ),
    .A2(\d13.count[1] ),
    .B1(\d13.count[2] ),
    .X(_0271_));
 sky130_fd_sc_hd__and3b_1 _2591_ (.A_N(_0270_),
    .B(_0271_),
    .C(_0266_),
    .X(_0272_));
 sky130_fd_sc_hd__clkbuf_1 _2592_ (.A(_0272_),
    .X(\d13.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2593_ (.A(\d13.count[3] ),
    .B(_0270_),
    .X(_0273_));
 sky130_fd_sc_hd__or2_1 _2594_ (.A(\d13.count[3] ),
    .B(_0270_),
    .X(_0274_));
 sky130_fd_sc_hd__and3b_1 _2595_ (.A_N(_0273_),
    .B(_0274_),
    .C(_0266_),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _2596_ (.A(_0275_),
    .X(\d13.nxt_count[3] ));
 sky130_fd_sc_hd__and3_1 _2597_ (.A(\d13.count[3] ),
    .B(\d13.count[4] ),
    .C(_0270_),
    .X(_0276_));
 sky130_fd_sc_hd__o21ai_1 _2598_ (.A1(net215),
    .A2(_0273_),
    .B1(_0266_),
    .Y(_0277_));
 sky130_fd_sc_hd__nor2_1 _2599_ (.A(_0276_),
    .B(_0277_),
    .Y(\d13.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2600_ (.A(\d13.count[5] ),
    .B(\d13.count[4] ),
    .C(_0273_),
    .X(_0278_));
 sky130_fd_sc_hd__o21ai_1 _2601_ (.A1(\d13.count[5] ),
    .A2(_0276_),
    .B1(_0266_),
    .Y(_0279_));
 sky130_fd_sc_hd__nor2_1 _2602_ (.A(_0278_),
    .B(_0279_),
    .Y(\d13.nxt_count[5] ));
 sky130_fd_sc_hd__and2_1 _2603_ (.A(\d13.count[6] ),
    .B(_0278_),
    .X(_0280_));
 sky130_fd_sc_hd__o21ai_1 _2604_ (.A1(\d13.count[6] ),
    .A2(_0278_),
    .B1(_0266_),
    .Y(_0281_));
 sky130_fd_sc_hd__nor2_1 _2605_ (.A(_0280_),
    .B(_0281_),
    .Y(\d13.nxt_count[6] ));
 sky130_fd_sc_hd__nand2_1 _2606_ (.A(\d13.count[7] ),
    .B(_0280_),
    .Y(_0282_));
 sky130_fd_sc_hd__or2_1 _2607_ (.A(\d13.count[7] ),
    .B(_0280_),
    .X(_0283_));
 sky130_fd_sc_hd__and3_1 _2608_ (.A(_0266_),
    .B(_0282_),
    .C(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__clkbuf_1 _2609_ (.A(_0284_),
    .X(\d13.nxt_count[7] ));
 sky130_fd_sc_hd__xnor2_1 _2610_ (.A(\d13.count[8] ),
    .B(_0282_),
    .Y(_0285_));
 sky130_fd_sc_hd__and2_1 _2611_ (.A(_0266_),
    .B(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _2612_ (.A(_0286_),
    .X(\d13.nxt_count[8] ));
 sky130_fd_sc_hd__inv_2 _2613_ (.A(net90),
    .Y(\p0.nxt_count[0] ));
 sky130_fd_sc_hd__xor2_1 _2614_ (.A(net134),
    .B(net90),
    .X(\p0.nxt_count[1] ));
 sky130_fd_sc_hd__and3_1 _2615_ (.A(\p0.count[2] ),
    .B(\p0.count[1] ),
    .C(\p0.count[0] ),
    .X(_0287_));
 sky130_fd_sc_hd__a21oi_1 _2616_ (.A1(\p0.count[1] ),
    .A2(\p0.count[0] ),
    .B1(net126),
    .Y(_0288_));
 sky130_fd_sc_hd__nor2_1 _2617_ (.A(_0287_),
    .B(net127),
    .Y(\p0.nxt_count[2] ));
 sky130_fd_sc_hd__and2_1 _2618_ (.A(\p0.count[3] ),
    .B(_0287_),
    .X(_0289_));
 sky130_fd_sc_hd__nor2_1 _2619_ (.A(net132),
    .B(_0287_),
    .Y(_0290_));
 sky130_fd_sc_hd__nor2_1 _2620_ (.A(_0289_),
    .B(_0290_),
    .Y(\p0.nxt_count[3] ));
 sky130_fd_sc_hd__inv_2 _2621_ (.A(net225),
    .Y(_0291_));
 sky130_fd_sc_hd__xnor2_1 _2622_ (.A(_0291_),
    .B(_0289_),
    .Y(\p0.nxt_count[4] ));
 sky130_fd_sc_hd__and3_1 _2623_ (.A(\p0.count[4] ),
    .B(\p0.count[5] ),
    .C(_0289_),
    .X(_0292_));
 sky130_fd_sc_hd__a21oi_1 _2624_ (.A1(\p0.count[4] ),
    .A2(_0289_),
    .B1(net121),
    .Y(_0293_));
 sky130_fd_sc_hd__nor2_1 _2625_ (.A(_0292_),
    .B(net122),
    .Y(\p0.nxt_count[5] ));
 sky130_fd_sc_hd__nand2_1 _2626_ (.A(\p0.count[6] ),
    .B(_0292_),
    .Y(_0294_));
 sky130_fd_sc_hd__or2_1 _2627_ (.A(\p0.count[6] ),
    .B(_0292_),
    .X(_0295_));
 sky130_fd_sc_hd__and2_1 _2628_ (.A(_0294_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _2629_ (.A(_0296_),
    .X(\p0.nxt_count[6] ));
 sky130_fd_sc_hd__xnor2_1 _2630_ (.A(net81),
    .B(_0294_),
    .Y(\p0.nxt_count[7] ));
 sky130_fd_sc_hd__or2b_1 _2631_ (.A(net220),
    .B_N(\m0.edgy.in ),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_1 _2632_ (.A(_1872_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__or2_1 _2633_ (.A(_1872_),
    .B(_0297_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _2634_ (.A(_0298_),
    .B(_0299_),
    .Y(\e0.next_q[0] ));
 sky130_fd_sc_hd__a22o_1 _2635_ (.A1(_1724_),
    .A2(_0297_),
    .B1(_0298_),
    .B2(_1726_),
    .X(\e0.next_q[1] ));
 sky130_fd_sc_hd__clkbuf_8 _2636_ (.A(\s0.type_switch[0] ),
    .X(_0300_));
 sky130_fd_sc_hd__buf_12 _2637_ (.A(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__and2b_1 _2638_ (.A_N(\m0.edgo.delay ),
    .B(\m0.edgo.in ),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _2639_ (.A(_0301_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__or2_1 _2640_ (.A(_0301_),
    .B(_0302_),
    .X(_0304_));
 sky130_fd_sc_hd__and2_1 _2641_ (.A(_0303_),
    .B(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _2642_ (.A(_0305_),
    .X(\s0.next_q[0] ));
 sky130_fd_sc_hd__buf_4 _2643_ (.A(\s0.type_switch[1] ),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_16 _2644_ (.A(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__and2b_1 _2645_ (.A_N(_0306_),
    .B(_0300_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_4 _2646_ (.A(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_8 _2647_ (.A(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _2648_ (.A1(_0307_),
    .A2(_0303_),
    .B1(_0310_),
    .B2(_0302_),
    .X(\s0.next_q[1] ));
 sky130_fd_sc_hd__inv_2 _2649_ (.A(\p0.count[7] ),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _2650_ (.A(\p0.count[6] ),
    .Y(_0312_));
 sky130_fd_sc_hd__or2_1 _2651_ (.A(_0312_),
    .B(\em0.mixed_sample[6] ),
    .X(_0313_));
 sky130_fd_sc_hd__inv_2 _2652_ (.A(\p0.count[5] ),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _2653_ (.A(\p0.count[3] ),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _2654_ (.A(\p0.count[2] ),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _2655_ (.A(\p0.count[1] ),
    .Y(_0317_));
 sky130_fd_sc_hd__or2_1 _2656_ (.A(_0317_),
    .B(\em0.mixed_sample[1] ),
    .X(_0318_));
 sky130_fd_sc_hd__a22o_1 _2657_ (.A1(_0316_),
    .A2(\em0.mixed_sample[2] ),
    .B1(\em0.mixed_sample[1] ),
    .B2(_0317_),
    .X(_0319_));
 sky130_fd_sc_hd__a31o_1 _2658_ (.A1(\p0.nxt_count[0] ),
    .A2(\em0.mixed_sample[0] ),
    .A3(_0318_),
    .B1(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__o221a_1 _2659_ (.A1(_0315_),
    .A2(\em0.mixed_sample[3] ),
    .B1(\em0.mixed_sample[2] ),
    .B2(_0316_),
    .C1(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__a221o_1 _2660_ (.A1(_0291_),
    .A2(\em0.mixed_sample[4] ),
    .B1(\em0.mixed_sample[3] ),
    .B2(_0315_),
    .C1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__o221a_1 _2661_ (.A1(_0314_),
    .A2(\em0.mixed_sample[5] ),
    .B1(\em0.mixed_sample[4] ),
    .B2(_0291_),
    .C1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__a221o_1 _2662_ (.A1(_0312_),
    .A2(\em0.mixed_sample[6] ),
    .B1(\em0.mixed_sample[5] ),
    .B2(_0314_),
    .C1(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _2663_ (.A1(_0311_),
    .A2(\em0.mixed_sample[7] ),
    .B1(_0313_),
    .B2(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__o21a_1 _2664_ (.A1(_0311_),
    .A2(net113),
    .B1(_0325_),
    .X(\p0.pwm ));
 sky130_fd_sc_hd__inv_2 _2665_ (.A(\em0.u1.state[1] ),
    .Y(_0326_));
 sky130_fd_sc_hd__nor2_1 _2666_ (.A(_0326_),
    .B(_1711_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _2667_ (.A(\em0.u1.state[2] ),
    .Y(_0327_));
 sky130_fd_sc_hd__buf_4 _2668_ (.A(net10),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_8 _2669_ (.A(net7),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_8 _2670_ (.A(net3),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _2671_ (.A(_0329_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__or2_1 _2672_ (.A(_0329_),
    .B(_0330_),
    .X(_0332_));
 sky130_fd_sc_hd__inv_2 _2673_ (.A(net12),
    .Y(_0333_));
 sky130_fd_sc_hd__clkbuf_4 _2674_ (.A(net4),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_4 _2675_ (.A(net14),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_4 _2676_ (.A(net15),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_4 _2677_ (.A(net13),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _2678_ (.A(_0336_),
    .B(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__nand2_1 _2679_ (.A(_0336_),
    .B(_0337_),
    .Y(_0339_));
 sky130_fd_sc_hd__clkbuf_4 _2680_ (.A(net5),
    .X(_0340_));
 sky130_fd_sc_hd__a21o_1 _2681_ (.A1(_0338_),
    .A2(_0339_),
    .B1(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__nand3_1 _2682_ (.A(_0340_),
    .B(_0338_),
    .C(_0339_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _2683_ (.A(_0341_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__clkbuf_4 _2684_ (.A(net6),
    .X(_0344_));
 sky130_fd_sc_hd__inv_2 _2685_ (.A(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__clkbuf_4 _2686_ (.A(net11),
    .X(_0346_));
 sky130_fd_sc_hd__buf_4 _2687_ (.A(net9),
    .X(_0347_));
 sky130_fd_sc_hd__buf_4 _2688_ (.A(net8),
    .X(_0348_));
 sky130_fd_sc_hd__or2_1 _2689_ (.A(_0347_),
    .B(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _2690_ (.A(_0347_),
    .B(_0348_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _2691_ (.A(_0349_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__xor2_1 _2692_ (.A(_0346_),
    .B(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__xnor2_1 _2693_ (.A(_0345_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _2694_ (.A(_0343_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__or2_1 _2695_ (.A(_0343_),
    .B(_0353_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _2696_ (.A(_0354_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _2697_ (.A(_0335_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_1 _2698_ (.A(_0335_),
    .B(_0356_),
    .Y(_0358_));
 sky130_fd_sc_hd__and2_1 _2699_ (.A(_0357_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _2700_ (.A(_0334_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__nand2_1 _2701_ (.A(_0334_),
    .B(_0359_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _2702_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__nor2_1 _2703_ (.A(_0333_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__and2_1 _2704_ (.A(_0333_),
    .B(_0362_),
    .X(_0364_));
 sky130_fd_sc_hd__o2bb2a_1 _2705_ (.A1_N(_0331_),
    .A2_N(_0332_),
    .B1(_0363_),
    .B2(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _2706_ (.A(_0363_),
    .B(_0364_),
    .X(_0366_));
 sky130_fd_sc_hd__and3b_1 _2707_ (.A_N(_0366_),
    .B(_0332_),
    .C(_0331_),
    .X(_0367_));
 sky130_fd_sc_hd__nor2_2 _2708_ (.A(_0365_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _2709_ (.A(_0328_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__o21a_1 _2710_ (.A1(_0328_),
    .A2(_0368_),
    .B1(\em0.u1.state[2] ),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _2711_ (.A1(_0327_),
    .A2(net147),
    .B1(_0369_),
    .B2(_0370_),
    .X(_0003_));
 sky130_fd_sc_hd__a21bo_1 _2712_ (.A1(_0346_),
    .A2(_0349_),
    .B1_N(_0350_),
    .X(_0371_));
 sky130_fd_sc_hd__and3_1 _2713_ (.A(_0329_),
    .B(_0330_),
    .C(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__and2b_1 _2714_ (.A_N(_0371_),
    .B(_0331_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _2715_ (.A(_0372_),
    .B(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__o21a_1 _2716_ (.A1(_0345_),
    .A2(_0352_),
    .B1(_0355_),
    .X(_0375_));
 sky130_fd_sc_hd__xnor2_1 _2717_ (.A(_0374_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__a21oi_1 _2718_ (.A1(_0339_),
    .A2(_0342_),
    .B1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__and3_1 _2719_ (.A(_0339_),
    .B(_0342_),
    .C(_0376_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_1 _2720_ (.A(_0377_),
    .B(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__a21oi_2 _2721_ (.A1(_0358_),
    .A2(_0361_),
    .B1(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__and3_1 _2722_ (.A(_0358_),
    .B(_0361_),
    .C(_0379_),
    .X(_0381_));
 sky130_fd_sc_hd__nor2_1 _2723_ (.A(_0380_),
    .B(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__o21a_1 _2724_ (.A1(_0363_),
    .A2(_0367_),
    .B1(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__nor3_1 _2725_ (.A(_0363_),
    .B(_0367_),
    .C(_0382_),
    .Y(_0384_));
 sky130_fd_sc_hd__or2_1 _2726_ (.A(_0383_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__a21o_1 _2727_ (.A1(_0369_),
    .A2(_0385_),
    .B1(_0327_),
    .X(_0386_));
 sky130_fd_sc_hd__nor2_1 _2728_ (.A(_0369_),
    .B(_0385_),
    .Y(_0387_));
 sky130_fd_sc_hd__a2bb2o_1 _2729_ (.A1_N(_0386_),
    .A2_N(_0387_),
    .B1(net116),
    .B2(_0327_),
    .X(_0004_));
 sky130_fd_sc_hd__xnor2_1 _2730_ (.A(_0372_),
    .B(_0377_),
    .Y(_0388_));
 sky130_fd_sc_hd__o21ai_2 _2731_ (.A1(_0374_),
    .A2(_0375_),
    .B1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__xor2_2 _2732_ (.A(_0380_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__o21ai_1 _2733_ (.A1(_0383_),
    .A2(_0387_),
    .B1(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__o31a_1 _2734_ (.A1(_0383_),
    .A2(_0387_),
    .A3(_0390_),
    .B1(\em0.u1.state[2] ),
    .X(_0392_));
 sky130_fd_sc_hd__a22o_1 _2735_ (.A1(_0327_),
    .A2(net244),
    .B1(_0391_),
    .B2(_0392_),
    .X(_0005_));
 sky130_fd_sc_hd__nand2_1 _2736_ (.A(\em0.u1.state[2] ),
    .B(_0391_),
    .Y(_0393_));
 sky130_fd_sc_hd__a22o_1 _2737_ (.A1(_0372_),
    .A2(_0377_),
    .B1(_0380_),
    .B2(_0389_),
    .X(_0394_));
 sky130_fd_sc_hd__o22a_1 _2738_ (.A1(\em0.u1.state[2] ),
    .A2(net158),
    .B1(_0393_),
    .B2(_0394_),
    .X(_0006_));
 sky130_fd_sc_hd__and2_1 _2739_ (.A(_0327_),
    .B(\em0.u1.D[12] ),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _2740_ (.A(_0395_),
    .X(_0007_));
 sky130_fd_sc_hd__o2bb2a_1 _2741_ (.A1_N(\d13.count[1] ),
    .A2_N(_1723_),
    .B1(_1718_),
    .B2(\d13.count[4] ),
    .X(_0396_));
 sky130_fd_sc_hd__o2bb2a_1 _2742_ (.A1_N(\d13.count[4] ),
    .A2_N(_1718_),
    .B1(_1722_),
    .B2(\d13.count[6] ),
    .X(_0397_));
 sky130_fd_sc_hd__a211o_1 _2743_ (.A1(\d13.count[8] ),
    .A2(_1714_),
    .B1(_0256_),
    .C1(\d13.count[9] ),
    .X(_0398_));
 sky130_fd_sc_hd__a21oi_1 _2744_ (.A1(\d13.count[0] ),
    .A2(_1732_),
    .B1(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__and3_1 _2745_ (.A(_0255_),
    .B(_0397_),
    .C(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__xnor2_1 _2746_ (.A(\d13.count[5] ),
    .B(_1733_),
    .Y(_0401_));
 sky130_fd_sc_hd__and4_1 _2747_ (.A(_0257_),
    .B(_0396_),
    .C(_0400_),
    .D(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__and3_1 _2748_ (.A(_0260_),
    .B(_0259_),
    .C(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__and4_1 _2749_ (.A(\d13.saw_temp[6] ),
    .B(\d13.saw_temp[5] ),
    .C(\d13.saw_temp[2] ),
    .D(\d13.saw_temp[1] ),
    .X(_0404_));
 sky130_fd_sc_hd__and4_1 _2750_ (.A(\d13.saw_temp[4] ),
    .B(\d13.saw_temp[3] ),
    .C(\d13.saw_temp[0] ),
    .D(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _2751_ (.A(\d13.saw_temp[7] ),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__o21a_1 _2752_ (.A1(_0406_),
    .A2(_0403_),
    .B1(\d13.saw_temp[0] ),
    .X(_0407_));
 sky130_fd_sc_hd__o21ba_1 _2753_ (.A1(net191),
    .A2(_0403_),
    .B1_N(_0407_),
    .X(_0008_));
 sky130_fd_sc_hd__xor2_1 _2754_ (.A(net153),
    .B(_0407_),
    .X(_0009_));
 sky130_fd_sc_hd__a21oi_1 _2755_ (.A1(\d13.saw_temp[1] ),
    .A2(_0407_),
    .B1(net219),
    .Y(_0408_));
 sky130_fd_sc_hd__and3_1 _2756_ (.A(\d13.saw_temp[2] ),
    .B(\d13.saw_temp[1] ),
    .C(_0407_),
    .X(_0409_));
 sky130_fd_sc_hd__nor2_1 _2757_ (.A(_0408_),
    .B(_0409_),
    .Y(_0010_));
 sky130_fd_sc_hd__xor2_1 _2758_ (.A(net145),
    .B(_0409_),
    .X(_0011_));
 sky130_fd_sc_hd__a21oi_1 _2759_ (.A1(\d13.saw_temp[3] ),
    .A2(_0409_),
    .B1(net210),
    .Y(_0410_));
 sky130_fd_sc_hd__and3_1 _2760_ (.A(\d13.saw_temp[4] ),
    .B(\d13.saw_temp[3] ),
    .C(_0409_),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _2761_ (.A(_0410_),
    .B(_0411_),
    .Y(_0012_));
 sky130_fd_sc_hd__or2_1 _2762_ (.A(\d13.saw_temp[5] ),
    .B(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__nand2_1 _2763_ (.A(\d13.saw_temp[5] ),
    .B(_0411_),
    .Y(_0413_));
 sky130_fd_sc_hd__and2_1 _2764_ (.A(_0412_),
    .B(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _2765_ (.A(_0414_),
    .X(_0013_));
 sky130_fd_sc_hd__xnor2_1 _2766_ (.A(net115),
    .B(_0413_),
    .Y(_0014_));
 sky130_fd_sc_hd__a21oi_1 _2767_ (.A1(_0405_),
    .A2(_0403_),
    .B1(\d13.saw_temp[7] ),
    .Y(_0415_));
 sky130_fd_sc_hd__nor2_1 _2768_ (.A(_0406_),
    .B(_0415_),
    .Y(_0015_));
 sky130_fd_sc_hd__or4bb_1 _2769_ (.A(_1767_),
    .B(_1770_),
    .C_N(_1771_),
    .D_N(_1776_),
    .X(_0416_));
 sky130_fd_sc_hd__o21a_1 _2770_ (.A1(\d2.count[1] ),
    .A2(\d2.count[6] ),
    .B1(_1732_),
    .X(_0417_));
 sky130_fd_sc_hd__o21ai_1 _2771_ (.A1(\d2.count[8] ),
    .A2(_1717_),
    .B1(_1768_),
    .Y(_0418_));
 sky130_fd_sc_hd__a2111o_1 _2772_ (.A1(_1712_),
    .A2(\d2.count[2] ),
    .B1(_1782_),
    .C1(_0418_),
    .D1(\d2.count[0] ),
    .X(_0419_));
 sky130_fd_sc_hd__or4_1 _2773_ (.A(_1779_),
    .B(_1773_),
    .C(_0417_),
    .D(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_2 _2774_ (.A(_0416_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__and4_1 _2775_ (.A(\d2.saw_temp[6] ),
    .B(\d2.saw_temp[5] ),
    .C(\d2.saw_temp[2] ),
    .D(\d2.saw_temp[1] ),
    .X(_0422_));
 sky130_fd_sc_hd__and4_1 _2776_ (.A(\d2.saw_temp[4] ),
    .B(\d2.saw_temp[3] ),
    .C(\d2.saw_temp[0] ),
    .D(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _2777_ (.A(\d2.saw_temp[7] ),
    .B(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__o21ai_2 _2778_ (.A1(_0424_),
    .A2(_0421_),
    .B1(\d2.saw_temp[0] ),
    .Y(_0425_));
 sky130_fd_sc_hd__o21a_1 _2779_ (.A1(net235),
    .A2(_0421_),
    .B1(_0425_),
    .X(_0016_));
 sky130_fd_sc_hd__xnor2_1 _2780_ (.A(net170),
    .B(_0425_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _2781_ (.A(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21oi_1 _2782_ (.A1(\d2.saw_temp[1] ),
    .A2(_0426_),
    .B1(net207),
    .Y(_0427_));
 sky130_fd_sc_hd__and3_1 _2783_ (.A(\d2.saw_temp[2] ),
    .B(\d2.saw_temp[1] ),
    .C(_0426_),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_1 _2784_ (.A(_0427_),
    .B(_0428_),
    .Y(_0018_));
 sky130_fd_sc_hd__xor2_1 _2785_ (.A(net174),
    .B(_0428_),
    .X(_0019_));
 sky130_fd_sc_hd__a21oi_1 _2786_ (.A1(\d2.saw_temp[3] ),
    .A2(_0428_),
    .B1(net218),
    .Y(_0429_));
 sky130_fd_sc_hd__and3_1 _2787_ (.A(\d2.saw_temp[4] ),
    .B(\d2.saw_temp[3] ),
    .C(_0428_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_1 _2788_ (.A(_0429_),
    .B(_0430_),
    .Y(_0020_));
 sky130_fd_sc_hd__or2_1 _2789_ (.A(\d2.saw_temp[5] ),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__nand2_1 _2790_ (.A(\d2.saw_temp[5] ),
    .B(_0430_),
    .Y(_0432_));
 sky130_fd_sc_hd__and2_1 _2791_ (.A(_0431_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _2792_ (.A(_0433_),
    .X(_0021_));
 sky130_fd_sc_hd__xnor2_1 _2793_ (.A(net123),
    .B(_0432_),
    .Y(_0022_));
 sky130_fd_sc_hd__a21oi_1 _2794_ (.A1(_0423_),
    .A2(_0421_),
    .B1(\d2.saw_temp[7] ),
    .Y(_0434_));
 sky130_fd_sc_hd__nor2_1 _2795_ (.A(_0424_),
    .B(_0434_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _2796_ (.A(net239),
    .Y(_0435_));
 sky130_fd_sc_hd__a21o_1 _2797_ (.A1(\d3.count[2] ),
    .A2(_1733_),
    .B1(_1807_),
    .X(_0436_));
 sky130_fd_sc_hd__a2111o_1 _2798_ (.A1(_1735_),
    .A2(\d3.count[1] ),
    .B1(\d3.count[5] ),
    .C1(_1810_),
    .D1(_1813_),
    .X(_0437_));
 sky130_fd_sc_hd__a211o_1 _2799_ (.A1(\d3.count[0] ),
    .A2(_1732_),
    .B1(_1812_),
    .C1(_1815_),
    .X(_0438_));
 sky130_fd_sc_hd__o22a_1 _2800_ (.A1(\d3.count[9] ),
    .A2(_1714_),
    .B1(_1732_),
    .B2(\d3.count[6] ),
    .X(_0439_));
 sky130_fd_sc_hd__or4b_1 _2801_ (.A(_1809_),
    .B(_1817_),
    .C(_0438_),
    .D_N(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__or4_2 _2802_ (.A(_1806_),
    .B(_0436_),
    .C(_0437_),
    .D(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__and3_1 _2803_ (.A(\d3.saw_temp[4] ),
    .B(\d3.saw_temp[3] ),
    .C(\d3.saw_temp[0] ),
    .X(_0442_));
 sky130_fd_sc_hd__and4_1 _2804_ (.A(\d3.saw_temp[6] ),
    .B(\d3.saw_temp[5] ),
    .C(\d3.saw_temp[2] ),
    .D(\d3.saw_temp[1] ),
    .X(_0443_));
 sky130_fd_sc_hd__and3_1 _2805_ (.A(\d3.saw_temp[7] ),
    .B(_0442_),
    .C(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__or2b_1 _2806_ (.A(_0444_),
    .B_N(_0441_),
    .X(_0445_));
 sky130_fd_sc_hd__and2_1 _2807_ (.A(\d3.saw_temp[0] ),
    .B(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__a21oi_1 _2808_ (.A1(_0435_),
    .A2(_0441_),
    .B1(_0446_),
    .Y(_0024_));
 sky130_fd_sc_hd__xor2_1 _2809_ (.A(net160),
    .B(_0446_),
    .X(_0025_));
 sky130_fd_sc_hd__a21oi_1 _2810_ (.A1(\d3.saw_temp[1] ),
    .A2(_0446_),
    .B1(net224),
    .Y(_0447_));
 sky130_fd_sc_hd__and3_1 _2811_ (.A(\d3.saw_temp[2] ),
    .B(\d3.saw_temp[1] ),
    .C(_0446_),
    .X(_0448_));
 sky130_fd_sc_hd__nor2_1 _2812_ (.A(_0447_),
    .B(_0448_),
    .Y(_0026_));
 sky130_fd_sc_hd__nor2_1 _2813_ (.A(net243),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__and2_1 _2814_ (.A(\d3.saw_temp[3] ),
    .B(_0448_),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_1 _2815_ (.A(_0449_),
    .B(_0450_),
    .Y(_0027_));
 sky130_fd_sc_hd__xor2_1 _2816_ (.A(net150),
    .B(_0450_),
    .X(_0028_));
 sky130_fd_sc_hd__a21oi_1 _2817_ (.A1(\d3.saw_temp[4] ),
    .A2(_0450_),
    .B1(net241),
    .Y(_0451_));
 sky130_fd_sc_hd__and3_1 _2818_ (.A(\d3.saw_temp[5] ),
    .B(\d3.saw_temp[4] ),
    .C(_0450_),
    .X(_0452_));
 sky130_fd_sc_hd__nor2_1 _2819_ (.A(_0451_),
    .B(_0452_),
    .Y(_0029_));
 sky130_fd_sc_hd__xor2_1 _2820_ (.A(net114),
    .B(_0452_),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_1 _2821_ (.A(_0442_),
    .B(_0443_),
    .Y(_0453_));
 sky130_fd_sc_hd__o21ba_1 _2822_ (.A1(_0453_),
    .A2(_0441_),
    .B1_N(\d3.saw_temp[7] ),
    .X(_0454_));
 sky130_fd_sc_hd__nor2_1 _2823_ (.A(_0444_),
    .B(_0454_),
    .Y(_0031_));
 sky130_fd_sc_hd__and4_1 _2824_ (.A(\d4.saw_temp[5] ),
    .B(\d4.saw_temp[4] ),
    .C(\d4.saw_temp[1] ),
    .D(\d4.saw_temp[2] ),
    .X(_0455_));
 sky130_fd_sc_hd__and4_1 _2825_ (.A(\d4.saw_temp[6] ),
    .B(\d4.saw_temp[0] ),
    .C(\d4.saw_temp[3] ),
    .D(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__and2_1 _2826_ (.A(\d4.saw_temp[7] ),
    .B(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__inv_2 _2827_ (.A(_1847_),
    .Y(_0458_));
 sky130_fd_sc_hd__a22o_1 _2828_ (.A1(\d4.count[2] ),
    .A2(_1724_),
    .B1(_1777_),
    .B2(\d4.count[0] ),
    .X(_0459_));
 sky130_fd_sc_hd__a221o_1 _2829_ (.A1(_1735_),
    .A2(\d4.count[1] ),
    .B1(_1869_),
    .B2(_1724_),
    .C1(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__a2111oi_4 _2830_ (.A1(\d4.count[8] ),
    .A2(_1805_),
    .B1(_0458_),
    .C1(_0460_),
    .D1(\d4.count[9] ),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_1 _2831_ (.A(_0457_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__xnor2_1 _2832_ (.A(net152),
    .B(_0462_),
    .Y(_0032_));
 sky130_fd_sc_hd__o211a_1 _2833_ (.A1(_0457_),
    .A2(_0461_),
    .B1(\d4.saw_temp[1] ),
    .C1(\d4.saw_temp[0] ),
    .X(_0463_));
 sky130_fd_sc_hd__inv_2 _2834_ (.A(\d4.saw_temp[0] ),
    .Y(_0464_));
 sky130_fd_sc_hd__o21ba_1 _2835_ (.A1(_0464_),
    .A2(_0462_),
    .B1_N(\d4.saw_temp[1] ),
    .X(_0465_));
 sky130_fd_sc_hd__nor2_1 _2836_ (.A(_0463_),
    .B(_0465_),
    .Y(_0033_));
 sky130_fd_sc_hd__and2_1 _2837_ (.A(\d4.saw_temp[2] ),
    .B(_0463_),
    .X(_0466_));
 sky130_fd_sc_hd__nor2_1 _2838_ (.A(net182),
    .B(_0463_),
    .Y(_0467_));
 sky130_fd_sc_hd__nor2_1 _2839_ (.A(_0466_),
    .B(_0467_),
    .Y(_0034_));
 sky130_fd_sc_hd__xor2_1 _2840_ (.A(net104),
    .B(_0466_),
    .X(_0035_));
 sky130_fd_sc_hd__and3_1 _2841_ (.A(\d4.saw_temp[4] ),
    .B(\d4.saw_temp[3] ),
    .C(_0466_),
    .X(_0468_));
 sky130_fd_sc_hd__a21oi_1 _2842_ (.A1(net104),
    .A2(_0466_),
    .B1(net161),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_1 _2843_ (.A(_0468_),
    .B(_0469_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand2_1 _2844_ (.A(\d4.saw_temp[5] ),
    .B(_0468_),
    .Y(_0470_));
 sky130_fd_sc_hd__or2_1 _2845_ (.A(\d4.saw_temp[5] ),
    .B(_0468_),
    .X(_0471_));
 sky130_fd_sc_hd__and2_1 _2846_ (.A(_0470_),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _2847_ (.A(_0472_),
    .X(_0037_));
 sky130_fd_sc_hd__xnor2_1 _2848_ (.A(net130),
    .B(_0470_),
    .Y(_0038_));
 sky130_fd_sc_hd__a21oi_1 _2849_ (.A1(_0456_),
    .A2(_0461_),
    .B1(\d4.saw_temp[7] ),
    .Y(_0473_));
 sky130_fd_sc_hd__nor2_1 _2850_ (.A(_0457_),
    .B(_0473_),
    .Y(_0039_));
 sky130_fd_sc_hd__a2bb2o_1 _2851_ (.A1_N(\d5.count[8] ),
    .A2_N(_1805_),
    .B1(_1735_),
    .B2(\d5.count[1] ),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_1 _2852_ (.A(_1945_),
    .B(_1877_),
    .Y(_0475_));
 sky130_fd_sc_hd__a211o_1 _2853_ (.A1(\d5.count[8] ),
    .A2(_1715_),
    .B1(_1871_),
    .C1(_1885_),
    .X(_0476_));
 sky130_fd_sc_hd__or4_1 _2854_ (.A(\d5.count[9] ),
    .B(_1876_),
    .C(_0475_),
    .D(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__a2111o_2 _2855_ (.A1(\d5.count[0] ),
    .A2(_1777_),
    .B1(_1882_),
    .C1(_0474_),
    .D1(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__inv_2 _2856_ (.A(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__and3_1 _2857_ (.A(\d5.saw_temp[4] ),
    .B(\d5.saw_temp[3] ),
    .C(\d5.saw_temp[0] ),
    .X(_0480_));
 sky130_fd_sc_hd__and2_1 _2858_ (.A(\d5.saw_temp[2] ),
    .B(\d5.saw_temp[1] ),
    .X(_0481_));
 sky130_fd_sc_hd__and4_1 _2859_ (.A(\d5.saw_temp[6] ),
    .B(\d5.saw_temp[5] ),
    .C(_0480_),
    .D(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _2860_ (.A(\d5.saw_temp[7] ),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__a21boi_2 _2861_ (.A1(_0483_),
    .A2(_0478_),
    .B1_N(\d5.saw_temp[0] ),
    .Y(_0484_));
 sky130_fd_sc_hd__o21ba_1 _2862_ (.A1(net196),
    .A2(_0479_),
    .B1_N(_0484_),
    .X(_0040_));
 sky130_fd_sc_hd__xor2_1 _2863_ (.A(net118),
    .B(_0484_),
    .X(_0041_));
 sky130_fd_sc_hd__a21oi_1 _2864_ (.A1(\d5.saw_temp[1] ),
    .A2(_0484_),
    .B1(net221),
    .Y(_0485_));
 sky130_fd_sc_hd__and2_1 _2865_ (.A(_0481_),
    .B(_0484_),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_1 _2866_ (.A(net222),
    .B(_0486_),
    .Y(_0042_));
 sky130_fd_sc_hd__nor2_1 _2867_ (.A(\d5.saw_temp[3] ),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__and3_1 _2868_ (.A(\d5.saw_temp[3] ),
    .B(_0481_),
    .C(_0484_),
    .X(_0488_));
 sky130_fd_sc_hd__nor2_1 _2869_ (.A(_0487_),
    .B(_0488_),
    .Y(_0043_));
 sky130_fd_sc_hd__nor2_1 _2870_ (.A(net229),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__and2_1 _2871_ (.A(\d5.saw_temp[4] ),
    .B(_0488_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_1 _2872_ (.A(_0489_),
    .B(_0490_),
    .Y(_0044_));
 sky130_fd_sc_hd__or2_1 _2873_ (.A(\d5.saw_temp[5] ),
    .B(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_1 _2874_ (.A(\d5.saw_temp[5] ),
    .B(_0490_),
    .Y(_0492_));
 sky130_fd_sc_hd__and2_1 _2875_ (.A(_0491_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _2876_ (.A(_0493_),
    .X(_0045_));
 sky130_fd_sc_hd__xnor2_1 _2877_ (.A(net105),
    .B(_0492_),
    .Y(_0046_));
 sky130_fd_sc_hd__a21o_1 _2878_ (.A1(_0482_),
    .A2(_0479_),
    .B1(\d5.saw_temp[7] ),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _2879_ (.A(_0483_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _2880_ (.A(_0495_),
    .X(_0047_));
 sky130_fd_sc_hd__a2111oi_1 _2881_ (.A1(\d6.count[3] ),
    .A2(_1777_),
    .B1(_1919_),
    .C1(_1923_),
    .D1(\d6.count[2] ),
    .Y(_0496_));
 sky130_fd_sc_hd__and3b_1 _2882_ (.A_N(_1918_),
    .B(_1921_),
    .C(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__and4_1 _2883_ (.A(\d6.saw_temp[6] ),
    .B(\d6.saw_temp[5] ),
    .C(\d6.saw_temp[2] ),
    .D(\d6.saw_temp[1] ),
    .X(_0498_));
 sky130_fd_sc_hd__and4_1 _2884_ (.A(\d6.saw_temp[4] ),
    .B(\d6.saw_temp[3] ),
    .C(\d6.saw_temp[0] ),
    .D(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__and2_1 _2885_ (.A(\d6.saw_temp[7] ),
    .B(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__o21ai_2 _2886_ (.A1(_0497_),
    .A2(_0500_),
    .B1(\d6.saw_temp[0] ),
    .Y(_0501_));
 sky130_fd_sc_hd__o21a_1 _2887_ (.A1(net206),
    .A2(_0497_),
    .B1(_0501_),
    .X(_0048_));
 sky130_fd_sc_hd__xnor2_1 _2888_ (.A(net139),
    .B(_0501_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _2889_ (.A(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__and3_1 _2890_ (.A(\d6.saw_temp[2] ),
    .B(\d6.saw_temp[1] ),
    .C(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__a21oi_1 _2891_ (.A1(\d6.saw_temp[1] ),
    .A2(_0502_),
    .B1(net171),
    .Y(_0504_));
 sky130_fd_sc_hd__nor2_1 _2892_ (.A(_0503_),
    .B(_0504_),
    .Y(_0050_));
 sky130_fd_sc_hd__xor2_1 _2893_ (.A(net146),
    .B(_0503_),
    .X(_0051_));
 sky130_fd_sc_hd__and3_1 _2894_ (.A(\d6.saw_temp[4] ),
    .B(\d6.saw_temp[3] ),
    .C(_0503_),
    .X(_0505_));
 sky130_fd_sc_hd__a21oi_1 _2895_ (.A1(\d6.saw_temp[3] ),
    .A2(_0503_),
    .B1(net168),
    .Y(_0506_));
 sky130_fd_sc_hd__nor2_1 _2896_ (.A(_0505_),
    .B(_0506_),
    .Y(_0052_));
 sky130_fd_sc_hd__xor2_1 _2897_ (.A(net140),
    .B(_0505_),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _2898_ (.A(\d6.saw_temp[5] ),
    .B(_0505_),
    .X(_0507_));
 sky130_fd_sc_hd__xor2_1 _2899_ (.A(net112),
    .B(_0507_),
    .X(_0054_));
 sky130_fd_sc_hd__a21oi_1 _2900_ (.A1(_0497_),
    .A2(_0499_),
    .B1(net202),
    .Y(_0508_));
 sky130_fd_sc_hd__nor2_1 _2901_ (.A(_0500_),
    .B(_0508_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _2902_ (.A(\d7.count[6] ),
    .Y(_0509_));
 sky130_fd_sc_hd__o221a_1 _2903_ (.A1(\d7.count[6] ),
    .A2(_1733_),
    .B1(_1950_),
    .B2(\d7.count[3] ),
    .C1(_1948_),
    .X(_0510_));
 sky130_fd_sc_hd__o211a_1 _2904_ (.A1(_0509_),
    .A2(_1726_),
    .B1(_1949_),
    .C1(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__a221o_1 _2905_ (.A1(\d7.count[1] ),
    .A2(_1723_),
    .B1(_1777_),
    .B2(\d7.count[0] ),
    .C1(_1955_),
    .X(_0512_));
 sky130_fd_sc_hd__a2111oi_1 _2906_ (.A1(\d7.count[8] ),
    .A2(_1805_),
    .B1(_1957_),
    .C1(_0512_),
    .D1(\d7.count[9] ),
    .Y(_0513_));
 sky130_fd_sc_hd__and3_2 _2907_ (.A(_1947_),
    .B(_0511_),
    .C(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__and4_1 _2908_ (.A(\d7.saw_temp[6] ),
    .B(\d7.saw_temp[5] ),
    .C(\d7.saw_temp[2] ),
    .D(\d7.saw_temp[1] ),
    .X(_0515_));
 sky130_fd_sc_hd__and4_1 _2909_ (.A(\d7.saw_temp[4] ),
    .B(\d7.saw_temp[3] ),
    .C(\d7.saw_temp[0] ),
    .D(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__and2_1 _2910_ (.A(\d7.saw_temp[7] ),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__o21ai_1 _2911_ (.A1(_0514_),
    .A2(_0517_),
    .B1(\d7.saw_temp[0] ),
    .Y(_0518_));
 sky130_fd_sc_hd__o21a_1 _2912_ (.A1(net189),
    .A2(_0514_),
    .B1(_0518_),
    .X(_0056_));
 sky130_fd_sc_hd__inv_2 _2913_ (.A(\d7.saw_temp[1] ),
    .Y(_0519_));
 sky130_fd_sc_hd__nor2_1 _2914_ (.A(_0519_),
    .B(_0518_),
    .Y(_0520_));
 sky130_fd_sc_hd__and2_1 _2915_ (.A(_0519_),
    .B(_0518_),
    .X(_0521_));
 sky130_fd_sc_hd__nor2_1 _2916_ (.A(_0520_),
    .B(_0521_),
    .Y(_0057_));
 sky130_fd_sc_hd__o2111a_1 _2917_ (.A1(_0514_),
    .A2(_0517_),
    .B1(\d7.saw_temp[2] ),
    .C1(\d7.saw_temp[1] ),
    .D1(\d7.saw_temp[0] ),
    .X(_0522_));
 sky130_fd_sc_hd__o21ba_1 _2918_ (.A1(net180),
    .A2(_0520_),
    .B1_N(_0522_),
    .X(_0058_));
 sky130_fd_sc_hd__nand2_1 _2919_ (.A(\d7.saw_temp[3] ),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__or2_1 _2920_ (.A(\d7.saw_temp[3] ),
    .B(_0522_),
    .X(_0524_));
 sky130_fd_sc_hd__and2_1 _2921_ (.A(_0523_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _2922_ (.A(_0525_),
    .X(_0059_));
 sky130_fd_sc_hd__xnor2_1 _2923_ (.A(net173),
    .B(_0523_),
    .Y(_0060_));
 sky130_fd_sc_hd__and4_1 _2924_ (.A(\d7.saw_temp[5] ),
    .B(\d7.saw_temp[4] ),
    .C(\d7.saw_temp[3] ),
    .D(_0522_),
    .X(_0526_));
 sky130_fd_sc_hd__a31oi_1 _2925_ (.A1(\d7.saw_temp[4] ),
    .A2(\d7.saw_temp[3] ),
    .A3(_0522_),
    .B1(net155),
    .Y(_0527_));
 sky130_fd_sc_hd__nor2_1 _2926_ (.A(_0526_),
    .B(_0527_),
    .Y(_0061_));
 sky130_fd_sc_hd__xor2_1 _2927_ (.A(net94),
    .B(_0526_),
    .X(_0062_));
 sky130_fd_sc_hd__a21oi_1 _2928_ (.A1(_0514_),
    .A2(_0516_),
    .B1(net192),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_1 _2929_ (.A(_0517_),
    .B(_0528_),
    .Y(_0063_));
 sky130_fd_sc_hd__and4_1 _2930_ (.A(\d8.saw_temp[5] ),
    .B(\d8.saw_temp[4] ),
    .C(\d8.saw_temp[1] ),
    .D(\d8.saw_temp[2] ),
    .X(_0529_));
 sky130_fd_sc_hd__and4_1 _2931_ (.A(\d8.saw_temp[6] ),
    .B(\d8.saw_temp[0] ),
    .C(\d8.saw_temp[3] ),
    .D(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__and2_1 _2932_ (.A(\d8.saw_temp[7] ),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__a211o_1 _2933_ (.A1(\d8.count[8] ),
    .A2(_1715_),
    .B1(_1980_),
    .C1(\d8.count[9] ),
    .X(_0532_));
 sky130_fd_sc_hd__a21oi_1 _2934_ (.A1(\d8.count[6] ),
    .A2(_1733_),
    .B1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__a22o_1 _2935_ (.A1(\d8.count[3] ),
    .A2(_1718_),
    .B1(_1723_),
    .B2(\d8.count[2] ),
    .X(_0534_));
 sky130_fd_sc_hd__a2bb2o_1 _2936_ (.A1_N(\d8.count[3] ),
    .A2_N(_1718_),
    .B1(_1777_),
    .B2(\d8.count[1] ),
    .X(_0535_));
 sky130_fd_sc_hd__nor2_1 _2937_ (.A(_0534_),
    .B(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_2 _2938_ (.A(\d8.count[0] ),
    .Y(_0537_));
 sky130_fd_sc_hd__o2111a_1 _2939_ (.A1(_1735_),
    .A2(\d8.count[5] ),
    .B1(_1988_),
    .C1(_1986_),
    .D1(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__o2111a_1 _2940_ (.A1(\d8.count[8] ),
    .A2(_1805_),
    .B1(_1981_),
    .C1(_0536_),
    .D1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__o2111a_2 _2941_ (.A1(\d8.count[6] ),
    .A2(_1733_),
    .B1(_1983_),
    .C1(_0533_),
    .D1(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__o21a_1 _2942_ (.A1(_0531_),
    .A2(_0540_),
    .B1(\d8.saw_temp[0] ),
    .X(_0541_));
 sky130_fd_sc_hd__nor3_1 _2943_ (.A(\d8.saw_temp[0] ),
    .B(_0531_),
    .C(_0540_),
    .Y(_0542_));
 sky130_fd_sc_hd__nor2_1 _2944_ (.A(_0541_),
    .B(_0542_),
    .Y(_0064_));
 sky130_fd_sc_hd__xor2_1 _2945_ (.A(net129),
    .B(_0541_),
    .X(_0065_));
 sky130_fd_sc_hd__and3_1 _2946_ (.A(\d8.saw_temp[1] ),
    .B(\d8.saw_temp[2] ),
    .C(_0541_),
    .X(_0543_));
 sky130_fd_sc_hd__a21oi_1 _2947_ (.A1(\d8.saw_temp[1] ),
    .A2(_0541_),
    .B1(net216),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_1 _2948_ (.A(_0543_),
    .B(net217),
    .Y(_0066_));
 sky130_fd_sc_hd__xor2_1 _2949_ (.A(net164),
    .B(_0543_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _2950_ (.A(\d8.saw_temp[4] ),
    .B(\d8.saw_temp[3] ),
    .C(_0543_),
    .X(_0545_));
 sky130_fd_sc_hd__a21oi_1 _2951_ (.A1(\d8.saw_temp[3] ),
    .A2(_0543_),
    .B1(net167),
    .Y(_0546_));
 sky130_fd_sc_hd__nor2_1 _2952_ (.A(_0545_),
    .B(_0546_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand2_1 _2953_ (.A(\d8.saw_temp[5] ),
    .B(_0545_),
    .Y(_0547_));
 sky130_fd_sc_hd__or2_1 _2954_ (.A(\d8.saw_temp[5] ),
    .B(_0545_),
    .X(_0548_));
 sky130_fd_sc_hd__and2_1 _2955_ (.A(_0547_),
    .B(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(_0549_),
    .X(_0069_));
 sky130_fd_sc_hd__xnor2_1 _2957_ (.A(net133),
    .B(_0547_),
    .Y(_0070_));
 sky130_fd_sc_hd__a21oi_1 _2958_ (.A1(_0530_),
    .A2(_0540_),
    .B1(\d8.saw_temp[7] ),
    .Y(_0550_));
 sky130_fd_sc_hd__nor2_1 _2959_ (.A(_0531_),
    .B(_0550_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _2960_ (.A(\d1.saw_temp[0] ),
    .Y(_0551_));
 sky130_fd_sc_hd__a2bb2o_1 _2961_ (.A1_N(\d1.count[5] ),
    .A2_N(_1720_),
    .B1(_1723_),
    .B2(\d1.count[7] ),
    .X(_0552_));
 sky130_fd_sc_hd__a221o_1 _2962_ (.A1(_1735_),
    .A2(\d1.count[1] ),
    .B1(_1744_),
    .B2(_1724_),
    .C1(_1738_),
    .X(_0553_));
 sky130_fd_sc_hd__a211o_1 _2963_ (.A1(\d1.count[0] ),
    .A2(_1777_),
    .B1(_0553_),
    .C1(_1719_),
    .X(_0554_));
 sky130_fd_sc_hd__o21ba_1 _2964_ (.A1(\d1.count[6] ),
    .A2(_1726_),
    .B1_N(_1728_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _2965_ (.A(\d1.count[6] ),
    .B(_1726_),
    .Y(_0556_));
 sky130_fd_sc_hd__o221a_1 _2966_ (.A1(\d1.count[8] ),
    .A2(_1720_),
    .B1(_1723_),
    .B2(\d1.count[7] ),
    .C1(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__o211ai_1 _2967_ (.A1(_1945_),
    .A2(_1730_),
    .B1(_0555_),
    .C1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__or4_2 _2968_ (.A(_1737_),
    .B(_0552_),
    .C(_0554_),
    .D(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__inv_2 _2969_ (.A(\d1.saw_temp[7] ),
    .Y(_0560_));
 sky130_fd_sc_hd__and4_1 _2970_ (.A(\d1.saw_temp[6] ),
    .B(\d1.saw_temp[5] ),
    .C(\d1.saw_temp[2] ),
    .D(\d1.saw_temp[1] ),
    .X(_0561_));
 sky130_fd_sc_hd__nand4_1 _2971_ (.A(\d1.saw_temp[4] ),
    .B(\d1.saw_temp[3] ),
    .C(\d1.saw_temp[0] ),
    .D(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__or2_1 _2972_ (.A(_0560_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a21oi_2 _2973_ (.A1(_0563_),
    .A2(_0559_),
    .B1(_0551_),
    .Y(_0564_));
 sky130_fd_sc_hd__a21oi_1 _2974_ (.A1(_0551_),
    .A2(_0559_),
    .B1(_0564_),
    .Y(_0072_));
 sky130_fd_sc_hd__xor2_1 _2975_ (.A(net177),
    .B(_0564_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_1 _2976_ (.A(\d1.saw_temp[2] ),
    .B(\d1.saw_temp[1] ),
    .C(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__a21oi_1 _2977_ (.A1(\d1.saw_temp[1] ),
    .A2(_0564_),
    .B1(net178),
    .Y(_0566_));
 sky130_fd_sc_hd__nor2_1 _2978_ (.A(_0565_),
    .B(_0566_),
    .Y(_0074_));
 sky130_fd_sc_hd__xor2_1 _2979_ (.A(net169),
    .B(_0565_),
    .X(_0075_));
 sky130_fd_sc_hd__and3_1 _2980_ (.A(\d1.saw_temp[4] ),
    .B(\d1.saw_temp[3] ),
    .C(_0565_),
    .X(_0567_));
 sky130_fd_sc_hd__a21oi_1 _2981_ (.A1(\d1.saw_temp[3] ),
    .A2(_0565_),
    .B1(net172),
    .Y(_0568_));
 sky130_fd_sc_hd__nor2_1 _2982_ (.A(_0567_),
    .B(_0568_),
    .Y(_0076_));
 sky130_fd_sc_hd__nand2_1 _2983_ (.A(\d1.saw_temp[5] ),
    .B(_0567_),
    .Y(_0569_));
 sky130_fd_sc_hd__or2_1 _2984_ (.A(\d1.saw_temp[5] ),
    .B(_0567_),
    .X(_0570_));
 sky130_fd_sc_hd__and2_1 _2985_ (.A(_0569_),
    .B(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _2986_ (.A(_0571_),
    .X(_0077_));
 sky130_fd_sc_hd__xnor2_1 _2987_ (.A(net108),
    .B(_0569_),
    .Y(_0078_));
 sky130_fd_sc_hd__nor2_1 _2988_ (.A(_0562_),
    .B(_0559_),
    .Y(_0572_));
 sky130_fd_sc_hd__o21a_1 _2989_ (.A1(\d1.saw_temp[7] ),
    .A2(_0572_),
    .B1(_0563_),
    .X(_0079_));
 sky130_fd_sc_hd__and4_1 _2990_ (.A(\d10.saw_temp[6] ),
    .B(\d10.saw_temp[5] ),
    .C(\d10.saw_temp[2] ),
    .D(\d10.saw_temp[1] ),
    .X(_0573_));
 sky130_fd_sc_hd__and4_1 _2991_ (.A(\d10.saw_temp[4] ),
    .B(\d10.saw_temp[3] ),
    .C(\d10.saw_temp[0] ),
    .D(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__and2_1 _2992_ (.A(\d10.saw_temp[7] ),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _2993_ (.A1(\d10.count[7] ),
    .A2(_1720_),
    .B1(_1777_),
    .B2(\d10.count[2] ),
    .X(_0576_));
 sky130_fd_sc_hd__nor2_1 _2994_ (.A(_1872_),
    .B(_0163_),
    .Y(_0577_));
 sky130_fd_sc_hd__a211o_1 _2995_ (.A1(_1735_),
    .A2(\d10.count[3] ),
    .B1(_0162_),
    .C1(_0173_),
    .X(_0578_));
 sky130_fd_sc_hd__or4b_1 _2996_ (.A(_0577_),
    .B(_0171_),
    .C(_0578_),
    .D_N(_0161_),
    .X(_0579_));
 sky130_fd_sc_hd__a2111oi_1 _2997_ (.A1(\d10.count[5] ),
    .A2(_1729_),
    .B1(_0168_),
    .C1(_0576_),
    .D1(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__o21a_1 _2998_ (.A1(_0575_),
    .A2(net18),
    .B1(\d10.saw_temp[0] ),
    .X(_0581_));
 sky130_fd_sc_hd__nor3_1 _2999_ (.A(net233),
    .B(_0575_),
    .C(net18),
    .Y(_0582_));
 sky130_fd_sc_hd__nor2_1 _3000_ (.A(_0581_),
    .B(_0582_),
    .Y(_0080_));
 sky130_fd_sc_hd__xor2_1 _3001_ (.A(net124),
    .B(_0581_),
    .X(_0081_));
 sky130_fd_sc_hd__and3_1 _3002_ (.A(\d10.saw_temp[2] ),
    .B(\d10.saw_temp[1] ),
    .C(_0581_),
    .X(_0583_));
 sky130_fd_sc_hd__a21oi_1 _3003_ (.A1(\d10.saw_temp[1] ),
    .A2(_0581_),
    .B1(net198),
    .Y(_0584_));
 sky130_fd_sc_hd__nor2_1 _3004_ (.A(_0583_),
    .B(net199),
    .Y(_0082_));
 sky130_fd_sc_hd__xor2_1 _3005_ (.A(net120),
    .B(_0583_),
    .X(_0083_));
 sky130_fd_sc_hd__and3_1 _3006_ (.A(\d10.saw_temp[4] ),
    .B(\d10.saw_temp[3] ),
    .C(_0583_),
    .X(_0585_));
 sky130_fd_sc_hd__a21oi_1 _3007_ (.A1(net120),
    .A2(_0583_),
    .B1(net144),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_1 _3008_ (.A(_0585_),
    .B(_0586_),
    .Y(_0084_));
 sky130_fd_sc_hd__xor2_1 _3009_ (.A(net142),
    .B(_0585_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _3010_ (.A(net252),
    .B(_0585_),
    .X(_0587_));
 sky130_fd_sc_hd__xor2_1 _3011_ (.A(net117),
    .B(_0587_),
    .X(_0086_));
 sky130_fd_sc_hd__a21oi_1 _3012_ (.A1(_0574_),
    .A2(net18),
    .B1(net183),
    .Y(_0588_));
 sky130_fd_sc_hd__nor2_1 _3013_ (.A(_0575_),
    .B(_0588_),
    .Y(_0087_));
 sky130_fd_sc_hd__and4b_1 _3014_ (.A_N(_0202_),
    .B(_0194_),
    .C(_0206_),
    .D(_0193_),
    .X(_0589_));
 sky130_fd_sc_hd__a211o_1 _3015_ (.A1(\d11.count[1] ),
    .A2(_1732_),
    .B1(_0201_),
    .C1(\d11.count[0] ),
    .X(_0590_));
 sky130_fd_sc_hd__a21oi_1 _3016_ (.A1(\d11.count[7] ),
    .A2(_1718_),
    .B1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__o21a_1 _3017_ (.A1(\d11.count[8] ),
    .A2(_1715_),
    .B1(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__and4_1 _3018_ (.A(\d11.saw_temp[6] ),
    .B(\d11.saw_temp[5] ),
    .C(\d11.saw_temp[2] ),
    .D(\d11.saw_temp[1] ),
    .X(_0593_));
 sky130_fd_sc_hd__and4_1 _3019_ (.A(\d11.saw_temp[4] ),
    .B(\d11.saw_temp[3] ),
    .C(\d11.saw_temp[0] ),
    .D(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__and2_1 _3020_ (.A(\d11.saw_temp[7] ),
    .B(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__a31o_2 _3021_ (.A1(_0198_),
    .A2(_0589_),
    .A3(_0592_),
    .B1(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__nor2_1 _3022_ (.A(net247),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _3023_ (.A(\d11.saw_temp[0] ),
    .B(_0596_),
    .Y(_0598_));
 sky130_fd_sc_hd__inv_2 _3024_ (.A(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__nor2_1 _3025_ (.A(_0597_),
    .B(_0599_),
    .Y(_0088_));
 sky130_fd_sc_hd__xnor2_1 _3026_ (.A(net135),
    .B(_0598_),
    .Y(_0089_));
 sky130_fd_sc_hd__a21oi_1 _3027_ (.A1(\d11.saw_temp[1] ),
    .A2(_0599_),
    .B1(\d11.saw_temp[2] ),
    .Y(_0600_));
 sky130_fd_sc_hd__and3_1 _3028_ (.A(\d11.saw_temp[2] ),
    .B(\d11.saw_temp[1] ),
    .C(_0599_),
    .X(_0601_));
 sky130_fd_sc_hd__nor2_1 _3029_ (.A(_0600_),
    .B(_0601_),
    .Y(_0090_));
 sky130_fd_sc_hd__xor2_1 _3030_ (.A(net136),
    .B(_0601_),
    .X(_0091_));
 sky130_fd_sc_hd__a21oi_1 _3031_ (.A1(\d11.saw_temp[3] ),
    .A2(_0601_),
    .B1(net231),
    .Y(_0602_));
 sky130_fd_sc_hd__and3_1 _3032_ (.A(\d11.saw_temp[4] ),
    .B(\d11.saw_temp[3] ),
    .C(_0601_),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_1 _3033_ (.A(_0602_),
    .B(_0603_),
    .Y(_0092_));
 sky130_fd_sc_hd__or2_1 _3034_ (.A(\d11.saw_temp[5] ),
    .B(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_1 _3035_ (.A(\d11.saw_temp[5] ),
    .B(_0603_),
    .Y(_0605_));
 sky130_fd_sc_hd__and2_1 _3036_ (.A(_0604_),
    .B(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_1 _3037_ (.A(_0606_),
    .X(_0093_));
 sky130_fd_sc_hd__xnor2_1 _3038_ (.A(net99),
    .B(_0605_),
    .Y(_0094_));
 sky130_fd_sc_hd__a41o_1 _3039_ (.A1(_0198_),
    .A2(_0594_),
    .A3(_0589_),
    .A4(_0592_),
    .B1(\d11.saw_temp[7] ),
    .X(_0607_));
 sky130_fd_sc_hd__and2b_1 _3040_ (.A_N(_0595_),
    .B(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_1 _3041_ (.A(_0608_),
    .X(_0095_));
 sky130_fd_sc_hd__or2b_1 _3042_ (.A(_0306_),
    .B_N(_0300_),
    .X(_0609_));
 sky130_fd_sc_hd__nor2b_2 _3043_ (.A(_0300_),
    .B_N(_0306_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand2_2 _3044_ (.A(\d2.saw_temp[7] ),
    .B(_0329_),
    .Y(_0611_));
 sky130_fd_sc_hd__o31a_1 _3045_ (.A1(\d2.saw_temp[5] ),
    .A2(\d2.saw_temp[4] ),
    .A3(\d2.saw_temp[3] ),
    .B1(net7),
    .X(_0612_));
 sky130_fd_sc_hd__nand2_1 _3046_ (.A(\d2.saw_temp[0] ),
    .B(_0329_),
    .Y(_0613_));
 sky130_fd_sc_hd__o21ai_1 _3047_ (.A1(\d2.saw_temp[2] ),
    .A2(\d2.saw_temp[1] ),
    .B1(_0329_),
    .Y(_0614_));
 sky130_fd_sc_hd__and4bb_2 _3048_ (.A_N(\d2.saw_temp[6] ),
    .B_N(_0612_),
    .C(_0613_),
    .D(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__or3_1 _3049_ (.A(_0610_),
    .B(_0611_),
    .C(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__or2b_1 _3050_ (.A(_0300_),
    .B_N(_0306_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_4 _3051_ (.A(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__or2_1 _3052_ (.A(_0618_),
    .B(_0613_),
    .X(_0619_));
 sky130_fd_sc_hd__a31oi_4 _3053_ (.A1(\d2.saw_temp[7] ),
    .A2(_0329_),
    .A3(_0300_),
    .B1(_0306_),
    .Y(_0620_));
 sky130_fd_sc_hd__a31o_1 _3054_ (.A1(_0609_),
    .A2(_0616_),
    .A3(_0619_),
    .B1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_8 _3055_ (.A(_0609_),
    .X(_0622_));
 sky130_fd_sc_hd__nand2_2 _3056_ (.A(\d1.saw_temp[7] ),
    .B(_0330_),
    .Y(_0623_));
 sky130_fd_sc_hd__o31a_1 _3057_ (.A1(\d1.saw_temp[5] ),
    .A2(\d1.saw_temp[4] ),
    .A3(\d1.saw_temp[3] ),
    .B1(_0330_),
    .X(_0624_));
 sky130_fd_sc_hd__nand2_1 _3058_ (.A(\d1.saw_temp[0] ),
    .B(_0330_),
    .Y(_0625_));
 sky130_fd_sc_hd__o21ai_1 _3059_ (.A1(\d1.saw_temp[2] ),
    .A2(\d1.saw_temp[1] ),
    .B1(_0330_),
    .Y(_0626_));
 sky130_fd_sc_hd__and4bb_2 _3060_ (.A_N(\d1.saw_temp[6] ),
    .B_N(_0624_),
    .C(_0625_),
    .D(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__or3_1 _3061_ (.A(_0610_),
    .B(_0623_),
    .C(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__or2_1 _3062_ (.A(_0618_),
    .B(_0625_),
    .X(_0629_));
 sky130_fd_sc_hd__a31oi_4 _3063_ (.A1(\d1.saw_temp[7] ),
    .A2(_0300_),
    .A3(_0330_),
    .B1(_0306_),
    .Y(_0630_));
 sky130_fd_sc_hd__a31o_1 _3064_ (.A1(_0622_),
    .A2(_0628_),
    .A3(_0629_),
    .B1(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__xor2_2 _3065_ (.A(_0621_),
    .B(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__a31o_2 _3066_ (.A1(\d13.saw_temp[7] ),
    .A2(_0301_),
    .A3(_0344_),
    .B1(_0307_),
    .X(_0633_));
 sky130_fd_sc_hd__buf_8 _3067_ (.A(_0618_),
    .X(_0634_));
 sky130_fd_sc_hd__and2_2 _3068_ (.A(\d13.saw_temp[7] ),
    .B(_0344_),
    .X(_0635_));
 sky130_fd_sc_hd__o31a_1 _3069_ (.A1(\d13.saw_temp[4] ),
    .A2(\d13.saw_temp[2] ),
    .A3(\d13.saw_temp[1] ),
    .B1(_0344_),
    .X(_0636_));
 sky130_fd_sc_hd__o21a_1 _3070_ (.A1(\d13.saw_temp[3] ),
    .A2(\d13.saw_temp[0] ),
    .B1(_0344_),
    .X(_0637_));
 sky130_fd_sc_hd__nand2_1 _3071_ (.A(\d13.saw_temp[5] ),
    .B(_0344_),
    .Y(_0638_));
 sky130_fd_sc_hd__or4b_2 _3072_ (.A(\d13.saw_temp[6] ),
    .B(_0636_),
    .C(_0637_),
    .D_N(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_8 _3073_ (.A(_0610_),
    .X(_0640_));
 sky130_fd_sc_hd__a31o_1 _3074_ (.A1(\d13.saw_temp[0] ),
    .A2(_0344_),
    .A3(_0640_),
    .B1(_0309_),
    .X(_0641_));
 sky130_fd_sc_hd__a31o_1 _3075_ (.A1(_0634_),
    .A2(_0635_),
    .A3(_0639_),
    .B1(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nand2_1 _3076_ (.A(_0633_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__xor2_1 _3077_ (.A(_0632_),
    .B(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__a31o_2 _3078_ (.A1(\d12.saw_temp[7] ),
    .A2(_0301_),
    .A3(_0340_),
    .B1(_0307_),
    .X(_0645_));
 sky130_fd_sc_hd__buf_8 _3079_ (.A(_0634_),
    .X(_0646_));
 sky130_fd_sc_hd__and2_2 _3080_ (.A(\d12.saw_temp[7] ),
    .B(_0340_),
    .X(_0647_));
 sky130_fd_sc_hd__o31a_1 _3081_ (.A1(\d12.saw_temp[4] ),
    .A2(\d12.saw_temp[2] ),
    .A3(\d12.saw_temp[1] ),
    .B1(_0340_),
    .X(_0648_));
 sky130_fd_sc_hd__o21a_1 _3082_ (.A1(\d12.saw_temp[3] ),
    .A2(\d12.saw_temp[0] ),
    .B1(_0340_),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_1 _3083_ (.A(\d12.saw_temp[5] ),
    .B(_0340_),
    .Y(_0650_));
 sky130_fd_sc_hd__or4b_2 _3084_ (.A(\d12.saw_temp[6] ),
    .B(_0648_),
    .C(_0649_),
    .D_N(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__a31o_1 _3085_ (.A1(\d12.saw_temp[0] ),
    .A2(_0340_),
    .A3(_0640_),
    .B1(_0309_),
    .X(_0652_));
 sky130_fd_sc_hd__a31o_1 _3086_ (.A1(_0646_),
    .A2(_0647_),
    .A3(_0651_),
    .B1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__nand2_1 _3087_ (.A(_0645_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__nor2_1 _3088_ (.A(_0644_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__and2_1 _3089_ (.A(_0644_),
    .B(_0654_),
    .X(_0656_));
 sky130_fd_sc_hd__or2_1 _3090_ (.A(_0655_),
    .B(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__and2_2 _3091_ (.A(\d11.saw_temp[7] ),
    .B(_0334_),
    .X(_0658_));
 sky130_fd_sc_hd__a21oi_4 _3092_ (.A1(_0301_),
    .A2(_0658_),
    .B1(_0307_),
    .Y(_0659_));
 sky130_fd_sc_hd__o31a_1 _3093_ (.A1(\d11.saw_temp[4] ),
    .A2(\d11.saw_temp[2] ),
    .A3(\d11.saw_temp[1] ),
    .B1(_0334_),
    .X(_0660_));
 sky130_fd_sc_hd__o21a_1 _3094_ (.A1(\d11.saw_temp[3] ),
    .A2(\d11.saw_temp[0] ),
    .B1(_0334_),
    .X(_0661_));
 sky130_fd_sc_hd__nand2_1 _3095_ (.A(\d11.saw_temp[5] ),
    .B(_0334_),
    .Y(_0662_));
 sky130_fd_sc_hd__or4b_1 _3096_ (.A(\d11.saw_temp[6] ),
    .B(_0660_),
    .C(_0661_),
    .D_N(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__nand2_2 _3097_ (.A(_0658_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__a31o_1 _3098_ (.A1(\d11.saw_temp[0] ),
    .A2(_0334_),
    .A3(_0640_),
    .B1(_0309_),
    .X(_0665_));
 sky130_fd_sc_hd__o21ba_1 _3099_ (.A1(_0640_),
    .A2(_0664_),
    .B1_N(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__or2_1 _3100_ (.A(_0659_),
    .B(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__and2_2 _3101_ (.A(\d10.saw_temp[7] ),
    .B(_0336_),
    .X(_0668_));
 sky130_fd_sc_hd__a21oi_4 _3102_ (.A1(_0301_),
    .A2(_0668_),
    .B1(_0307_),
    .Y(_0669_));
 sky130_fd_sc_hd__o31a_1 _3103_ (.A1(\d10.saw_temp[4] ),
    .A2(\d10.saw_temp[2] ),
    .A3(\d10.saw_temp[1] ),
    .B1(_0336_),
    .X(_0670_));
 sky130_fd_sc_hd__o21a_1 _3104_ (.A1(\d10.saw_temp[3] ),
    .A2(\d10.saw_temp[0] ),
    .B1(_0336_),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _3105_ (.A(\d10.saw_temp[5] ),
    .B(_0336_),
    .Y(_0672_));
 sky130_fd_sc_hd__or4b_1 _3106_ (.A(\d10.saw_temp[6] ),
    .B(_0670_),
    .C(_0671_),
    .D_N(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_2 _3107_ (.A(_0668_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__a31o_1 _3108_ (.A1(\d10.saw_temp[0] ),
    .A2(_0336_),
    .A3(_0640_),
    .B1(_0309_),
    .X(_0675_));
 sky130_fd_sc_hd__o21ba_1 _3109_ (.A1(_0640_),
    .A2(_0674_),
    .B1_N(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__or2_1 _3110_ (.A(_0669_),
    .B(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__xor2_1 _3111_ (.A(_0667_),
    .B(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__inv_2 _3112_ (.A(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__and2_2 _3113_ (.A(\d9.saw_temp[7] ),
    .B(_0335_),
    .X(_0680_));
 sky130_fd_sc_hd__a21oi_4 _3114_ (.A1(_0301_),
    .A2(_0680_),
    .B1(_0307_),
    .Y(_0681_));
 sky130_fd_sc_hd__clkbuf_8 _3115_ (.A(_0640_),
    .X(_0682_));
 sky130_fd_sc_hd__buf_6 _3116_ (.A(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__o31a_1 _3117_ (.A1(\d9.saw_temp[4] ),
    .A2(\d9.saw_temp[1] ),
    .A3(\d9.saw_temp[2] ),
    .B1(_0335_),
    .X(_0684_));
 sky130_fd_sc_hd__o21a_1 _3118_ (.A1(\d9.saw_temp[0] ),
    .A2(\d9.saw_temp[3] ),
    .B1(_0335_),
    .X(_0685_));
 sky130_fd_sc_hd__nand2_1 _3119_ (.A(\d9.saw_temp[5] ),
    .B(_0335_),
    .Y(_0686_));
 sky130_fd_sc_hd__or4b_1 _3120_ (.A(\d9.saw_temp[6] ),
    .B(_0684_),
    .C(_0685_),
    .D_N(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__nand2_2 _3121_ (.A(_0680_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__a31o_1 _3122_ (.A1(\d9.saw_temp[0] ),
    .A2(_0335_),
    .A3(_0682_),
    .B1(_0309_),
    .X(_0689_));
 sky130_fd_sc_hd__o21ba_1 _3123_ (.A1(_0683_),
    .A2(_0688_),
    .B1_N(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__or2_1 _3124_ (.A(_0681_),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__nor2_1 _3125_ (.A(_0679_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__and2_1 _3126_ (.A(_0679_),
    .B(_0691_),
    .X(_0693_));
 sky130_fd_sc_hd__or2_1 _3127_ (.A(_0692_),
    .B(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__nor2_1 _3128_ (.A(_0657_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__and2_1 _3129_ (.A(_0657_),
    .B(_0694_),
    .X(_0696_));
 sky130_fd_sc_hd__and2_1 _3130_ (.A(\d8.saw_temp[7] ),
    .B(_0337_),
    .X(_0697_));
 sky130_fd_sc_hd__o31a_1 _3131_ (.A1(\d8.saw_temp[4] ),
    .A2(\d8.saw_temp[1] ),
    .A3(\d8.saw_temp[2] ),
    .B1(_0337_),
    .X(_0698_));
 sky130_fd_sc_hd__o21a_1 _3132_ (.A1(\d8.saw_temp[0] ),
    .A2(\d8.saw_temp[3] ),
    .B1(_0337_),
    .X(_0699_));
 sky130_fd_sc_hd__nand2_1 _3133_ (.A(\d8.saw_temp[5] ),
    .B(_0337_),
    .Y(_0700_));
 sky130_fd_sc_hd__or4b_2 _3134_ (.A(\d8.saw_temp[6] ),
    .B(_0698_),
    .C(_0699_),
    .D_N(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_2 _3135_ (.A(_0697_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__nor2_1 _3136_ (.A(_0683_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__a31o_1 _3137_ (.A1(\d8.saw_temp[0] ),
    .A2(_0337_),
    .A3(_0682_),
    .B1(_0310_),
    .X(_0704_));
 sky130_fd_sc_hd__a31o_2 _3138_ (.A1(\d8.saw_temp[7] ),
    .A2(_0301_),
    .A3(_0337_),
    .B1(_0307_),
    .X(_0705_));
 sky130_fd_sc_hd__o21ai_2 _3139_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__and2_2 _3140_ (.A(\d7.saw_temp[7] ),
    .B(net12),
    .X(_0707_));
 sky130_fd_sc_hd__a21oi_4 _3141_ (.A1(_0301_),
    .A2(_0707_),
    .B1(_0307_),
    .Y(_0708_));
 sky130_fd_sc_hd__o31a_1 _3142_ (.A1(\d7.saw_temp[4] ),
    .A2(\d7.saw_temp[2] ),
    .A3(\d7.saw_temp[1] ),
    .B1(net12),
    .X(_0709_));
 sky130_fd_sc_hd__o21a_1 _3143_ (.A1(\d7.saw_temp[3] ),
    .A2(\d7.saw_temp[0] ),
    .B1(net12),
    .X(_0710_));
 sky130_fd_sc_hd__nand2_1 _3144_ (.A(\d7.saw_temp[5] ),
    .B(net12),
    .Y(_0711_));
 sky130_fd_sc_hd__or4b_1 _3145_ (.A(\d7.saw_temp[6] ),
    .B(_0709_),
    .C(_0710_),
    .D_N(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_2 _3146_ (.A(_0707_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__a31o_1 _3147_ (.A1(\d7.saw_temp[0] ),
    .A2(net12),
    .A3(_0640_),
    .B1(_0309_),
    .X(_0714_));
 sky130_fd_sc_hd__o21ba_1 _3148_ (.A1(_0682_),
    .A2(_0713_),
    .B1_N(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__or2_1 _3149_ (.A(_0708_),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__nor2_1 _3150_ (.A(_0706_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__and2_1 _3151_ (.A(_0706_),
    .B(_0716_),
    .X(_0718_));
 sky130_fd_sc_hd__nor2_1 _3152_ (.A(_0717_),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__inv_2 _3153_ (.A(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__and2_2 _3154_ (.A(\d6.saw_temp[7] ),
    .B(_0346_),
    .X(_0721_));
 sky130_fd_sc_hd__a21oi_4 _3155_ (.A1(_0301_),
    .A2(_0721_),
    .B1(_0307_),
    .Y(_0722_));
 sky130_fd_sc_hd__buf_6 _3156_ (.A(_0683_),
    .X(_0723_));
 sky130_fd_sc_hd__o31a_1 _3157_ (.A1(\d6.saw_temp[4] ),
    .A2(\d6.saw_temp[2] ),
    .A3(\d6.saw_temp[1] ),
    .B1(_0346_),
    .X(_0724_));
 sky130_fd_sc_hd__o21a_1 _3158_ (.A1(\d6.saw_temp[3] ),
    .A2(\d6.saw_temp[0] ),
    .B1(_0346_),
    .X(_0725_));
 sky130_fd_sc_hd__nand2_1 _3159_ (.A(\d6.saw_temp[5] ),
    .B(_0346_),
    .Y(_0726_));
 sky130_fd_sc_hd__or4b_1 _3160_ (.A(\d6.saw_temp[6] ),
    .B(_0724_),
    .C(_0725_),
    .D_N(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__nand2_2 _3161_ (.A(_0721_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__a31o_1 _3162_ (.A1(\d6.saw_temp[0] ),
    .A2(_0346_),
    .A3(_0683_),
    .B1(_0310_),
    .X(_0729_));
 sky130_fd_sc_hd__o21ba_1 _3163_ (.A1(_0723_),
    .A2(_0728_),
    .B1_N(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__or2_1 _3164_ (.A(_0722_),
    .B(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__nor2_1 _3165_ (.A(_0720_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__and2_1 _3166_ (.A(_0720_),
    .B(_0731_),
    .X(_0733_));
 sky130_fd_sc_hd__or2_1 _3167_ (.A(_0732_),
    .B(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__or3_2 _3168_ (.A(_0695_),
    .B(_0696_),
    .C(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__inv_2 _3169_ (.A(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__o21a_1 _3170_ (.A1(_0695_),
    .A2(_0696_),
    .B1(_0734_),
    .X(_0737_));
 sky130_fd_sc_hd__buf_6 _3171_ (.A(_0723_),
    .X(_0738_));
 sky130_fd_sc_hd__nand2_1 _3172_ (.A(\d5.saw_temp[7] ),
    .B(_0328_),
    .Y(_0739_));
 sky130_fd_sc_hd__o31a_1 _3173_ (.A1(\d5.saw_temp[4] ),
    .A2(\d5.saw_temp[2] ),
    .A3(\d5.saw_temp[1] ),
    .B1(_0328_),
    .X(_0740_));
 sky130_fd_sc_hd__o21a_1 _3174_ (.A1(\d5.saw_temp[3] ),
    .A2(\d5.saw_temp[0] ),
    .B1(_0328_),
    .X(_0741_));
 sky130_fd_sc_hd__nand2_1 _3175_ (.A(\d5.saw_temp[5] ),
    .B(_0328_),
    .Y(_0742_));
 sky130_fd_sc_hd__or4b_1 _3176_ (.A(\d5.saw_temp[6] ),
    .B(_0740_),
    .C(_0741_),
    .D_N(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__nand2b_2 _3177_ (.A_N(_0739_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__nor2_1 _3178_ (.A(_0738_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__a31o_1 _3179_ (.A1(\d5.saw_temp[0] ),
    .A2(_0328_),
    .A3(_0723_),
    .B1(_0310_),
    .X(_0746_));
 sky130_fd_sc_hd__a31o_2 _3180_ (.A1(\d5.saw_temp[7] ),
    .A2(_0301_),
    .A3(_0328_),
    .B1(_0307_),
    .X(_0747_));
 sky130_fd_sc_hd__o21ai_1 _3181_ (.A1(_0745_),
    .A2(_0746_),
    .B1(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__clkbuf_8 _3182_ (.A(_0622_),
    .X(_0749_));
 sky130_fd_sc_hd__buf_6 _3183_ (.A(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__buf_6 _3184_ (.A(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__nand2_1 _3185_ (.A(\d4.saw_temp[0] ),
    .B(_0347_),
    .Y(_0752_));
 sky130_fd_sc_hd__and2_1 _3186_ (.A(\d4.saw_temp[7] ),
    .B(_0347_),
    .X(_0753_));
 sky130_fd_sc_hd__o31a_1 _3187_ (.A1(\d4.saw_temp[5] ),
    .A2(\d4.saw_temp[4] ),
    .A3(\d4.saw_temp[1] ),
    .B1(_0347_),
    .X(_0754_));
 sky130_fd_sc_hd__nand2_1 _3188_ (.A(\d4.saw_temp[3] ),
    .B(_0347_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _3189_ (.A(\d4.saw_temp[2] ),
    .B(_0347_),
    .Y(_0756_));
 sky130_fd_sc_hd__nand2_1 _3190_ (.A(_0755_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__or4b_1 _3191_ (.A(\d4.saw_temp[6] ),
    .B(_0754_),
    .C(_0757_),
    .D_N(_0752_),
    .X(_0758_));
 sky130_fd_sc_hd__nand2_2 _3192_ (.A(_0753_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__clkbuf_8 _3193_ (.A(_0646_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(_0752_),
    .A1(_0759_),
    .S(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__a31o_2 _3195_ (.A1(\d4.saw_temp[7] ),
    .A2(_0301_),
    .A3(_0347_),
    .B1(_0307_),
    .X(_0762_));
 sky130_fd_sc_hd__a21bo_1 _3196_ (.A1(_0751_),
    .A2(_0761_),
    .B1_N(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__nor2_1 _3197_ (.A(_0748_),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__and2_1 _3198_ (.A(_0748_),
    .B(_0763_),
    .X(_0765_));
 sky130_fd_sc_hd__nor2_1 _3199_ (.A(_0764_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__a31o_2 _3200_ (.A1(\d3.saw_temp[7] ),
    .A2(_0301_),
    .A3(_0348_),
    .B1(_0307_),
    .X(_0767_));
 sky130_fd_sc_hd__and2_1 _3201_ (.A(\d3.saw_temp[7] ),
    .B(_0348_),
    .X(_0768_));
 sky130_fd_sc_hd__o31a_1 _3202_ (.A1(\d3.saw_temp[4] ),
    .A2(\d3.saw_temp[2] ),
    .A3(\d3.saw_temp[1] ),
    .B1(_0348_),
    .X(_0769_));
 sky130_fd_sc_hd__o21a_1 _3203_ (.A1(\d3.saw_temp[3] ),
    .A2(\d3.saw_temp[0] ),
    .B1(_0348_),
    .X(_0770_));
 sky130_fd_sc_hd__nand2_1 _3204_ (.A(\d3.saw_temp[5] ),
    .B(_0348_),
    .Y(_0771_));
 sky130_fd_sc_hd__or4b_2 _3205_ (.A(\d3.saw_temp[6] ),
    .B(_0769_),
    .C(_0770_),
    .D_N(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__a31o_1 _3206_ (.A1(\d3.saw_temp[0] ),
    .A2(_0348_),
    .A3(_0738_),
    .B1(_0310_),
    .X(_0773_));
 sky130_fd_sc_hd__a31o_1 _3207_ (.A1(_0760_),
    .A2(_0768_),
    .A3(_0772_),
    .B1(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__and3_1 _3208_ (.A(_0766_),
    .B(_0767_),
    .C(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__a21oi_1 _3209_ (.A1(_0767_),
    .A2(_0774_),
    .B1(_0766_),
    .Y(_0776_));
 sky130_fd_sc_hd__or2_1 _3210_ (.A(_0775_),
    .B(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__o21ai_1 _3211_ (.A1(_0736_),
    .A2(_0737_),
    .B1(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nor2_2 _3212_ (.A(_0327_),
    .B(\em0.u1.state[1] ),
    .Y(_0779_));
 sky130_fd_sc_hd__or3_1 _3213_ (.A(_0777_),
    .B(_0736_),
    .C(_0737_),
    .X(_0780_));
 sky130_fd_sc_hd__nor2_1 _3214_ (.A(\em0.u1.state[2] ),
    .B(\em0.u1.state[1] ),
    .Y(_0781_));
 sky130_fd_sc_hd__clkbuf_8 _3215_ (.A(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__a32o_1 _3216_ (.A1(_0778_),
    .A2(_0779_),
    .A3(_0780_),
    .B1(_0782_),
    .B2(net66),
    .X(_0096_));
 sky130_fd_sc_hd__nand2_1 _3217_ (.A(\d5.saw_temp[1] ),
    .B(_0328_),
    .Y(_0783_));
 sky130_fd_sc_hd__or2b_1 _3218_ (.A(\d5.saw_temp[7] ),
    .B_N(_0328_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(_0744_),
    .A1(_0784_),
    .S(\d5.saw_temp[0] ),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(_0783_),
    .A1(_0785_),
    .S(_0760_),
    .X(_0786_));
 sky130_fd_sc_hd__a21boi_1 _3221_ (.A1(_0751_),
    .A2(_0786_),
    .B1_N(_0747_),
    .Y(_0787_));
 sky130_fd_sc_hd__nand2_1 _3222_ (.A(\d4.saw_temp[1] ),
    .B(_0347_),
    .Y(_0788_));
 sky130_fd_sc_hd__o22a_1 _3223_ (.A1(\d4.saw_temp[7] ),
    .A2(_0752_),
    .B1(_0759_),
    .B2(\d4.saw_temp[0] ),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(_0788_),
    .A1(_0789_),
    .S(_0760_),
    .X(_0790_));
 sky130_fd_sc_hd__a21boi_1 _3225_ (.A1(_0751_),
    .A2(_0790_),
    .B1_N(_0762_),
    .Y(_0791_));
 sky130_fd_sc_hd__xor2_1 _3226_ (.A(_0787_),
    .B(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__nand2_2 _3227_ (.A(_0768_),
    .B(_0772_),
    .Y(_0793_));
 sky130_fd_sc_hd__or2b_1 _3228_ (.A(\d3.saw_temp[7] ),
    .B_N(_0348_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(_0793_),
    .A1(_0794_),
    .S(\d3.saw_temp[0] ),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_1 _3230_ (.A(\d3.saw_temp[1] ),
    .B(_0348_),
    .Y(_0796_));
 sky130_fd_sc_hd__o21a_1 _3231_ (.A1(_0760_),
    .A2(_0796_),
    .B1(_0751_),
    .X(_0797_));
 sky130_fd_sc_hd__o21ai_1 _3232_ (.A1(_0738_),
    .A2(_0795_),
    .B1(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_1 _3233_ (.A(_0767_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__xnor2_1 _3234_ (.A(_0792_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__o21ai_2 _3235_ (.A1(_0764_),
    .A2(_0775_),
    .B1(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__or3_1 _3236_ (.A(_0764_),
    .B(_0775_),
    .C(_0800_),
    .X(_0802_));
 sky130_fd_sc_hd__nand2_1 _3237_ (.A(_0801_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_1 _3238_ (.A(_0667_),
    .B(_0677_),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_1 _3239_ (.A(\d8.saw_temp[1] ),
    .B(_0337_),
    .Y(_0805_));
 sky130_fd_sc_hd__or2b_1 _3240_ (.A(\d8.saw_temp[7] ),
    .B_N(_0337_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _3241_ (.A0(_0702_),
    .A1(_0806_),
    .S(\d8.saw_temp[0] ),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(_0805_),
    .A1(_0807_),
    .S(_0634_),
    .X(_0808_));
 sky130_fd_sc_hd__a21oi_2 _3243_ (.A1(_0301_),
    .A2(_0697_),
    .B1(_0307_),
    .Y(_0809_));
 sky130_fd_sc_hd__a21o_1 _3244_ (.A1(_0749_),
    .A2(_0808_),
    .B1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_1 _3245_ (.A(\d7.saw_temp[1] ),
    .B(net12),
    .Y(_0811_));
 sky130_fd_sc_hd__or2_1 _3246_ (.A(\d7.saw_temp[7] ),
    .B(_0333_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(_0713_),
    .A1(_0812_),
    .S(\d7.saw_temp[0] ),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(_0811_),
    .A1(_0813_),
    .S(_0646_),
    .X(_0814_));
 sky130_fd_sc_hd__a21o_1 _3249_ (.A1(_0749_),
    .A2(_0814_),
    .B1(_0708_),
    .X(_0815_));
 sky130_fd_sc_hd__xor2_2 _3250_ (.A(_0810_),
    .B(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__nand2_1 _3251_ (.A(\d6.saw_temp[1] ),
    .B(_0346_),
    .Y(_0817_));
 sky130_fd_sc_hd__or2b_1 _3252_ (.A(\d6.saw_temp[7] ),
    .B_N(_0346_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(_0728_),
    .A1(_0818_),
    .S(\d6.saw_temp[0] ),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(_0817_),
    .A1(_0819_),
    .S(_0646_),
    .X(_0820_));
 sky130_fd_sc_hd__a21o_1 _3255_ (.A1(_0750_),
    .A2(_0820_),
    .B1(_0722_),
    .X(_0821_));
 sky130_fd_sc_hd__xnor2_1 _3256_ (.A(_0816_),
    .B(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__o21ai_2 _3257_ (.A1(_0804_),
    .A2(_0692_),
    .B1(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__or3_1 _3258_ (.A(_0804_),
    .B(_0692_),
    .C(_0822_),
    .X(_0824_));
 sky130_fd_sc_hd__a211o_1 _3259_ (.A1(_0823_),
    .A2(_0824_),
    .B1(_0717_),
    .C1(_0732_),
    .X(_0825_));
 sky130_fd_sc_hd__o211ai_2 _3260_ (.A1(_0717_),
    .A2(_0732_),
    .B1(_0823_),
    .C1(_0824_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand2_1 _3261_ (.A(_0825_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__nand2_1 _3262_ (.A(\d11.saw_temp[1] ),
    .B(_0334_),
    .Y(_0828_));
 sky130_fd_sc_hd__or2b_1 _3263_ (.A(\d11.saw_temp[7] ),
    .B_N(_0334_),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(_0664_),
    .A1(_0829_),
    .S(\d11.saw_temp[0] ),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(_0828_),
    .A1(_0830_),
    .S(_0634_),
    .X(_0831_));
 sky130_fd_sc_hd__a21o_1 _3266_ (.A1(_0622_),
    .A2(_0831_),
    .B1(_0659_),
    .X(_0832_));
 sky130_fd_sc_hd__nand2_1 _3267_ (.A(\d10.saw_temp[1] ),
    .B(_0336_),
    .Y(_0833_));
 sky130_fd_sc_hd__or2b_1 _3268_ (.A(\d10.saw_temp[7] ),
    .B_N(_0336_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(_0674_),
    .A1(_0834_),
    .S(\d10.saw_temp[0] ),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(_0833_),
    .A1(_0835_),
    .S(_0634_),
    .X(_0836_));
 sky130_fd_sc_hd__a21o_1 _3271_ (.A1(_0622_),
    .A2(_0836_),
    .B1(_0669_),
    .X(_0837_));
 sky130_fd_sc_hd__xor2_1 _3272_ (.A(_0832_),
    .B(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__nand2_1 _3273_ (.A(\d9.saw_temp[1] ),
    .B(_0335_),
    .Y(_0839_));
 sky130_fd_sc_hd__or2b_1 _3274_ (.A(\d9.saw_temp[7] ),
    .B_N(_0335_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(_0688_),
    .A1(_0840_),
    .S(\d9.saw_temp[0] ),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(_0839_),
    .A1(_0841_),
    .S(_0634_),
    .X(_0842_));
 sky130_fd_sc_hd__a21o_1 _3277_ (.A1(_0622_),
    .A2(_0842_),
    .B1(_0681_),
    .X(_0843_));
 sky130_fd_sc_hd__inv_2 _3278_ (.A(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _3279_ (.A(_0838_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__or2_1 _3280_ (.A(_0838_),
    .B(_0844_),
    .X(_0846_));
 sky130_fd_sc_hd__nand2_1 _3281_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor2_1 _3282_ (.A(_0621_),
    .B(_0631_),
    .Y(_0848_));
 sky130_fd_sc_hd__a21oi_1 _3283_ (.A1(\d2.saw_temp[1] ),
    .A2(_0329_),
    .B1(_0300_),
    .Y(_0849_));
 sky130_fd_sc_hd__or2_1 _3284_ (.A(\d2.saw_temp[7] ),
    .B(_0613_),
    .X(_0850_));
 sky130_fd_sc_hd__o311a_1 _3285_ (.A1(\d2.saw_temp[0] ),
    .A2(_0611_),
    .A3(_0615_),
    .B1(_0850_),
    .C1(_0618_),
    .X(_0851_));
 sky130_fd_sc_hd__o21a_1 _3286_ (.A1(_0849_),
    .A2(_0851_),
    .B1(_0306_),
    .X(_0852_));
 sky130_fd_sc_hd__a21oi_1 _3287_ (.A1(\d1.saw_temp[1] ),
    .A2(_0330_),
    .B1(_0300_),
    .Y(_0853_));
 sky130_fd_sc_hd__or2_1 _3288_ (.A(\d1.saw_temp[7] ),
    .B(_0625_),
    .X(_0854_));
 sky130_fd_sc_hd__o311a_1 _3289_ (.A1(\d1.saw_temp[0] ),
    .A2(_0623_),
    .A3(_0627_),
    .B1(_0854_),
    .C1(_0618_),
    .X(_0855_));
 sky130_fd_sc_hd__o21a_1 _3290_ (.A1(_0853_),
    .A2(_0855_),
    .B1(_0306_),
    .X(_0856_));
 sky130_fd_sc_hd__or4_1 _3291_ (.A(_0620_),
    .B(_0630_),
    .C(_0852_),
    .D(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__o22ai_2 _3292_ (.A1(_0620_),
    .A2(_0852_),
    .B1(_0856_),
    .B2(_0630_),
    .Y(_0858_));
 sky130_fd_sc_hd__nand3_1 _3293_ (.A(_0848_),
    .B(_0857_),
    .C(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__a21o_1 _3294_ (.A1(_0857_),
    .A2(_0858_),
    .B1(_0848_),
    .X(_0860_));
 sky130_fd_sc_hd__nand2_1 _3295_ (.A(\d13.saw_temp[1] ),
    .B(_0344_),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2_2 _3296_ (.A(_0635_),
    .B(_0639_),
    .Y(_0862_));
 sky130_fd_sc_hd__or2_1 _3297_ (.A(\d13.saw_temp[7] ),
    .B(_0345_),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(_0862_),
    .A1(_0863_),
    .S(\d13.saw_temp[0] ),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(_0861_),
    .A1(_0864_),
    .S(_0634_),
    .X(_0865_));
 sky130_fd_sc_hd__a21oi_2 _3300_ (.A1(_0301_),
    .A2(_0635_),
    .B1(_0307_),
    .Y(_0866_));
 sky130_fd_sc_hd__a21oi_1 _3301_ (.A1(_0622_),
    .A2(_0865_),
    .B1(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand3_1 _3302_ (.A(_0859_),
    .B(_0860_),
    .C(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__a21o_1 _3303_ (.A1(_0859_),
    .A2(_0860_),
    .B1(_0867_),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_1 _3304_ (.A(\d12.saw_temp[1] ),
    .B(_0340_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_2 _3305_ (.A(_0647_),
    .B(_0651_),
    .Y(_0871_));
 sky130_fd_sc_hd__or2b_1 _3306_ (.A(\d12.saw_temp[7] ),
    .B_N(_0340_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(_0871_),
    .A1(_0872_),
    .S(\d12.saw_temp[0] ),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _3308_ (.A0(_0870_),
    .A1(_0873_),
    .S(_0646_),
    .X(_0874_));
 sky130_fd_sc_hd__a21oi_2 _3309_ (.A1(_0301_),
    .A2(_0647_),
    .B1(_0307_),
    .Y(_0875_));
 sky130_fd_sc_hd__a21oi_1 _3310_ (.A1(_0749_),
    .A2(_0874_),
    .B1(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__nand3_1 _3311_ (.A(_0868_),
    .B(_0869_),
    .C(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__a21o_1 _3312_ (.A1(_0868_),
    .A2(_0869_),
    .B1(_0876_),
    .X(_0878_));
 sky130_fd_sc_hd__a31o_1 _3313_ (.A1(_0632_),
    .A2(_0633_),
    .A3(_0642_),
    .B1(_0655_),
    .X(_0879_));
 sky130_fd_sc_hd__and3_1 _3314_ (.A(_0877_),
    .B(_0878_),
    .C(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__a21oi_1 _3315_ (.A1(_0877_),
    .A2(_0878_),
    .B1(_0879_),
    .Y(_0881_));
 sky130_fd_sc_hd__or3_1 _3316_ (.A(_0847_),
    .B(_0880_),
    .C(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__o21ai_1 _3317_ (.A1(_0880_),
    .A2(_0881_),
    .B1(_0847_),
    .Y(_0883_));
 sky130_fd_sc_hd__and3_1 _3318_ (.A(_0695_),
    .B(_0882_),
    .C(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__a21oi_1 _3319_ (.A1(_0882_),
    .A2(_0883_),
    .B1(_0695_),
    .Y(_0885_));
 sky130_fd_sc_hd__nor3_1 _3320_ (.A(_0827_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__o21a_1 _3321_ (.A1(_0884_),
    .A2(_0885_),
    .B1(_0827_),
    .X(_0887_));
 sky130_fd_sc_hd__or3_1 _3322_ (.A(_0735_),
    .B(_0886_),
    .C(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__o21ai_1 _3323_ (.A1(_0886_),
    .A2(_0887_),
    .B1(_0735_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_1 _3324_ (.A(_0888_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__xnor2_1 _3325_ (.A(_0803_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__nor2_1 _3326_ (.A(_0780_),
    .B(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_2 _3327_ (.A(\em0.u1.state[2] ),
    .B(_0326_),
    .Y(_0893_));
 sky130_fd_sc_hd__a21o_1 _3328_ (.A1(_0780_),
    .A2(_0891_),
    .B1(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__a22oi_1 _3329_ (.A1(_1710_),
    .A2(net66),
    .B1(_0782_),
    .B2(net95),
    .Y(_0895_));
 sky130_fd_sc_hd__o21ai_1 _3330_ (.A1(_0892_),
    .A2(_0894_),
    .B1(_0895_),
    .Y(_0097_));
 sky130_fd_sc_hd__a32o_1 _3331_ (.A1(_0767_),
    .A2(_0792_),
    .A3(_0798_),
    .B1(_0787_),
    .B2(_0791_),
    .X(_0896_));
 sky130_fd_sc_hd__nand2_1 _3332_ (.A(\d5.saw_temp[2] ),
    .B(_0328_),
    .Y(_0897_));
 sky130_fd_sc_hd__o22a_1 _3333_ (.A1(\d5.saw_temp[7] ),
    .A2(_0783_),
    .B1(_0744_),
    .B2(\d5.saw_temp[1] ),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(_0897_),
    .A1(_0898_),
    .S(_0760_),
    .X(_0899_));
 sky130_fd_sc_hd__a21boi_1 _3335_ (.A1(_0750_),
    .A2(_0899_),
    .B1_N(_0747_),
    .Y(_0900_));
 sky130_fd_sc_hd__o22a_1 _3336_ (.A1(\d4.saw_temp[7] ),
    .A2(_0788_),
    .B1(_0759_),
    .B2(\d4.saw_temp[1] ),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(_0756_),
    .A1(_0901_),
    .S(_0646_),
    .X(_0902_));
 sky130_fd_sc_hd__a21boi_1 _3338_ (.A1(_0750_),
    .A2(_0902_),
    .B1_N(_0762_),
    .Y(_0903_));
 sky130_fd_sc_hd__nand2_1 _3339_ (.A(_0900_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__or2_1 _3340_ (.A(_0900_),
    .B(_0903_),
    .X(_0905_));
 sky130_fd_sc_hd__and2_1 _3341_ (.A(_0904_),
    .B(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__nand2_1 _3342_ (.A(\d3.saw_temp[2] ),
    .B(_0348_),
    .Y(_0907_));
 sky130_fd_sc_hd__o22a_1 _3343_ (.A1(\d3.saw_temp[7] ),
    .A2(_0796_),
    .B1(_0793_),
    .B2(\d3.saw_temp[1] ),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(_0907_),
    .A1(_0908_),
    .S(_0760_),
    .X(_0909_));
 sky130_fd_sc_hd__a21boi_2 _3345_ (.A1(_0751_),
    .A2(_0909_),
    .B1_N(_0767_),
    .Y(_0910_));
 sky130_fd_sc_hd__xnor2_1 _3346_ (.A(_0906_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__a21oi_1 _3347_ (.A1(_0823_),
    .A2(_0826_),
    .B1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__and3_1 _3348_ (.A(_0823_),
    .B(_0826_),
    .C(_0911_),
    .X(_0913_));
 sky130_fd_sc_hd__nor2_1 _3349_ (.A(_0912_),
    .B(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__xnor2_1 _3350_ (.A(_0896_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__or2_1 _3351_ (.A(_0832_),
    .B(_0837_),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _3352_ (.A(\d8.saw_temp[2] ),
    .B(_0337_),
    .Y(_0917_));
 sky130_fd_sc_hd__o22a_1 _3353_ (.A1(\d8.saw_temp[7] ),
    .A2(_0805_),
    .B1(_0702_),
    .B2(\d8.saw_temp[1] ),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _3354_ (.A0(_0917_),
    .A1(_0918_),
    .S(_0634_),
    .X(_0919_));
 sky130_fd_sc_hd__a21o_1 _3355_ (.A1(_0749_),
    .A2(_0919_),
    .B1(_0809_),
    .X(_0920_));
 sky130_fd_sc_hd__nand2_1 _3356_ (.A(\d7.saw_temp[2] ),
    .B(net12),
    .Y(_0921_));
 sky130_fd_sc_hd__o22a_1 _3357_ (.A1(\d7.saw_temp[7] ),
    .A2(_0811_),
    .B1(_0713_),
    .B2(\d7.saw_temp[1] ),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(_0921_),
    .A1(_0922_),
    .S(_0634_),
    .X(_0923_));
 sky130_fd_sc_hd__a21o_1 _3359_ (.A1(_0749_),
    .A2(_0923_),
    .B1(_0708_),
    .X(_0924_));
 sky130_fd_sc_hd__xor2_1 _3360_ (.A(_0920_),
    .B(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__nand2_1 _3361_ (.A(\d6.saw_temp[2] ),
    .B(_0346_),
    .Y(_0926_));
 sky130_fd_sc_hd__o22a_1 _3362_ (.A1(\d6.saw_temp[7] ),
    .A2(_0817_),
    .B1(_0728_),
    .B2(\d6.saw_temp[1] ),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _3363_ (.A0(_0926_),
    .A1(_0927_),
    .S(_0634_),
    .X(_0928_));
 sky130_fd_sc_hd__a21o_1 _3364_ (.A1(_0749_),
    .A2(_0928_),
    .B1(_0722_),
    .X(_0929_));
 sky130_fd_sc_hd__inv_2 _3365_ (.A(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_1 _3366_ (.A(_0925_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__or2_1 _3367_ (.A(_0925_),
    .B(_0930_),
    .X(_0932_));
 sky130_fd_sc_hd__nand2_1 _3368_ (.A(_0931_),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__a21o_1 _3369_ (.A1(_0916_),
    .A2(_0845_),
    .B1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__nand3_1 _3370_ (.A(_0916_),
    .B(_0845_),
    .C(_0933_),
    .Y(_0935_));
 sky130_fd_sc_hd__nor2_1 _3371_ (.A(_0810_),
    .B(_0815_),
    .Y(_0936_));
 sky130_fd_sc_hd__inv_2 _3372_ (.A(_0816_),
    .Y(_0937_));
 sky130_fd_sc_hd__nor2_1 _3373_ (.A(_0937_),
    .B(_0821_),
    .Y(_0938_));
 sky130_fd_sc_hd__a211o_1 _3374_ (.A1(_0934_),
    .A2(_0935_),
    .B1(_0936_),
    .C1(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__o211ai_2 _3375_ (.A1(_0936_),
    .A2(_0938_),
    .B1(_0934_),
    .C1(_0935_),
    .Y(_0940_));
 sky130_fd_sc_hd__and2_1 _3376_ (.A(_0939_),
    .B(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__nand2_1 _3377_ (.A(\d11.saw_temp[2] ),
    .B(_0334_),
    .Y(_0942_));
 sky130_fd_sc_hd__o22a_1 _3378_ (.A1(\d11.saw_temp[7] ),
    .A2(_0828_),
    .B1(_0664_),
    .B2(\d11.saw_temp[1] ),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(_0942_),
    .A1(_0943_),
    .S(_0618_),
    .X(_0944_));
 sky130_fd_sc_hd__a21o_1 _3380_ (.A1(_0622_),
    .A2(_0944_),
    .B1(_0659_),
    .X(_0945_));
 sky130_fd_sc_hd__nand2_1 _3381_ (.A(\d10.saw_temp[2] ),
    .B(_0336_),
    .Y(_0946_));
 sky130_fd_sc_hd__o22a_1 _3382_ (.A1(\d10.saw_temp[7] ),
    .A2(_0833_),
    .B1(_0674_),
    .B2(\d10.saw_temp[1] ),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(_0946_),
    .A1(_0947_),
    .S(_0618_),
    .X(_0948_));
 sky130_fd_sc_hd__a21o_1 _3384_ (.A1(_0622_),
    .A2(_0948_),
    .B1(_0669_),
    .X(_0949_));
 sky130_fd_sc_hd__xor2_2 _3385_ (.A(_0945_),
    .B(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(\d9.saw_temp[2] ),
    .B(_0335_),
    .Y(_0951_));
 sky130_fd_sc_hd__o22a_1 _3387_ (.A1(\d9.saw_temp[7] ),
    .A2(_0839_),
    .B1(_0688_),
    .B2(\d9.saw_temp[1] ),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _3388_ (.A0(_0951_),
    .A1(_0952_),
    .S(_0646_),
    .X(_0953_));
 sky130_fd_sc_hd__a21o_1 _3389_ (.A1(_0749_),
    .A2(_0953_),
    .B1(_0681_),
    .X(_0954_));
 sky130_fd_sc_hd__xnor2_2 _3390_ (.A(_0950_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__a21bo_1 _3391_ (.A1(_0848_),
    .A2(_0858_),
    .B1_N(_0857_),
    .X(_0956_));
 sky130_fd_sc_hd__or3_1 _3392_ (.A(\d2.saw_temp[1] ),
    .B(_0611_),
    .C(_0615_),
    .X(_0957_));
 sky130_fd_sc_hd__nand3b_1 _3393_ (.A_N(\d2.saw_temp[7] ),
    .B(\d2.saw_temp[1] ),
    .C(_0329_),
    .Y(_0958_));
 sky130_fd_sc_hd__a21oi_1 _3394_ (.A1(\d2.saw_temp[2] ),
    .A2(_0329_),
    .B1(_0300_),
    .Y(_0959_));
 sky130_fd_sc_hd__a31o_1 _3395_ (.A1(_0618_),
    .A2(_0957_),
    .A3(_0958_),
    .B1(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__a21o_1 _3396_ (.A1(_0307_),
    .A2(_0960_),
    .B1(_0620_),
    .X(_0961_));
 sky130_fd_sc_hd__a21oi_1 _3397_ (.A1(\d1.saw_temp[2] ),
    .A2(_0330_),
    .B1(_0301_),
    .Y(_0962_));
 sky130_fd_sc_hd__nand3_1 _3398_ (.A(_0560_),
    .B(\d1.saw_temp[1] ),
    .C(_0330_),
    .Y(_0963_));
 sky130_fd_sc_hd__o311a_1 _3399_ (.A1(\d1.saw_temp[1] ),
    .A2(_0623_),
    .A3(_0627_),
    .B1(_0963_),
    .C1(_0618_),
    .X(_0964_));
 sky130_fd_sc_hd__o21a_1 _3400_ (.A1(_0962_),
    .A2(_0964_),
    .B1(_0307_),
    .X(_0965_));
 sky130_fd_sc_hd__nor2_1 _3401_ (.A(_0630_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__xnor2_2 _3402_ (.A(_0961_),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__xor2_2 _3403_ (.A(_0956_),
    .B(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__o22a_1 _3404_ (.A1(\d13.saw_temp[7] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\d13.saw_temp[1] ),
    .X(_0969_));
 sky130_fd_sc_hd__nor2_1 _3405_ (.A(_0682_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__nand2_1 _3406_ (.A(\d13.saw_temp[2] ),
    .B(_0344_),
    .Y(_0971_));
 sky130_fd_sc_hd__o21ai_1 _3407_ (.A1(_0646_),
    .A2(_0971_),
    .B1(_0622_),
    .Y(_0972_));
 sky130_fd_sc_hd__o21ai_2 _3408_ (.A1(_0970_),
    .A2(_0972_),
    .B1(_0633_),
    .Y(_0973_));
 sky130_fd_sc_hd__xnor2_2 _3409_ (.A(_0968_),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__o22a_1 _3410_ (.A1(\d12.saw_temp[7] ),
    .A2(_0870_),
    .B1(_0871_),
    .B2(\d12.saw_temp[1] ),
    .X(_0975_));
 sky130_fd_sc_hd__nor2_1 _3411_ (.A(_0683_),
    .B(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__nand2_1 _3412_ (.A(\d12.saw_temp[2] ),
    .B(_0340_),
    .Y(_0977_));
 sky130_fd_sc_hd__o21ai_1 _3413_ (.A1(_0760_),
    .A2(_0977_),
    .B1(_0750_),
    .Y(_0978_));
 sky130_fd_sc_hd__o21ai_1 _3414_ (.A1(_0976_),
    .A2(_0978_),
    .B1(_0645_),
    .Y(_0979_));
 sky130_fd_sc_hd__xor2_2 _3415_ (.A(_0974_),
    .B(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__and2_1 _3416_ (.A(_0868_),
    .B(_0877_),
    .X(_0981_));
 sky130_fd_sc_hd__xor2_2 _3417_ (.A(_0980_),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__xor2_1 _3418_ (.A(_0955_),
    .B(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__and2b_1 _3419_ (.A_N(_0880_),
    .B(_0882_),
    .X(_0984_));
 sky130_fd_sc_hd__xnor2_1 _3420_ (.A(_0983_),
    .B(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__xnor2_1 _3421_ (.A(_0941_),
    .B(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__nor2_1 _3422_ (.A(_0884_),
    .B(_0886_),
    .Y(_0987_));
 sky130_fd_sc_hd__xnor2_1 _3423_ (.A(_0986_),
    .B(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__xnor2_1 _3424_ (.A(_0915_),
    .B(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__o21a_1 _3425_ (.A1(_0803_),
    .A2(_0890_),
    .B1(_0888_),
    .X(_0990_));
 sky130_fd_sc_hd__or2_1 _3426_ (.A(_0989_),
    .B(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_1 _3427_ (.A(_0989_),
    .B(_0990_),
    .Y(_0992_));
 sky130_fd_sc_hd__nand2_1 _3428_ (.A(_0991_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__xor2_1 _3429_ (.A(_0801_),
    .B(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__nand2_1 _3430_ (.A(_0892_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__or2_1 _3431_ (.A(_0892_),
    .B(_0994_),
    .X(_0996_));
 sky130_fd_sc_hd__a22o_1 _3432_ (.A1(\em0.u1.state[1] ),
    .A2(net95),
    .B1(net96),
    .B2(_0781_),
    .X(_0997_));
 sky130_fd_sc_hd__a31o_1 _3433_ (.A1(_0779_),
    .A2(_0995_),
    .A3(_0996_),
    .B1(_0997_),
    .X(_0098_));
 sky130_fd_sc_hd__a21oi_2 _3434_ (.A1(_0896_),
    .A2(_0914_),
    .B1(_0912_),
    .Y(_0998_));
 sky130_fd_sc_hd__a21bo_1 _3435_ (.A1(_0905_),
    .A2(_0910_),
    .B1_N(_0904_),
    .X(_0999_));
 sky130_fd_sc_hd__nand2_1 _3436_ (.A(\d5.saw_temp[3] ),
    .B(_0328_),
    .Y(_1000_));
 sky130_fd_sc_hd__o22a_1 _3437_ (.A1(\d5.saw_temp[7] ),
    .A2(_0897_),
    .B1(_0744_),
    .B2(\d5.saw_temp[2] ),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(_1000_),
    .A1(_1001_),
    .S(_0760_),
    .X(_1002_));
 sky130_fd_sc_hd__a21boi_1 _3439_ (.A1(_0751_),
    .A2(_1002_),
    .B1_N(_0747_),
    .Y(_1003_));
 sky130_fd_sc_hd__o22a_1 _3440_ (.A1(\d4.saw_temp[7] ),
    .A2(_0756_),
    .B1(_0759_),
    .B2(\d4.saw_temp[2] ),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(_0755_),
    .A1(_1004_),
    .S(_0760_),
    .X(_1005_));
 sky130_fd_sc_hd__a21boi_1 _3442_ (.A1(_0750_),
    .A2(_1005_),
    .B1_N(_0762_),
    .Y(_1006_));
 sky130_fd_sc_hd__nand2_1 _3443_ (.A(_1003_),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__or2_1 _3444_ (.A(_1003_),
    .B(_1006_),
    .X(_1008_));
 sky130_fd_sc_hd__and2_1 _3445_ (.A(_1007_),
    .B(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_1 _3446_ (.A(\d3.saw_temp[3] ),
    .B(_0348_),
    .Y(_1010_));
 sky130_fd_sc_hd__o22a_1 _3447_ (.A1(\d3.saw_temp[7] ),
    .A2(_0907_),
    .B1(_0793_),
    .B2(\d3.saw_temp[2] ),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(_1010_),
    .A1(_1011_),
    .S(_0760_),
    .X(_1012_));
 sky130_fd_sc_hd__a21boi_2 _3449_ (.A1(_0751_),
    .A2(_1012_),
    .B1_N(_0767_),
    .Y(_1013_));
 sky130_fd_sc_hd__xnor2_1 _3450_ (.A(_1009_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__a21oi_1 _3451_ (.A1(_0934_),
    .A2(_0940_),
    .B1(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__and3_1 _3452_ (.A(_0934_),
    .B(_0940_),
    .C(_1014_),
    .X(_1016_));
 sky130_fd_sc_hd__nor2_1 _3453_ (.A(_1015_),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__xnor2_1 _3454_ (.A(_0999_),
    .B(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__o21a_1 _3455_ (.A1(_0920_),
    .A2(_0924_),
    .B1(_0931_),
    .X(_1019_));
 sky130_fd_sc_hd__or2_1 _3456_ (.A(_0945_),
    .B(_0949_),
    .X(_1020_));
 sky130_fd_sc_hd__inv_2 _3457_ (.A(_0950_),
    .Y(_1021_));
 sky130_fd_sc_hd__or2_1 _3458_ (.A(_1021_),
    .B(_0954_),
    .X(_1022_));
 sky130_fd_sc_hd__nand2_1 _3459_ (.A(\d8.saw_temp[3] ),
    .B(_0337_),
    .Y(_1023_));
 sky130_fd_sc_hd__o22a_1 _3460_ (.A1(\d8.saw_temp[7] ),
    .A2(_0917_),
    .B1(_0702_),
    .B2(\d8.saw_temp[2] ),
    .X(_1024_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(_1023_),
    .A1(_1024_),
    .S(_0634_),
    .X(_1025_));
 sky130_fd_sc_hd__a21o_1 _3462_ (.A1(_0622_),
    .A2(_1025_),
    .B1(_0809_),
    .X(_1026_));
 sky130_fd_sc_hd__nand2_1 _3463_ (.A(\d7.saw_temp[3] ),
    .B(net12),
    .Y(_1027_));
 sky130_fd_sc_hd__o22a_1 _3464_ (.A1(\d7.saw_temp[7] ),
    .A2(_0921_),
    .B1(_0713_),
    .B2(\d7.saw_temp[2] ),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _3465_ (.A0(_1027_),
    .A1(_1028_),
    .S(_0634_),
    .X(_1029_));
 sky130_fd_sc_hd__a21o_1 _3466_ (.A1(_0622_),
    .A2(_1029_),
    .B1(_0708_),
    .X(_1030_));
 sky130_fd_sc_hd__nor2_1 _3467_ (.A(_1026_),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__and2_1 _3468_ (.A(_1026_),
    .B(_1030_),
    .X(_1032_));
 sky130_fd_sc_hd__nor2_1 _3469_ (.A(_1031_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _3470_ (.A(\d6.saw_temp[3] ),
    .B(_0346_),
    .Y(_1034_));
 sky130_fd_sc_hd__o22a_1 _3471_ (.A1(\d6.saw_temp[7] ),
    .A2(_0926_),
    .B1(_0728_),
    .B2(\d6.saw_temp[2] ),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _3472_ (.A0(_1034_),
    .A1(_1035_),
    .S(_0646_),
    .X(_1036_));
 sky130_fd_sc_hd__a21o_1 _3473_ (.A1(_0750_),
    .A2(_1036_),
    .B1(_0722_),
    .X(_1037_));
 sky130_fd_sc_hd__xor2_1 _3474_ (.A(_1033_),
    .B(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__a21o_1 _3475_ (.A1(_1020_),
    .A2(_1022_),
    .B1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__inv_2 _3476_ (.A(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__and3_1 _3477_ (.A(_1020_),
    .B(_1022_),
    .C(_1038_),
    .X(_1041_));
 sky130_fd_sc_hd__nor2_1 _3478_ (.A(_1040_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__xnor2_2 _3479_ (.A(_1019_),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _3480_ (.A(\d11.saw_temp[3] ),
    .B(_0334_),
    .Y(_1044_));
 sky130_fd_sc_hd__o22a_1 _3481_ (.A1(\d11.saw_temp[7] ),
    .A2(_0942_),
    .B1(_0664_),
    .B2(\d11.saw_temp[2] ),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(_1044_),
    .A1(_1045_),
    .S(_0634_),
    .X(_1046_));
 sky130_fd_sc_hd__a21o_1 _3483_ (.A1(_0749_),
    .A2(_1046_),
    .B1(_0659_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_1 _3484_ (.A(\d10.saw_temp[3] ),
    .B(_0336_),
    .Y(_1048_));
 sky130_fd_sc_hd__o22a_1 _3485_ (.A1(\d10.saw_temp[7] ),
    .A2(_0946_),
    .B1(_0674_),
    .B2(\d10.saw_temp[2] ),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(_1048_),
    .A1(_1049_),
    .S(_0634_),
    .X(_1050_));
 sky130_fd_sc_hd__a21o_1 _3487_ (.A1(_0749_),
    .A2(_1050_),
    .B1(_0669_),
    .X(_1051_));
 sky130_fd_sc_hd__or2_1 _3488_ (.A(_1047_),
    .B(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__nand2_1 _3489_ (.A(_1047_),
    .B(_1051_),
    .Y(_1053_));
 sky130_fd_sc_hd__and2_1 _3490_ (.A(_1052_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nand2_1 _3491_ (.A(\d9.saw_temp[3] ),
    .B(_0335_),
    .Y(_1055_));
 sky130_fd_sc_hd__o22a_1 _3492_ (.A1(\d9.saw_temp[7] ),
    .A2(_0951_),
    .B1(_0688_),
    .B2(\d9.saw_temp[2] ),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(_1055_),
    .A1(_1056_),
    .S(_0646_),
    .X(_1057_));
 sky130_fd_sc_hd__a21o_1 _3494_ (.A1(_0750_),
    .A2(_1057_),
    .B1(_0681_),
    .X(_1058_));
 sky130_fd_sc_hd__inv_2 _3495_ (.A(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__nand2_1 _3496_ (.A(_1054_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__or2_1 _3497_ (.A(_1054_),
    .B(_1059_),
    .X(_1061_));
 sky130_fd_sc_hd__nand2_2 _3498_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a31o_1 _3499_ (.A1(\d2.saw_temp[7] ),
    .A2(_0329_),
    .A3(_0301_),
    .B1(_0306_),
    .X(_1063_));
 sky130_fd_sc_hd__a31o_2 _3500_ (.A1(\d1.saw_temp[7] ),
    .A2(_0300_),
    .A3(_0330_),
    .B1(_0306_),
    .X(_1064_));
 sky130_fd_sc_hd__a21oi_1 _3501_ (.A1(\d2.saw_temp[3] ),
    .A2(_0329_),
    .B1(_0300_),
    .Y(_1065_));
 sky130_fd_sc_hd__nand3b_1 _3502_ (.A_N(\d2.saw_temp[7] ),
    .B(\d2.saw_temp[2] ),
    .C(_0329_),
    .Y(_1066_));
 sky130_fd_sc_hd__o311a_1 _3503_ (.A1(\d2.saw_temp[2] ),
    .A2(_0611_),
    .A3(_0615_),
    .B1(_1066_),
    .C1(_0618_),
    .X(_1067_));
 sky130_fd_sc_hd__o21ai_1 _3504_ (.A1(_1065_),
    .A2(_1067_),
    .B1(_0306_),
    .Y(_1068_));
 sky130_fd_sc_hd__a21oi_1 _3505_ (.A1(\d1.saw_temp[3] ),
    .A2(_0330_),
    .B1(_0300_),
    .Y(_1069_));
 sky130_fd_sc_hd__nand3_1 _3506_ (.A(_0560_),
    .B(\d1.saw_temp[2] ),
    .C(_0330_),
    .Y(_1070_));
 sky130_fd_sc_hd__o311a_1 _3507_ (.A1(\d1.saw_temp[2] ),
    .A2(_0623_),
    .A3(_0627_),
    .B1(_1070_),
    .C1(_0618_),
    .X(_1071_));
 sky130_fd_sc_hd__o21ai_1 _3508_ (.A1(_1069_),
    .A2(_1071_),
    .B1(_0306_),
    .Y(_1072_));
 sky130_fd_sc_hd__and4_1 _3509_ (.A(_1063_),
    .B(_1064_),
    .C(_1068_),
    .D(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__a22o_1 _3510_ (.A1(_1063_),
    .A2(_1068_),
    .B1(_1072_),
    .B2(_1064_),
    .X(_1074_));
 sky130_fd_sc_hd__and2b_1 _3511_ (.A_N(_1073_),
    .B(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__a2111oi_1 _3512_ (.A1(_0307_),
    .A2(_0960_),
    .B1(_0965_),
    .C1(_0620_),
    .D1(_0630_),
    .Y(_1076_));
 sky130_fd_sc_hd__a21oi_1 _3513_ (.A1(_0956_),
    .A2(_0967_),
    .B1(net20),
    .Y(_1077_));
 sky130_fd_sc_hd__xnor2_2 _3514_ (.A(_1075_),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__o22a_1 _3515_ (.A1(\d13.saw_temp[7] ),
    .A2(_0971_),
    .B1(_0862_),
    .B2(\d13.saw_temp[2] ),
    .X(_1079_));
 sky130_fd_sc_hd__nor2_1 _3516_ (.A(_0682_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2_1 _3517_ (.A(\d13.saw_temp[3] ),
    .B(_0344_),
    .Y(_1081_));
 sky130_fd_sc_hd__nor2_1 _3518_ (.A(_0646_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__o31a_1 _3519_ (.A1(_0310_),
    .A2(_1080_),
    .A3(_1082_),
    .B1(_0633_),
    .X(_1083_));
 sky130_fd_sc_hd__xor2_2 _3520_ (.A(_1078_),
    .B(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__nand2_1 _3521_ (.A(\d12.saw_temp[3] ),
    .B(_0340_),
    .Y(_1085_));
 sky130_fd_sc_hd__o22a_1 _3522_ (.A1(\d12.saw_temp[7] ),
    .A2(_0977_),
    .B1(_0871_),
    .B2(\d12.saw_temp[2] ),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(_1085_),
    .A1(_1086_),
    .S(_0646_),
    .X(_1087_));
 sky130_fd_sc_hd__a21oi_2 _3524_ (.A1(_0750_),
    .A2(_1087_),
    .B1(_0875_),
    .Y(_1088_));
 sky130_fd_sc_hd__xnor2_2 _3525_ (.A(_1084_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__o211a_1 _3526_ (.A1(_0970_),
    .A2(_0972_),
    .B1(_0633_),
    .C1(_0968_),
    .X(_1090_));
 sky130_fd_sc_hd__o211a_1 _3527_ (.A1(_0976_),
    .A2(_0978_),
    .B1(_0645_),
    .C1(_0974_),
    .X(_1091_));
 sky130_fd_sc_hd__nor2_1 _3528_ (.A(_1090_),
    .B(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__xnor2_2 _3529_ (.A(_1089_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__xor2_2 _3530_ (.A(_1062_),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _3531_ (.A(_0980_),
    .B(_0981_),
    .Y(_1095_));
 sky130_fd_sc_hd__a21oi_2 _3532_ (.A1(_0955_),
    .A2(_0982_),
    .B1(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__xnor2_2 _3533_ (.A(_1094_),
    .B(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__xnor2_1 _3534_ (.A(_1043_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__and2b_1 _3535_ (.A_N(_0984_),
    .B(_0983_),
    .X(_1099_));
 sky130_fd_sc_hd__a21o_1 _3536_ (.A1(_0941_),
    .A2(_0985_),
    .B1(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__xor2_1 _3537_ (.A(_1098_),
    .B(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__xor2_1 _3538_ (.A(_1018_),
    .B(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__or2_1 _3539_ (.A(_0986_),
    .B(_0987_),
    .X(_1103_));
 sky130_fd_sc_hd__o21a_1 _3540_ (.A1(_0915_),
    .A2(_0988_),
    .B1(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__xnor2_1 _3541_ (.A(_1102_),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__xnor2_2 _3542_ (.A(_0998_),
    .B(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__o21a_1 _3543_ (.A1(_0801_),
    .A2(_0993_),
    .B1(_0991_),
    .X(_1107_));
 sky130_fd_sc_hd__xor2_2 _3544_ (.A(_1106_),
    .B(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__a21oi_1 _3545_ (.A1(_0995_),
    .A2(_1108_),
    .B1(_0893_),
    .Y(_1109_));
 sky130_fd_sc_hd__o21a_1 _3546_ (.A1(_0995_),
    .A2(_1108_),
    .B1(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__a221o_1 _3547_ (.A1(_1710_),
    .A2(net96),
    .B1(_0782_),
    .B2(\em0.u1.R[11] ),
    .C1(_1110_),
    .X(_0099_));
 sky130_fd_sc_hd__a21o_1 _3548_ (.A1(_0999_),
    .A2(_1017_),
    .B1(_1015_),
    .X(_1111_));
 sky130_fd_sc_hd__and2b_1 _3549_ (.A_N(_1098_),
    .B(_1100_),
    .X(_1112_));
 sky130_fd_sc_hd__nor2_1 _3550_ (.A(_1018_),
    .B(_1101_),
    .Y(_1113_));
 sky130_fd_sc_hd__a21bo_1 _3551_ (.A1(_1008_),
    .A2(_1013_),
    .B1_N(_1007_),
    .X(_1114_));
 sky130_fd_sc_hd__or3_1 _3552_ (.A(_1019_),
    .B(_1040_),
    .C(_1041_),
    .X(_1115_));
 sky130_fd_sc_hd__o22a_1 _3553_ (.A1(\d5.saw_temp[7] ),
    .A2(_1000_),
    .B1(_0744_),
    .B2(\d5.saw_temp[3] ),
    .X(_1116_));
 sky130_fd_sc_hd__nor2_1 _3554_ (.A(_0723_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__a31o_1 _3555_ (.A1(\d5.saw_temp[4] ),
    .A2(_0328_),
    .A3(_0683_),
    .B1(_0310_),
    .X(_1118_));
 sky130_fd_sc_hd__o21a_1 _3556_ (.A1(_1117_),
    .A2(_1118_),
    .B1(_0747_),
    .X(_1119_));
 sky130_fd_sc_hd__o22a_1 _3557_ (.A1(\d4.saw_temp[7] ),
    .A2(_0755_),
    .B1(_0759_),
    .B2(\d4.saw_temp[3] ),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_1 _3558_ (.A(_0723_),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__a31o_1 _3559_ (.A1(\d4.saw_temp[4] ),
    .A2(_0347_),
    .A3(_0683_),
    .B1(_0310_),
    .X(_1122_));
 sky130_fd_sc_hd__o21a_1 _3560_ (.A1(_1121_),
    .A2(_1122_),
    .B1(_0762_),
    .X(_1123_));
 sky130_fd_sc_hd__nand2_1 _3561_ (.A(_1119_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__or2_1 _3562_ (.A(_1119_),
    .B(_1123_),
    .X(_1125_));
 sky130_fd_sc_hd__and2_1 _3563_ (.A(_1124_),
    .B(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__o22a_1 _3564_ (.A1(\d3.saw_temp[7] ),
    .A2(_1010_),
    .B1(_0793_),
    .B2(\d3.saw_temp[3] ),
    .X(_1127_));
 sky130_fd_sc_hd__nor2_1 _3565_ (.A(_0738_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__a31o_1 _3566_ (.A1(\d3.saw_temp[4] ),
    .A2(_0348_),
    .A3(_0738_),
    .B1(_0310_),
    .X(_1129_));
 sky130_fd_sc_hd__o21a_1 _3567_ (.A1(_1128_),
    .A2(_1129_),
    .B1(_0767_),
    .X(_1130_));
 sky130_fd_sc_hd__xnor2_1 _3568_ (.A(_1126_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__a21oi_1 _3569_ (.A1(_1039_),
    .A2(_1115_),
    .B1(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__and3_1 _3570_ (.A(_1039_),
    .B(_1115_),
    .C(_1131_),
    .X(_1133_));
 sky130_fd_sc_hd__nor2_1 _3571_ (.A(_1132_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__xor2_1 _3572_ (.A(_1114_),
    .B(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__inv_2 _3573_ (.A(_1033_),
    .Y(_1136_));
 sky130_fd_sc_hd__o21bai_2 _3574_ (.A1(_1136_),
    .A2(_1037_),
    .B1_N(_1031_),
    .Y(_1137_));
 sky130_fd_sc_hd__o22a_1 _3575_ (.A1(\d8.saw_temp[7] ),
    .A2(_1023_),
    .B1(_0702_),
    .B2(\d8.saw_temp[3] ),
    .X(_1138_));
 sky130_fd_sc_hd__nor2_1 _3576_ (.A(_0683_),
    .B(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__a31o_1 _3577_ (.A1(\d8.saw_temp[4] ),
    .A2(_0337_),
    .A3(_0682_),
    .B1(_0310_),
    .X(_1140_));
 sky130_fd_sc_hd__o21ai_2 _3578_ (.A1(_1139_),
    .A2(_1140_),
    .B1(_0705_),
    .Y(_1141_));
 sky130_fd_sc_hd__o22a_1 _3579_ (.A1(\d7.saw_temp[7] ),
    .A2(_1027_),
    .B1(_0713_),
    .B2(\d7.saw_temp[3] ),
    .X(_1142_));
 sky130_fd_sc_hd__or2_1 _3580_ (.A(_0682_),
    .B(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nand3_1 _3581_ (.A(\d7.saw_temp[4] ),
    .B(net12),
    .C(_0683_),
    .Y(_1144_));
 sky130_fd_sc_hd__a31o_1 _3582_ (.A1(_0749_),
    .A2(_1143_),
    .A3(_1144_),
    .B1(_0708_),
    .X(_1145_));
 sky130_fd_sc_hd__xor2_1 _3583_ (.A(_1141_),
    .B(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__o22a_1 _3584_ (.A1(\d6.saw_temp[7] ),
    .A2(_1034_),
    .B1(_0728_),
    .B2(\d6.saw_temp[3] ),
    .X(_1147_));
 sky130_fd_sc_hd__a31o_1 _3585_ (.A1(\d6.saw_temp[4] ),
    .A2(_0346_),
    .A3(_0640_),
    .B1(_0309_),
    .X(_1148_));
 sky130_fd_sc_hd__o21ba_1 _3586_ (.A1(_0682_),
    .A2(_1147_),
    .B1_N(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__or2_1 _3587_ (.A(_0722_),
    .B(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__inv_2 _3588_ (.A(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand2_1 _3589_ (.A(_1146_),
    .B(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__or2_1 _3590_ (.A(_1146_),
    .B(_1151_),
    .X(_1153_));
 sky130_fd_sc_hd__nand2_1 _3591_ (.A(_1152_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__a21o_1 _3592_ (.A1(_1052_),
    .A2(_1060_),
    .B1(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__nand3_1 _3593_ (.A(_1052_),
    .B(_1060_),
    .C(_1154_),
    .Y(_1156_));
 sky130_fd_sc_hd__nand2_1 _3594_ (.A(_1155_),
    .B(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__xnor2_2 _3595_ (.A(_1137_),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__o22a_1 _3596_ (.A1(\d11.saw_temp[7] ),
    .A2(_1044_),
    .B1(_0664_),
    .B2(\d11.saw_temp[3] ),
    .X(_1159_));
 sky130_fd_sc_hd__or2_1 _3597_ (.A(_0682_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__nand3_1 _3598_ (.A(\d11.saw_temp[4] ),
    .B(_0334_),
    .C(_0682_),
    .Y(_1161_));
 sky130_fd_sc_hd__a31o_1 _3599_ (.A1(_0622_),
    .A2(_1160_),
    .A3(_1161_),
    .B1(_0659_),
    .X(_1162_));
 sky130_fd_sc_hd__o22a_1 _3600_ (.A1(\d10.saw_temp[7] ),
    .A2(_1048_),
    .B1(_0674_),
    .B2(\d10.saw_temp[3] ),
    .X(_1163_));
 sky130_fd_sc_hd__or2_1 _3601_ (.A(_0640_),
    .B(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__nand3_1 _3602_ (.A(\d10.saw_temp[4] ),
    .B(_0336_),
    .C(_0682_),
    .Y(_1165_));
 sky130_fd_sc_hd__a31o_1 _3603_ (.A1(_0622_),
    .A2(_1164_),
    .A3(_1165_),
    .B1(_0669_),
    .X(_1166_));
 sky130_fd_sc_hd__or2_1 _3604_ (.A(_1162_),
    .B(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__nand2_1 _3605_ (.A(_1162_),
    .B(_1166_),
    .Y(_1168_));
 sky130_fd_sc_hd__and2_1 _3606_ (.A(_1167_),
    .B(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__o22a_1 _3607_ (.A1(\d9.saw_temp[7] ),
    .A2(_1055_),
    .B1(_0688_),
    .B2(\d9.saw_temp[3] ),
    .X(_1170_));
 sky130_fd_sc_hd__a31o_1 _3608_ (.A1(\d9.saw_temp[4] ),
    .A2(_0335_),
    .A3(_0682_),
    .B1(_0309_),
    .X(_1171_));
 sky130_fd_sc_hd__o21ba_1 _3609_ (.A1(_0683_),
    .A2(_1170_),
    .B1_N(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__or2_1 _3610_ (.A(_0681_),
    .B(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__inv_2 _3611_ (.A(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_2 _3612_ (.A(_1169_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__or2_1 _3613_ (.A(_1169_),
    .B(_1174_),
    .X(_1176_));
 sky130_fd_sc_hd__nand2_1 _3614_ (.A(_1175_),
    .B(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__nand3b_1 _3615_ (.A_N(\d2.saw_temp[7] ),
    .B(\d2.saw_temp[3] ),
    .C(_0329_),
    .Y(_1178_));
 sky130_fd_sc_hd__o31a_1 _3616_ (.A1(\d2.saw_temp[3] ),
    .A2(_0611_),
    .A3(_0615_),
    .B1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__a31o_1 _3617_ (.A1(\d2.saw_temp[4] ),
    .A2(_0329_),
    .A3(_0610_),
    .B1(_0309_),
    .X(_1180_));
 sky130_fd_sc_hd__o21ba_1 _3618_ (.A1(_0640_),
    .A2(_1179_),
    .B1_N(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__nor2_2 _3619_ (.A(_0620_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__and2b_1 _3620_ (.A_N(\d1.saw_temp[7] ),
    .B(_0330_),
    .X(_1183_));
 sky130_fd_sc_hd__nand2_1 _3621_ (.A(\d1.saw_temp[3] ),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__o31a_1 _3622_ (.A1(\d1.saw_temp[3] ),
    .A2(_0623_),
    .A3(_0627_),
    .B1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__nor2_1 _3623_ (.A(_0640_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a31o_1 _3624_ (.A1(\d1.saw_temp[4] ),
    .A2(_0330_),
    .A3(_0640_),
    .B1(_0309_),
    .X(_1187_));
 sky130_fd_sc_hd__o21ai_4 _3625_ (.A1(_1186_),
    .A2(_1187_),
    .B1(_1064_),
    .Y(_1188_));
 sky130_fd_sc_hd__xnor2_4 _3626_ (.A(_1182_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__o21a_1 _3627_ (.A1(net21),
    .A2(_1073_),
    .B1(_1074_),
    .X(_1190_));
 sky130_fd_sc_hd__a31o_2 _3628_ (.A1(_0956_),
    .A2(_0967_),
    .A3(_1075_),
    .B1(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__xor2_4 _3629_ (.A(_1189_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__o22a_1 _3630_ (.A1(\d13.saw_temp[7] ),
    .A2(_1081_),
    .B1(_0862_),
    .B2(\d13.saw_temp[3] ),
    .X(_1193_));
 sky130_fd_sc_hd__nor2_1 _3631_ (.A(_0682_),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__a311o_1 _3632_ (.A1(\d13.saw_temp[4] ),
    .A2(_0344_),
    .A3(_0682_),
    .B1(_1194_),
    .C1(_0309_),
    .X(_1195_));
 sky130_fd_sc_hd__nand2_1 _3633_ (.A(_0633_),
    .B(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__xnor2_2 _3634_ (.A(_1192_),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__o22a_1 _3635_ (.A1(\d12.saw_temp[7] ),
    .A2(_1085_),
    .B1(_0871_),
    .B2(\d12.saw_temp[3] ),
    .X(_1198_));
 sky130_fd_sc_hd__nor2_1 _3636_ (.A(_0683_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__a31o_1 _3637_ (.A1(\d12.saw_temp[4] ),
    .A2(_0340_),
    .A3(_0683_),
    .B1(_0310_),
    .X(_1200_));
 sky130_fd_sc_hd__o21a_2 _3638_ (.A1(_1199_),
    .A2(_1200_),
    .B1(_0645_),
    .X(_1201_));
 sky130_fd_sc_hd__xor2_2 _3639_ (.A(_1197_),
    .B(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__nand2_1 _3640_ (.A(_1078_),
    .B(_1083_),
    .Y(_1203_));
 sky130_fd_sc_hd__a21boi_2 _3641_ (.A1(_1084_),
    .A2(_1088_),
    .B1_N(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__xnor2_2 _3642_ (.A(_1202_),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__xnor2_2 _3643_ (.A(_1177_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__nor2_1 _3644_ (.A(_1089_),
    .B(_1092_),
    .Y(_1207_));
 sky130_fd_sc_hd__o21bai_2 _3645_ (.A1(_1062_),
    .A2(_1093_),
    .B1_N(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__xor2_2 _3646_ (.A(_1206_),
    .B(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__xnor2_2 _3647_ (.A(_1158_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__and2b_1 _3648_ (.A_N(_1096_),
    .B(_1094_),
    .X(_1211_));
 sky130_fd_sc_hd__a21oi_2 _3649_ (.A1(_1043_),
    .A2(_1097_),
    .B1(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__xnor2_1 _3650_ (.A(_1210_),
    .B(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__xnor2_1 _3651_ (.A(_1135_),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__o21ai_1 _3652_ (.A1(_1112_),
    .A2(_1113_),
    .B1(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__or3_1 _3653_ (.A(_1112_),
    .B(_1113_),
    .C(_1214_),
    .X(_1216_));
 sky130_fd_sc_hd__and2_1 _3654_ (.A(_1215_),
    .B(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__xnor2_2 _3655_ (.A(_1111_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__or2b_1 _3656_ (.A(_1104_),
    .B_N(_1102_),
    .X(_1219_));
 sky130_fd_sc_hd__or2b_1 _3657_ (.A(_0998_),
    .B_N(_1105_),
    .X(_1220_));
 sky130_fd_sc_hd__and2_1 _3658_ (.A(_1219_),
    .B(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__xor2_2 _3659_ (.A(_1218_),
    .B(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__or2b_1 _3660_ (.A(_1107_),
    .B_N(_1106_),
    .X(_1223_));
 sky130_fd_sc_hd__o21ai_2 _3661_ (.A1(_0995_),
    .A2(_1108_),
    .B1(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2_1 _3662_ (.A(_1222_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__or2_1 _3663_ (.A(_1222_),
    .B(_1224_),
    .X(_1226_));
 sky130_fd_sc_hd__a22o_1 _3664_ (.A1(\em0.u1.state[1] ),
    .A2(\em0.u1.R[11] ),
    .B1(net61),
    .B2(_0781_),
    .X(_1227_));
 sky130_fd_sc_hd__a31o_1 _3665_ (.A1(_0779_),
    .A2(_1225_),
    .A3(_1226_),
    .B1(_1227_),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _3666_ (.A(_1111_),
    .B(_1217_),
    .Y(_1228_));
 sky130_fd_sc_hd__a21o_1 _3667_ (.A1(_1114_),
    .A2(_1134_),
    .B1(_1132_),
    .X(_1229_));
 sky130_fd_sc_hd__a21bo_1 _3668_ (.A1(_1125_),
    .A2(_1130_),
    .B1_N(_1124_),
    .X(_1230_));
 sky130_fd_sc_hd__or2b_1 _3669_ (.A(_1157_),
    .B_N(_1137_),
    .X(_1231_));
 sky130_fd_sc_hd__mux2_1 _3670_ (.A0(_0744_),
    .A1(_0784_),
    .S(\d5.saw_temp[4] ),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _3671_ (.A0(_0742_),
    .A1(_1232_),
    .S(_0760_),
    .X(_1233_));
 sky130_fd_sc_hd__a21boi_1 _3672_ (.A1(_0751_),
    .A2(_1233_),
    .B1_N(_0747_),
    .Y(_1234_));
 sky130_fd_sc_hd__or2b_1 _3673_ (.A(\d4.saw_temp[7] ),
    .B_N(_0347_),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _3674_ (.A0(_0759_),
    .A1(_1235_),
    .S(\d4.saw_temp[4] ),
    .X(_1236_));
 sky130_fd_sc_hd__nor2_1 _3675_ (.A(_0738_),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__a31o_1 _3676_ (.A1(\d4.saw_temp[5] ),
    .A2(_0347_),
    .A3(_0723_),
    .B1(_0310_),
    .X(_1238_));
 sky130_fd_sc_hd__o21a_1 _3677_ (.A1(_1237_),
    .A2(_1238_),
    .B1(_0762_),
    .X(_1239_));
 sky130_fd_sc_hd__nand2_1 _3678_ (.A(_1234_),
    .B(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__or2_1 _3679_ (.A(_1234_),
    .B(_1239_),
    .X(_1241_));
 sky130_fd_sc_hd__and2_1 _3680_ (.A(_1240_),
    .B(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(_0793_),
    .A1(_0794_),
    .S(\d3.saw_temp[4] ),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _3682_ (.A0(_0771_),
    .A1(_1243_),
    .S(_0760_),
    .X(_1244_));
 sky130_fd_sc_hd__a21boi_1 _3683_ (.A1(_0751_),
    .A2(_1244_),
    .B1_N(_0767_),
    .Y(_1245_));
 sky130_fd_sc_hd__xnor2_1 _3684_ (.A(_1242_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a21oi_1 _3685_ (.A1(_1155_),
    .A2(_1231_),
    .B1(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__and3_1 _3686_ (.A(_1155_),
    .B(_1231_),
    .C(_1246_),
    .X(_1248_));
 sky130_fd_sc_hd__nor2_1 _3687_ (.A(_1247_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__xnor2_1 _3688_ (.A(_1230_),
    .B(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__mux2_1 _3689_ (.A0(_0702_),
    .A1(_0806_),
    .S(\d8.saw_temp[4] ),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_1 _3690_ (.A0(_0700_),
    .A1(_1251_),
    .S(_0646_),
    .X(_1252_));
 sky130_fd_sc_hd__a21o_1 _3691_ (.A1(_0749_),
    .A2(_1252_),
    .B1(_0809_),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_1 _3692_ (.A0(_0713_),
    .A1(_0812_),
    .S(\d7.saw_temp[4] ),
    .X(_1254_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(_0711_),
    .A1(_1254_),
    .S(_0634_),
    .X(_1255_));
 sky130_fd_sc_hd__a21o_1 _3694_ (.A1(_0749_),
    .A2(_1255_),
    .B1(_0708_),
    .X(_1256_));
 sky130_fd_sc_hd__nor2_1 _3695_ (.A(_1253_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__and2_1 _3696_ (.A(_1253_),
    .B(_1256_),
    .X(_1258_));
 sky130_fd_sc_hd__nor2_1 _3697_ (.A(_1257_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__mux2_1 _3698_ (.A0(_0728_),
    .A1(_0818_),
    .S(\d6.saw_temp[4] ),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_1 _3699_ (.A0(_0726_),
    .A1(_1260_),
    .S(_0646_),
    .X(_1261_));
 sky130_fd_sc_hd__a21o_1 _3700_ (.A1(_0750_),
    .A2(_1261_),
    .B1(_0722_),
    .X(_1262_));
 sky130_fd_sc_hd__xor2_1 _3701_ (.A(_1259_),
    .B(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__a21o_1 _3702_ (.A1(_1167_),
    .A2(_1175_),
    .B1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__inv_2 _3703_ (.A(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__and3_1 _3704_ (.A(_1167_),
    .B(_1175_),
    .C(_1263_),
    .X(_1266_));
 sky130_fd_sc_hd__o21a_1 _3705_ (.A1(_1141_),
    .A2(_1145_),
    .B1(_1152_),
    .X(_1267_));
 sky130_fd_sc_hd__o21a_1 _3706_ (.A1(_1265_),
    .A2(_1266_),
    .B1(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__or3_1 _3707_ (.A(_1267_),
    .B(_1265_),
    .C(_1266_),
    .X(_1269_));
 sky130_fd_sc_hd__and2b_1 _3708_ (.A_N(_1268_),
    .B(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _3709_ (.A0(_0664_),
    .A1(_0829_),
    .S(\d11.saw_temp[4] ),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_1 _3710_ (.A0(_0662_),
    .A1(_1271_),
    .S(_0646_),
    .X(_1272_));
 sky130_fd_sc_hd__a21o_1 _3711_ (.A1(_0749_),
    .A2(_1272_),
    .B1(_0659_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _3712_ (.A0(_0674_),
    .A1(_0834_),
    .S(\d10.saw_temp[4] ),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _3713_ (.A0(_0672_),
    .A1(_1274_),
    .S(_0646_),
    .X(_1275_));
 sky130_fd_sc_hd__a21o_1 _3714_ (.A1(_0749_),
    .A2(_1275_),
    .B1(_0669_),
    .X(_1276_));
 sky130_fd_sc_hd__or2_1 _3715_ (.A(_1273_),
    .B(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__nand2_1 _3716_ (.A(_1273_),
    .B(_1276_),
    .Y(_1278_));
 sky130_fd_sc_hd__and2_1 _3717_ (.A(_1277_),
    .B(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _3718_ (.A0(_0688_),
    .A1(_0840_),
    .S(\d9.saw_temp[4] ),
    .X(_1280_));
 sky130_fd_sc_hd__mux2_1 _3719_ (.A0(_0686_),
    .A1(_1280_),
    .S(_0646_),
    .X(_1281_));
 sky130_fd_sc_hd__a21o_1 _3720_ (.A1(_0750_),
    .A2(_1281_),
    .B1(_0681_),
    .X(_1282_));
 sky130_fd_sc_hd__inv_2 _3721_ (.A(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__nand2_1 _3722_ (.A(_1279_),
    .B(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__or2_1 _3723_ (.A(_1279_),
    .B(_1283_),
    .X(_1285_));
 sky130_fd_sc_hd__nand2_2 _3724_ (.A(_1284_),
    .B(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_1 _3725_ (.A(\d2.saw_temp[5] ),
    .B(_0329_),
    .Y(_1287_));
 sky130_fd_sc_hd__nand3b_1 _3726_ (.A_N(\d2.saw_temp[7] ),
    .B(\d2.saw_temp[4] ),
    .C(_0329_),
    .Y(_1288_));
 sky130_fd_sc_hd__o311a_1 _3727_ (.A1(\d2.saw_temp[4] ),
    .A2(_0611_),
    .A3(_0615_),
    .B1(_1288_),
    .C1(_0618_),
    .X(_1289_));
 sky130_fd_sc_hd__a21o_1 _3728_ (.A1(_0610_),
    .A2(_1287_),
    .B1(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__nand2_1 _3729_ (.A(_0622_),
    .B(_1290_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2_1 _3730_ (.A(\d1.saw_temp[5] ),
    .B(_0330_),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _3731_ (.A(\d1.saw_temp[4] ),
    .B(_1183_),
    .Y(_1293_));
 sky130_fd_sc_hd__o311a_1 _3732_ (.A1(\d1.saw_temp[4] ),
    .A2(_0623_),
    .A3(_0627_),
    .B1(_1293_),
    .C1(_0618_),
    .X(_1294_));
 sky130_fd_sc_hd__a21o_1 _3733_ (.A1(_0640_),
    .A2(_1292_),
    .B1(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__nand2_1 _3734_ (.A(_0622_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__and4_1 _3735_ (.A(_1063_),
    .B(_1064_),
    .C(_1291_),
    .D(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__a22oi_2 _3736_ (.A1(_1063_),
    .A2(_1291_),
    .B1(_1296_),
    .B2(_1064_),
    .Y(_1298_));
 sky130_fd_sc_hd__nor2_1 _3737_ (.A(_1297_),
    .B(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__nor3_1 _3738_ (.A(_0620_),
    .B(_1181_),
    .C(_1188_),
    .Y(_1300_));
 sky130_fd_sc_hd__a21o_1 _3739_ (.A1(_1189_),
    .A2(_1191_),
    .B1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__xnor2_2 _3740_ (.A(_1299_),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(_0862_),
    .A1(_0863_),
    .S(\d13.saw_temp[4] ),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _3742_ (.A0(_0638_),
    .A1(_1303_),
    .S(_0646_),
    .X(_1304_));
 sky130_fd_sc_hd__a21o_1 _3743_ (.A1(_0750_),
    .A2(_1304_),
    .B1(_0866_),
    .X(_1305_));
 sky130_fd_sc_hd__xor2_2 _3744_ (.A(_1302_),
    .B(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__mux2_1 _3745_ (.A0(_0871_),
    .A1(_0872_),
    .S(\d12.saw_temp[4] ),
    .X(_1307_));
 sky130_fd_sc_hd__mux2_1 _3746_ (.A0(_0650_),
    .A1(_1307_),
    .S(_0760_),
    .X(_1308_));
 sky130_fd_sc_hd__a21oi_2 _3747_ (.A1(_0751_),
    .A2(_1308_),
    .B1(_0875_),
    .Y(_1309_));
 sky130_fd_sc_hd__xnor2_2 _3748_ (.A(_1306_),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__a32oi_4 _3749_ (.A1(_0633_),
    .A2(_1192_),
    .A3(_1195_),
    .B1(_1197_),
    .B2(_1201_),
    .Y(_1311_));
 sky130_fd_sc_hd__xnor2_2 _3750_ (.A(_1310_),
    .B(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__xor2_2 _3751_ (.A(_1286_),
    .B(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__and2b_1 _3752_ (.A_N(_1204_),
    .B(_1202_),
    .X(_1314_));
 sky130_fd_sc_hd__a31oi_2 _3753_ (.A1(_1175_),
    .A2(_1176_),
    .A3(_1205_),
    .B1(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__xnor2_2 _3754_ (.A(_1313_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__xnor2_1 _3755_ (.A(_1270_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__and2_1 _3756_ (.A(_1206_),
    .B(_1208_),
    .X(_1318_));
 sky130_fd_sc_hd__a21oi_1 _3757_ (.A1(_1158_),
    .A2(_1209_),
    .B1(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__xnor2_1 _3758_ (.A(_1317_),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__xor2_1 _3759_ (.A(_1250_),
    .B(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__nand2_1 _3760_ (.A(_1210_),
    .B(_1212_),
    .Y(_1322_));
 sky130_fd_sc_hd__nor2_1 _3761_ (.A(_1210_),
    .B(_1212_),
    .Y(_1323_));
 sky130_fd_sc_hd__a21oi_1 _3762_ (.A1(_1135_),
    .A2(_1322_),
    .B1(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__xnor2_1 _3763_ (.A(_1321_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__xnor2_1 _3764_ (.A(_1229_),
    .B(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__and3_1 _3765_ (.A(_1215_),
    .B(_1228_),
    .C(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__a21oi_1 _3766_ (.A1(_1215_),
    .A2(_1228_),
    .B1(_1326_),
    .Y(_1328_));
 sky130_fd_sc_hd__nor2_1 _3767_ (.A(_1218_),
    .B(_1221_),
    .Y(_1329_));
 sky130_fd_sc_hd__a21o_1 _3768_ (.A1(_1222_),
    .A2(_1224_),
    .B1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__o21ai_1 _3769_ (.A1(_1327_),
    .A2(_1328_),
    .B1(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__a211o_1 _3770_ (.A1(_1222_),
    .A2(_1224_),
    .B1(_1328_),
    .C1(_1329_),
    .X(_1332_));
 sky130_fd_sc_hd__or2_1 _3771_ (.A(_1327_),
    .B(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__a21oi_1 _3772_ (.A1(_1331_),
    .A2(_1333_),
    .B1(_0893_),
    .Y(_1334_));
 sky130_fd_sc_hd__a221o_1 _3773_ (.A1(_1710_),
    .A2(net61),
    .B1(_0782_),
    .B2(\em0.u1.R[13] ),
    .C1(_1334_),
    .X(_0101_));
 sky130_fd_sc_hd__a21o_1 _3774_ (.A1(_1230_),
    .A2(_1249_),
    .B1(_1247_),
    .X(_1335_));
 sky130_fd_sc_hd__nor2_1 _3775_ (.A(_1317_),
    .B(_1319_),
    .Y(_1336_));
 sky130_fd_sc_hd__nor2_1 _3776_ (.A(_1250_),
    .B(_1320_),
    .Y(_1337_));
 sky130_fd_sc_hd__a21bo_1 _3777_ (.A1(_1241_),
    .A2(_1245_),
    .B1_N(_1240_),
    .X(_1338_));
 sky130_fd_sc_hd__o22a_1 _3778_ (.A1(\d5.saw_temp[7] ),
    .A2(_0742_),
    .B1(_0744_),
    .B2(\d5.saw_temp[5] ),
    .X(_1339_));
 sky130_fd_sc_hd__nand2_1 _3779_ (.A(\d5.saw_temp[6] ),
    .B(_0328_),
    .Y(_1340_));
 sky130_fd_sc_hd__o21a_1 _3780_ (.A1(_0760_),
    .A2(_1340_),
    .B1(_0751_),
    .X(_1341_));
 sky130_fd_sc_hd__o21ai_1 _3781_ (.A1(_0738_),
    .A2(_1339_),
    .B1(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__nand2_1 _3782_ (.A(_0747_),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__mux2_1 _3783_ (.A0(_0759_),
    .A1(_1235_),
    .S(\d4.saw_temp[5] ),
    .X(_1344_));
 sky130_fd_sc_hd__nor2_1 _3784_ (.A(_0738_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__a31o_1 _3785_ (.A1(\d4.saw_temp[6] ),
    .A2(_0347_),
    .A3(_0738_),
    .B1(_0310_),
    .X(_1346_));
 sky130_fd_sc_hd__o21a_1 _3786_ (.A1(_1345_),
    .A2(_1346_),
    .B1(_0762_),
    .X(_1347_));
 sky130_fd_sc_hd__xnor2_1 _3787_ (.A(_1343_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__o22a_1 _3788_ (.A1(\d3.saw_temp[7] ),
    .A2(_0771_),
    .B1(_0793_),
    .B2(\d3.saw_temp[5] ),
    .X(_1349_));
 sky130_fd_sc_hd__nor2_1 _3789_ (.A(_0738_),
    .B(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__a31o_1 _3790_ (.A1(\d3.saw_temp[6] ),
    .A2(_0348_),
    .A3(_0738_),
    .B1(_0310_),
    .X(_1351_));
 sky130_fd_sc_hd__o21a_1 _3791_ (.A1(_1350_),
    .A2(_1351_),
    .B1(_0767_),
    .X(_1352_));
 sky130_fd_sc_hd__xnor2_1 _3792_ (.A(_1348_),
    .B(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__a21oi_1 _3793_ (.A1(_1264_),
    .A2(_1269_),
    .B1(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__and3_1 _3794_ (.A(_1264_),
    .B(_1269_),
    .C(_1353_),
    .X(_1355_));
 sky130_fd_sc_hd__nor2_1 _3795_ (.A(_1354_),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__xor2_1 _3796_ (.A(_1338_),
    .B(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__nor3_1 _3797_ (.A(_1257_),
    .B(_1258_),
    .C(_1262_),
    .Y(_1358_));
 sky130_fd_sc_hd__o22a_1 _3798_ (.A1(\d8.saw_temp[7] ),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\d8.saw_temp[5] ),
    .X(_1359_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(\d8.saw_temp[6] ),
    .B(_0337_),
    .Y(_1360_));
 sky130_fd_sc_hd__o21a_1 _3800_ (.A1(_0634_),
    .A2(_1360_),
    .B1(_0622_),
    .X(_1361_));
 sky130_fd_sc_hd__o21ai_2 _3801_ (.A1(_0682_),
    .A2(_1359_),
    .B1(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__nand2_1 _3802_ (.A(_0705_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__o22a_1 _3803_ (.A1(\d7.saw_temp[7] ),
    .A2(_0711_),
    .B1(_0713_),
    .B2(\d7.saw_temp[5] ),
    .X(_1364_));
 sky130_fd_sc_hd__nand2_1 _3804_ (.A(\d7.saw_temp[6] ),
    .B(net12),
    .Y(_1365_));
 sky130_fd_sc_hd__mux2_1 _3805_ (.A0(_1364_),
    .A1(_1365_),
    .S(_0682_),
    .X(_1366_));
 sky130_fd_sc_hd__a21oi_4 _3806_ (.A1(_0749_),
    .A2(_1366_),
    .B1(_0708_),
    .Y(_1367_));
 sky130_fd_sc_hd__xnor2_1 _3807_ (.A(_1363_),
    .B(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__inv_2 _3808_ (.A(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__o22a_1 _3809_ (.A1(\d6.saw_temp[7] ),
    .A2(_0726_),
    .B1(_0728_),
    .B2(\d6.saw_temp[5] ),
    .X(_1370_));
 sky130_fd_sc_hd__nand2_1 _3810_ (.A(\d6.saw_temp[6] ),
    .B(_0346_),
    .Y(_1371_));
 sky130_fd_sc_hd__mux2_1 _3811_ (.A0(_1370_),
    .A1(_1371_),
    .S(_0683_),
    .X(_1372_));
 sky130_fd_sc_hd__a21o_1 _3812_ (.A1(_0750_),
    .A2(_1372_),
    .B1(_0722_),
    .X(_1373_));
 sky130_fd_sc_hd__nor2_1 _3813_ (.A(_1369_),
    .B(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__and2_1 _3814_ (.A(_1369_),
    .B(_1373_),
    .X(_1375_));
 sky130_fd_sc_hd__or2_1 _3815_ (.A(_1374_),
    .B(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__a21o_1 _3816_ (.A1(_1277_),
    .A2(_1284_),
    .B1(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__nand3_1 _3817_ (.A(_1277_),
    .B(_1284_),
    .C(_1376_),
    .Y(_1378_));
 sky130_fd_sc_hd__o211ai_2 _3818_ (.A1(_1257_),
    .A2(_1358_),
    .B1(_1377_),
    .C1(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__a211o_1 _3819_ (.A1(_1377_),
    .A2(_1378_),
    .B1(_1257_),
    .C1(_1358_),
    .X(_1380_));
 sky130_fd_sc_hd__and2_1 _3820_ (.A(_1379_),
    .B(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__o22a_1 _3821_ (.A1(\d11.saw_temp[7] ),
    .A2(_0662_),
    .B1(_0664_),
    .B2(\d11.saw_temp[5] ),
    .X(_1382_));
 sky130_fd_sc_hd__nand2_1 _3822_ (.A(\d11.saw_temp[6] ),
    .B(_0334_),
    .Y(_1383_));
 sky130_fd_sc_hd__mux2_1 _3823_ (.A0(_1382_),
    .A1(_1383_),
    .S(_0683_),
    .X(_1384_));
 sky130_fd_sc_hd__a21o_1 _3824_ (.A1(_0750_),
    .A2(_1384_),
    .B1(_0659_),
    .X(_1385_));
 sky130_fd_sc_hd__o22a_1 _3825_ (.A1(\d10.saw_temp[7] ),
    .A2(_0672_),
    .B1(_0674_),
    .B2(\d10.saw_temp[5] ),
    .X(_1386_));
 sky130_fd_sc_hd__nand2_1 _3826_ (.A(\d10.saw_temp[6] ),
    .B(_0336_),
    .Y(_1387_));
 sky130_fd_sc_hd__mux2_1 _3827_ (.A0(_1386_),
    .A1(_1387_),
    .S(_0683_),
    .X(_1388_));
 sky130_fd_sc_hd__a21o_1 _3828_ (.A1(_0750_),
    .A2(_1388_),
    .B1(_0669_),
    .X(_1389_));
 sky130_fd_sc_hd__xor2_1 _3829_ (.A(_1385_),
    .B(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__o22a_1 _3830_ (.A1(\d9.saw_temp[7] ),
    .A2(_0686_),
    .B1(_0688_),
    .B2(\d9.saw_temp[5] ),
    .X(_1391_));
 sky130_fd_sc_hd__nand2_1 _3831_ (.A(\d9.saw_temp[6] ),
    .B(_0335_),
    .Y(_1392_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(_1391_),
    .A1(_1392_),
    .S(_0723_),
    .X(_1393_));
 sky130_fd_sc_hd__a21oi_1 _3833_ (.A1(_0751_),
    .A2(_1393_),
    .B1(_0681_),
    .Y(_1394_));
 sky130_fd_sc_hd__and2_1 _3834_ (.A(_1390_),
    .B(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__or2_1 _3835_ (.A(_1390_),
    .B(_1394_),
    .X(_1396_));
 sky130_fd_sc_hd__or2b_2 _3836_ (.A(_1395_),
    .B_N(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__o32a_1 _3837_ (.A1(\d2.saw_temp[5] ),
    .A2(_0611_),
    .A3(_0615_),
    .B1(_1287_),
    .B2(\d2.saw_temp[7] ),
    .X(_1398_));
 sky130_fd_sc_hd__nand2_1 _3838_ (.A(\d2.saw_temp[6] ),
    .B(_0329_),
    .Y(_1399_));
 sky130_fd_sc_hd__mux2_1 _3839_ (.A0(_1398_),
    .A1(_1399_),
    .S(_0640_),
    .X(_1400_));
 sky130_fd_sc_hd__a21o_1 _3840_ (.A1(_0622_),
    .A2(_1400_),
    .B1(_0620_),
    .X(_1401_));
 sky130_fd_sc_hd__o32a_1 _3841_ (.A1(\d1.saw_temp[5] ),
    .A2(_0623_),
    .A3(_0627_),
    .B1(_1292_),
    .B2(\d1.saw_temp[7] ),
    .X(_1402_));
 sky130_fd_sc_hd__nand2_1 _3842_ (.A(\d1.saw_temp[6] ),
    .B(_0330_),
    .Y(_1403_));
 sky130_fd_sc_hd__mux2_1 _3843_ (.A0(_1402_),
    .A1(_1403_),
    .S(_0640_),
    .X(_1404_));
 sky130_fd_sc_hd__a21o_1 _3844_ (.A1(_0622_),
    .A2(_1404_),
    .B1(_0630_),
    .X(_1405_));
 sky130_fd_sc_hd__or2_1 _3845_ (.A(_1401_),
    .B(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__nand2_1 _3846_ (.A(_1401_),
    .B(_1405_),
    .Y(_1407_));
 sky130_fd_sc_hd__and2_1 _3847_ (.A(_1406_),
    .B(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__o21ba_1 _3848_ (.A1(_1300_),
    .A2(_1297_),
    .B1_N(_1298_),
    .X(_1409_));
 sky130_fd_sc_hd__a31o_1 _3849_ (.A1(_1189_),
    .A2(_1191_),
    .A3(_1299_),
    .B1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__xnor2_2 _3850_ (.A(_1408_),
    .B(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__o22a_1 _3851_ (.A1(\d13.saw_temp[7] ),
    .A2(_0638_),
    .B1(_0862_),
    .B2(\d13.saw_temp[5] ),
    .X(_1412_));
 sky130_fd_sc_hd__nand2_1 _3852_ (.A(\d13.saw_temp[6] ),
    .B(_0344_),
    .Y(_1413_));
 sky130_fd_sc_hd__mux2_1 _3853_ (.A0(_1412_),
    .A1(_1413_),
    .S(_0683_),
    .X(_1414_));
 sky130_fd_sc_hd__a21o_1 _3854_ (.A1(_0750_),
    .A2(_1414_),
    .B1(_0866_),
    .X(_1415_));
 sky130_fd_sc_hd__xor2_2 _3855_ (.A(_1411_),
    .B(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__o22a_1 _3856_ (.A1(\d12.saw_temp[7] ),
    .A2(_0650_),
    .B1(_0871_),
    .B2(\d12.saw_temp[5] ),
    .X(_1417_));
 sky130_fd_sc_hd__nand2_1 _3857_ (.A(\d12.saw_temp[6] ),
    .B(_0340_),
    .Y(_1418_));
 sky130_fd_sc_hd__mux2_1 _3858_ (.A0(_1417_),
    .A1(_1418_),
    .S(_0683_),
    .X(_1419_));
 sky130_fd_sc_hd__a21oi_2 _3859_ (.A1(_0751_),
    .A2(_1419_),
    .B1(_0875_),
    .Y(_1420_));
 sky130_fd_sc_hd__xnor2_2 _3860_ (.A(_1416_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__nor2_1 _3861_ (.A(_1302_),
    .B(_1305_),
    .Y(_1422_));
 sky130_fd_sc_hd__a21oi_2 _3862_ (.A1(_1306_),
    .A2(_1309_),
    .B1(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__xnor2_2 _3863_ (.A(_1421_),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__xor2_2 _3864_ (.A(_1397_),
    .B(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__nor2_1 _3865_ (.A(_1310_),
    .B(_1311_),
    .Y(_1426_));
 sky130_fd_sc_hd__o21ba_1 _3866_ (.A1(_1286_),
    .A2(_1312_),
    .B1_N(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__xnor2_2 _3867_ (.A(_1425_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__xnor2_1 _3868_ (.A(_1381_),
    .B(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__and2b_1 _3869_ (.A_N(_1315_),
    .B(_1313_),
    .X(_1430_));
 sky130_fd_sc_hd__a21oi_2 _3870_ (.A1(_1270_),
    .A2(_1316_),
    .B1(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__xnor2_1 _3871_ (.A(_1429_),
    .B(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__xnor2_1 _3872_ (.A(_1357_),
    .B(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__o21ai_1 _3873_ (.A1(_1336_),
    .A2(_1337_),
    .B1(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__or3_1 _3874_ (.A(_1336_),
    .B(_1337_),
    .C(_1433_),
    .X(_1435_));
 sky130_fd_sc_hd__and2_1 _3875_ (.A(_1434_),
    .B(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__xnor2_1 _3876_ (.A(_1335_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__or2b_1 _3877_ (.A(_1324_),
    .B_N(_1321_),
    .X(_1438_));
 sky130_fd_sc_hd__a21boi_1 _3878_ (.A1(_1229_),
    .A2(_1325_),
    .B1_N(_1438_),
    .Y(_1439_));
 sky130_fd_sc_hd__xor2_1 _3879_ (.A(_1437_),
    .B(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__nand3b_2 _3880_ (.A_N(_1327_),
    .B(_1332_),
    .C(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__and2b_1 _3881_ (.A_N(_1327_),
    .B(_1332_),
    .X(_1442_));
 sky130_fd_sc_hd__o21a_1 _3882_ (.A1(_1442_),
    .A2(_1440_),
    .B1(_0779_),
    .X(_1443_));
 sky130_fd_sc_hd__a22o_1 _3883_ (.A1(\em0.u1.state[1] ),
    .A2(\em0.u1.R[13] ),
    .B1(net56),
    .B2(_0782_),
    .X(_1444_));
 sky130_fd_sc_hd__a21o_1 _3884_ (.A1(_1441_),
    .A2(_1443_),
    .B1(_1444_),
    .X(_0102_));
 sky130_fd_sc_hd__nor2_1 _3885_ (.A(_1437_),
    .B(_1439_),
    .Y(_1445_));
 sky130_fd_sc_hd__inv_2 _3886_ (.A(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__nand2_1 _3887_ (.A(_1335_),
    .B(_1436_),
    .Y(_1447_));
 sky130_fd_sc_hd__a21o_1 _3888_ (.A1(_1338_),
    .A2(_1356_),
    .B1(_1354_),
    .X(_1448_));
 sky130_fd_sc_hd__a32o_1 _3889_ (.A1(_0747_),
    .A2(_1342_),
    .A3(_1347_),
    .B1(_1348_),
    .B2(_1352_),
    .X(_1449_));
 sky130_fd_sc_hd__a21oi_1 _3890_ (.A1(_0743_),
    .A2(_1340_),
    .B1(_0738_),
    .Y(_1450_));
 sky130_fd_sc_hd__nor2_1 _3891_ (.A(_0739_),
    .B(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__a41o_1 _3892_ (.A1(\d5.saw_temp[6] ),
    .A2(_0328_),
    .A3(_0739_),
    .A4(_0760_),
    .B1(_0310_),
    .X(_1452_));
 sky130_fd_sc_hd__o21a_1 _3893_ (.A1(_1451_),
    .A2(_1452_),
    .B1(_0747_),
    .X(_1453_));
 sky130_fd_sc_hd__a21boi_1 _3894_ (.A1(\d4.saw_temp[6] ),
    .A2(_0347_),
    .B1_N(_0758_),
    .Y(_1454_));
 sky130_fd_sc_hd__o21a_1 _3895_ (.A1(_0738_),
    .A2(_1454_),
    .B1(_0753_),
    .X(_1455_));
 sky130_fd_sc_hd__and4b_1 _3896_ (.A_N(\d4.saw_temp[7] ),
    .B(\d4.saw_temp[6] ),
    .C(_0347_),
    .D(_0760_),
    .X(_1456_));
 sky130_fd_sc_hd__o31a_1 _3897_ (.A1(_0310_),
    .A2(_1455_),
    .A3(_1456_),
    .B1(_0762_),
    .X(_1457_));
 sky130_fd_sc_hd__xor2_1 _3898_ (.A(_1453_),
    .B(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__a21boi_1 _3899_ (.A1(\d3.saw_temp[6] ),
    .A2(_0348_),
    .B1_N(_0772_),
    .Y(_1459_));
 sky130_fd_sc_hd__o21a_1 _3900_ (.A1(_0738_),
    .A2(_1459_),
    .B1(_0768_),
    .X(_1460_));
 sky130_fd_sc_hd__and4b_1 _3901_ (.A_N(\d3.saw_temp[7] ),
    .B(\d3.saw_temp[6] ),
    .C(_0348_),
    .D(_0760_),
    .X(_1461_));
 sky130_fd_sc_hd__o31a_1 _3902_ (.A1(_0310_),
    .A2(_1460_),
    .A3(_1461_),
    .B1(_0767_),
    .X(_1462_));
 sky130_fd_sc_hd__and2_1 _3903_ (.A(_1458_),
    .B(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__nor2_1 _3904_ (.A(_1458_),
    .B(_1462_),
    .Y(_1464_));
 sky130_fd_sc_hd__or2_1 _3905_ (.A(_1463_),
    .B(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__a21oi_1 _3906_ (.A1(_1377_),
    .A2(_1379_),
    .B1(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__and3_1 _3907_ (.A(_1377_),
    .B(_1379_),
    .C(_1465_),
    .X(_1467_));
 sky130_fd_sc_hd__nor2_1 _3908_ (.A(_1466_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__xnor2_1 _3909_ (.A(_1449_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__a31oi_4 _3910_ (.A1(_0705_),
    .A2(_1362_),
    .A3(_1367_),
    .B1(_1374_),
    .Y(_1470_));
 sky130_fd_sc_hd__nor2_1 _3911_ (.A(_1385_),
    .B(_1389_),
    .Y(_1471_));
 sky130_fd_sc_hd__a21o_1 _3912_ (.A1(_0701_),
    .A2(_1360_),
    .B1(_0723_),
    .X(_1472_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(_0697_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__or3_1 _3914_ (.A(_0683_),
    .B(_0697_),
    .C(_1360_),
    .X(_1474_));
 sky130_fd_sc_hd__a31o_1 _3915_ (.A1(_0751_),
    .A2(_1473_),
    .A3(_1474_),
    .B1(_0809_),
    .X(_1475_));
 sky130_fd_sc_hd__a21o_1 _3916_ (.A1(_0712_),
    .A2(_1365_),
    .B1(_0723_),
    .X(_1476_));
 sky130_fd_sc_hd__nand2_1 _3917_ (.A(_0707_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__o31a_1 _3918_ (.A1(_0723_),
    .A2(_0707_),
    .A3(_1365_),
    .B1(_0750_),
    .X(_1478_));
 sky130_fd_sc_hd__a21oi_2 _3919_ (.A1(_1477_),
    .A2(_1478_),
    .B1(_0708_),
    .Y(_1479_));
 sky130_fd_sc_hd__xor2_1 _3920_ (.A(_1475_),
    .B(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__a21o_1 _3921_ (.A1(_0727_),
    .A2(_1371_),
    .B1(_0723_),
    .X(_1481_));
 sky130_fd_sc_hd__nand2_1 _3922_ (.A(_0721_),
    .B(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__o311a_1 _3923_ (.A1(_0738_),
    .A2(_0721_),
    .A3(_1371_),
    .B1(_1482_),
    .C1(_0751_),
    .X(_1483_));
 sky130_fd_sc_hd__nor2_1 _3924_ (.A(_0722_),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__xnor2_1 _3925_ (.A(_1480_),
    .B(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__o21ai_2 _3926_ (.A1(_1471_),
    .A2(_1395_),
    .B1(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__or3_1 _3927_ (.A(_1471_),
    .B(_1395_),
    .C(_1485_),
    .X(_1487_));
 sky130_fd_sc_hd__and2_1 _3928_ (.A(_1486_),
    .B(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__xnor2_2 _3929_ (.A(_1470_),
    .B(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__a21o_1 _3930_ (.A1(_0663_),
    .A2(_1383_),
    .B1(_0723_),
    .X(_1490_));
 sky130_fd_sc_hd__nand2_1 _3931_ (.A(_0658_),
    .B(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__or3_1 _3932_ (.A(_0723_),
    .B(_0658_),
    .C(_1383_),
    .X(_1492_));
 sky130_fd_sc_hd__a31o_1 _3933_ (.A1(_0751_),
    .A2(_1491_),
    .A3(_1492_),
    .B1(_0659_),
    .X(_1493_));
 sky130_fd_sc_hd__a21o_1 _3934_ (.A1(_0673_),
    .A2(_1387_),
    .B1(_0723_),
    .X(_1494_));
 sky130_fd_sc_hd__nand2_1 _3935_ (.A(_0668_),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__o31a_1 _3936_ (.A1(_0723_),
    .A2(_0668_),
    .A3(_1387_),
    .B1(_0750_),
    .X(_1496_));
 sky130_fd_sc_hd__a21oi_1 _3937_ (.A1(_1495_),
    .A2(_1496_),
    .B1(_0669_),
    .Y(_1497_));
 sky130_fd_sc_hd__xnor2_1 _3938_ (.A(_1493_),
    .B(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__a21o_1 _3939_ (.A1(_0687_),
    .A2(_1392_),
    .B1(_0738_),
    .X(_1499_));
 sky130_fd_sc_hd__nand2_1 _3940_ (.A(_0680_),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__o31a_1 _3941_ (.A1(_0738_),
    .A2(_0680_),
    .A3(_1392_),
    .B1(_0751_),
    .X(_1501_));
 sky130_fd_sc_hd__a21oi_1 _3942_ (.A1(_1500_),
    .A2(_1501_),
    .B1(_0681_),
    .Y(_1502_));
 sky130_fd_sc_hd__nand2_1 _3943_ (.A(_1498_),
    .B(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__or2_1 _3944_ (.A(_1498_),
    .B(_1502_),
    .X(_1504_));
 sky130_fd_sc_hd__and2_1 _3945_ (.A(_1503_),
    .B(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__nor2_1 _3946_ (.A(_0640_),
    .B(_1399_),
    .Y(_1506_));
 sky130_fd_sc_hd__a211o_1 _3947_ (.A1(_0634_),
    .A2(_0615_),
    .B1(_1506_),
    .C1(_0611_),
    .X(_1507_));
 sky130_fd_sc_hd__or3_1 _3948_ (.A(\d2.saw_temp[7] ),
    .B(_0682_),
    .C(_1399_),
    .X(_1508_));
 sky130_fd_sc_hd__a31o_1 _3949_ (.A1(_0749_),
    .A2(_1507_),
    .A3(_1508_),
    .B1(_0620_),
    .X(_1509_));
 sky130_fd_sc_hd__nor2_1 _3950_ (.A(_0640_),
    .B(_1403_),
    .Y(_1510_));
 sky130_fd_sc_hd__a211o_1 _3951_ (.A1(_0634_),
    .A2(_0627_),
    .B1(_1510_),
    .C1(_0623_),
    .X(_1511_));
 sky130_fd_sc_hd__nand2_1 _3952_ (.A(_0560_),
    .B(_1510_),
    .Y(_1512_));
 sky130_fd_sc_hd__a31o_1 _3953_ (.A1(_0749_),
    .A2(_1511_),
    .A3(_1512_),
    .B1(_0630_),
    .X(_1513_));
 sky130_fd_sc_hd__nand2_1 _3954_ (.A(_1509_),
    .B(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__or2_1 _3955_ (.A(_1509_),
    .B(_1513_),
    .X(_1515_));
 sky130_fd_sc_hd__nand2_1 _3956_ (.A(_1514_),
    .B(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__a21bo_1 _3957_ (.A1(_1408_),
    .A2(_1410_),
    .B1_N(_1406_),
    .X(_1517_));
 sky130_fd_sc_hd__xnor2_2 _3958_ (.A(_1516_),
    .B(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__a21o_1 _3959_ (.A1(_0639_),
    .A2(_1413_),
    .B1(_0723_),
    .X(_1519_));
 sky130_fd_sc_hd__nand2_1 _3960_ (.A(_0635_),
    .B(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__or3_1 _3961_ (.A(_0723_),
    .B(_0635_),
    .C(_1413_),
    .X(_1521_));
 sky130_fd_sc_hd__a31o_1 _3962_ (.A1(_0751_),
    .A2(_1520_),
    .A3(_1521_),
    .B1(_0866_),
    .X(_1522_));
 sky130_fd_sc_hd__xor2_2 _3963_ (.A(_1518_),
    .B(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__a21o_1 _3964_ (.A1(_0651_),
    .A2(_1418_),
    .B1(_0723_),
    .X(_1524_));
 sky130_fd_sc_hd__nand2_1 _3965_ (.A(_0647_),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__o31ai_1 _3966_ (.A1(_0738_),
    .A2(_0647_),
    .A3(_1418_),
    .B1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__o21a_1 _3967_ (.A1(_0310_),
    .A2(_1526_),
    .B1(_0645_),
    .X(_1527_));
 sky130_fd_sc_hd__xnor2_2 _3968_ (.A(_1523_),
    .B(_1527_),
    .Y(_1528_));
 sky130_fd_sc_hd__nor2_1 _3969_ (.A(_1411_),
    .B(_1415_),
    .Y(_1529_));
 sky130_fd_sc_hd__a21oi_2 _3970_ (.A1(_1416_),
    .A2(_1420_),
    .B1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__xnor2_2 _3971_ (.A(_1528_),
    .B(_1530_),
    .Y(_1531_));
 sky130_fd_sc_hd__xor2_2 _3972_ (.A(_1505_),
    .B(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__or2_1 _3973_ (.A(_1397_),
    .B(_1424_),
    .X(_1533_));
 sky130_fd_sc_hd__o21a_1 _3974_ (.A1(_1421_),
    .A2(_1423_),
    .B1(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__xnor2_2 _3975_ (.A(_1532_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__xnor2_2 _3976_ (.A(_1489_),
    .B(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__or2b_1 _3977_ (.A(_1427_),
    .B_N(_1425_),
    .X(_1537_));
 sky130_fd_sc_hd__a21boi_2 _3978_ (.A1(_1381_),
    .A2(_1428_),
    .B1_N(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__xor2_1 _3979_ (.A(_1536_),
    .B(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__xnor2_1 _3980_ (.A(_1469_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__nand2_1 _3981_ (.A(_1429_),
    .B(_1431_),
    .Y(_1541_));
 sky130_fd_sc_hd__nor2_1 _3982_ (.A(_1429_),
    .B(_1431_),
    .Y(_1542_));
 sky130_fd_sc_hd__a21oi_1 _3983_ (.A1(_1357_),
    .A2(_1541_),
    .B1(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__xnor2_1 _3984_ (.A(_1540_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__xnor2_1 _3985_ (.A(_1448_),
    .B(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__a21o_1 _3986_ (.A1(_1434_),
    .A2(_1447_),
    .B1(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__nand3_1 _3987_ (.A(_1434_),
    .B(_1447_),
    .C(_1545_),
    .Y(_1547_));
 sky130_fd_sc_hd__and2_1 _3988_ (.A(_1546_),
    .B(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__and3_1 _3989_ (.A(_1446_),
    .B(_1441_),
    .C(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__a21oi_1 _3990_ (.A1(_1446_),
    .A2(_1441_),
    .B1(_1548_),
    .Y(_1550_));
 sky130_fd_sc_hd__o21a_1 _3991_ (.A1(_1549_),
    .A2(_1550_),
    .B1(_0779_),
    .X(_1551_));
 sky130_fd_sc_hd__a221o_1 _3992_ (.A1(_1710_),
    .A2(net56),
    .B1(_0782_),
    .B2(\em0.u1.R[15] ),
    .C1(_1551_),
    .X(_0103_));
 sky130_fd_sc_hd__inv_2 _3993_ (.A(_1547_),
    .Y(_1552_));
 sky130_fd_sc_hd__a21o_1 _3994_ (.A1(_1449_),
    .A2(_1468_),
    .B1(_1466_),
    .X(_1553_));
 sky130_fd_sc_hd__or2b_1 _3995_ (.A(_1470_),
    .B_N(_1488_),
    .X(_1554_));
 sky130_fd_sc_hd__a21oi_1 _3996_ (.A1(_1453_),
    .A2(_1457_),
    .B1(_1463_),
    .Y(_1555_));
 sky130_fd_sc_hd__a21o_1 _3997_ (.A1(_1486_),
    .A2(_1554_),
    .B1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__nand3_1 _3998_ (.A(_1486_),
    .B(_1554_),
    .C(_1555_),
    .Y(_1557_));
 sky130_fd_sc_hd__and2_1 _3999_ (.A(_1556_),
    .B(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__or2b_1 _4000_ (.A(_1493_),
    .B_N(_1497_),
    .X(_1559_));
 sky130_fd_sc_hd__or2b_1 _4001_ (.A(_1475_),
    .B_N(_1479_),
    .X(_1560_));
 sky130_fd_sc_hd__o31a_1 _4002_ (.A1(_0722_),
    .A2(_1480_),
    .A3(_1483_),
    .B1(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__a21o_1 _4003_ (.A1(_1559_),
    .A2(_1503_),
    .B1(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__nand3_1 _4004_ (.A(_1559_),
    .B(_1503_),
    .C(_1561_),
    .Y(_1563_));
 sky130_fd_sc_hd__and2_1 _4005_ (.A(_1562_),
    .B(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__inv_2 _4006_ (.A(_1518_),
    .Y(_1565_));
 sky130_fd_sc_hd__or2_1 _4007_ (.A(_1565_),
    .B(_1522_),
    .X(_1566_));
 sky130_fd_sc_hd__or2b_1 _4008_ (.A(_1523_),
    .B_N(_1527_),
    .X(_1567_));
 sky130_fd_sc_hd__a21boi_1 _4009_ (.A1(_1514_),
    .A2(_1517_),
    .B1_N(_1515_),
    .Y(_1568_));
 sky130_fd_sc_hd__a21oi_2 _4010_ (.A1(_1566_),
    .A2(_1567_),
    .B1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__and3_1 _4011_ (.A(_1566_),
    .B(_1567_),
    .C(_1568_),
    .X(_1570_));
 sky130_fd_sc_hd__or2_1 _4012_ (.A(_1569_),
    .B(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__and2b_1 _4013_ (.A_N(_1530_),
    .B(_1528_),
    .X(_1572_));
 sky130_fd_sc_hd__a21oi_1 _4014_ (.A1(_1505_),
    .A2(_1531_),
    .B1(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__xor2_1 _4015_ (.A(_1571_),
    .B(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__xnor2_1 _4016_ (.A(_1564_),
    .B(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__or2b_1 _4017_ (.A(_1534_),
    .B_N(_1532_),
    .X(_1576_));
 sky130_fd_sc_hd__a21boi_1 _4018_ (.A1(_1489_),
    .A2(_1535_),
    .B1_N(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__nor2_1 _4019_ (.A(_1575_),
    .B(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_1575_),
    .B(_1577_),
    .Y(_1579_));
 sky130_fd_sc_hd__and2b_1 _4021_ (.A_N(_1578_),
    .B(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__xnor2_1 _4022_ (.A(_1558_),
    .B(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__or2b_1 _4023_ (.A(_1469_),
    .B_N(_1539_),
    .X(_1582_));
 sky130_fd_sc_hd__o21a_1 _4024_ (.A1(_1536_),
    .A2(_1538_),
    .B1(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__xnor2_1 _4025_ (.A(_1581_),
    .B(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__xor2_1 _4026_ (.A(_1553_),
    .B(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__or2b_1 _4027_ (.A(_1543_),
    .B_N(_1540_),
    .X(_1586_));
 sky130_fd_sc_hd__a21boi_1 _4028_ (.A1(_1448_),
    .A2(_1544_),
    .B1_N(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__xnor2_1 _4029_ (.A(_1585_),
    .B(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__a311o_1 _4030_ (.A1(_1446_),
    .A2(_1441_),
    .A3(_1546_),
    .B1(_1552_),
    .C1(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__a31o_1 _4031_ (.A1(_1446_),
    .A2(_1441_),
    .A3(_1546_),
    .B1(_1552_),
    .X(_1590_));
 sky130_fd_sc_hd__a21oi_1 _4032_ (.A1(_1588_),
    .A2(_1590_),
    .B1(_0893_),
    .Y(_1591_));
 sky130_fd_sc_hd__and2b_1 _4033_ (.A_N(\em0.u1.D[12] ),
    .B(\em0.u1.R[19] ),
    .X(_1592_));
 sky130_fd_sc_hd__and2b_1 _4034_ (.A_N(\em0.u1.R[19] ),
    .B(\em0.u1.D[12] ),
    .X(_1593_));
 sky130_fd_sc_hd__inv_2 _4035_ (.A(\em0.u1.D[11] ),
    .Y(_1594_));
 sky130_fd_sc_hd__inv_2 _4036_ (.A(\em0.u1.D[10] ),
    .Y(_1595_));
 sky130_fd_sc_hd__or2b_1 _4037_ (.A(\em0.u1.D[9] ),
    .B_N(\em0.u1.R[16] ),
    .X(_1596_));
 sky130_fd_sc_hd__or2b_1 _4038_ (.A(\em0.u1.R[16] ),
    .B_N(\em0.u1.D[9] ),
    .X(_1597_));
 sky130_fd_sc_hd__nand2_1 _4039_ (.A(_1596_),
    .B(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__and2b_1 _4040_ (.A_N(\em0.u1.R[15] ),
    .B(\em0.u1.D[8] ),
    .X(_1599_));
 sky130_fd_sc_hd__o21ai_1 _4041_ (.A1(_1598_),
    .A2(_1599_),
    .B1(_1596_),
    .Y(_1600_));
 sky130_fd_sc_hd__o21a_1 _4042_ (.A1(_1595_),
    .A2(\em0.u1.R[17] ),
    .B1(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__a21o_1 _4043_ (.A1(_1595_),
    .A2(\em0.u1.R[17] ),
    .B1(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__o21a_1 _4044_ (.A1(_1594_),
    .A2(\em0.u1.R[18] ),
    .B1(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__a21oi_1 _4045_ (.A1(_1594_),
    .A2(\em0.u1.R[18] ),
    .B1(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__or3_1 _4046_ (.A(_1592_),
    .B(_1593_),
    .C(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__or3b_1 _4047_ (.A(\em0.u1.R[20] ),
    .B(_1592_),
    .C_N(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__or2_1 _4048_ (.A(\em0.u1.R[21] ),
    .B(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__or2_1 _4049_ (.A(\em0.u1.R[22] ),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_4 _4050_ (.A(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__a21oi_1 _4051_ (.A1(\em0.u1.D[8] ),
    .A2(_1609_),
    .B1(\em0.u1.R[15] ),
    .Y(_1610_));
 sky130_fd_sc_hd__a31o_1 _4052_ (.A1(\em0.u1.D[8] ),
    .A2(\em0.u1.R[15] ),
    .A3(_1609_),
    .B1(_0326_),
    .X(_1611_));
 sky130_fd_sc_hd__a2bb2o_1 _4053_ (.A1_N(_1610_),
    .A2_N(_1611_),
    .B1(\em0.u1.R[16] ),
    .B2(_0782_),
    .X(_1612_));
 sky130_fd_sc_hd__a21o_1 _4054_ (.A1(_1589_),
    .A2(_1591_),
    .B1(_1612_),
    .X(_0104_));
 sky130_fd_sc_hd__or2_1 _4055_ (.A(_1585_),
    .B(_1587_),
    .X(_1613_));
 sky130_fd_sc_hd__or2_1 _4056_ (.A(_1581_),
    .B(_1583_),
    .X(_1614_));
 sky130_fd_sc_hd__or2b_1 _4057_ (.A(_1584_),
    .B_N(_1553_),
    .X(_1615_));
 sky130_fd_sc_hd__and2_1 _4058_ (.A(_1564_),
    .B(_1574_),
    .X(_1616_));
 sky130_fd_sc_hd__nand2_1 _4059_ (.A(_1569_),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__or2_1 _4060_ (.A(_1569_),
    .B(_1616_),
    .X(_1618_));
 sky130_fd_sc_hd__o2bb2a_1 _4061_ (.A1_N(_1617_),
    .A2_N(_1618_),
    .B1(_1571_),
    .B2(_1573_),
    .X(_1619_));
 sky130_fd_sc_hd__xnor2_2 _4062_ (.A(_1562_),
    .B(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__a21oi_1 _4063_ (.A1(_1558_),
    .A2(_1579_),
    .B1(_1578_),
    .Y(_1621_));
 sky130_fd_sc_hd__xor2_1 _4064_ (.A(_1620_),
    .B(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__xor2_1 _4065_ (.A(_1556_),
    .B(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__and3_1 _4066_ (.A(_1614_),
    .B(_1615_),
    .C(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__a21oi_1 _4067_ (.A1(_1614_),
    .A2(_1615_),
    .B1(_1623_),
    .Y(_1625_));
 sky130_fd_sc_hd__or2_1 _4068_ (.A(_1624_),
    .B(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__a21o_1 _4069_ (.A1(_1613_),
    .A2(_1589_),
    .B1(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__nand3_1 _4070_ (.A(_1613_),
    .B(_1589_),
    .C(_1626_),
    .Y(_1628_));
 sky130_fd_sc_hd__xnor2_1 _4071_ (.A(_1598_),
    .B(_1599_),
    .Y(_1629_));
 sky130_fd_sc_hd__nand2_1 _4072_ (.A(_1609_),
    .B(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__o211a_1 _4073_ (.A1(\em0.u1.R[16] ),
    .A2(_1609_),
    .B1(_1630_),
    .C1(\em0.u1.state[1] ),
    .X(_1631_));
 sky130_fd_sc_hd__a31o_1 _4074_ (.A1(_0326_),
    .A2(_1627_),
    .A3(_1628_),
    .B1(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__or2_1 _4075_ (.A(\em0.u1.state[2] ),
    .B(\em0.u1.state[1] ),
    .X(_1633_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(\em0.u1.R[17] ),
    .A1(_1632_),
    .S(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__clkbuf_1 _4077_ (.A(_1634_),
    .X(_0105_));
 sky130_fd_sc_hd__a2bb2o_2 _4078_ (.A1_N(_1562_),
    .A2_N(_1619_),
    .B1(_1616_),
    .B2(_1569_),
    .X(_1635_));
 sky130_fd_sc_hd__nor2_1 _4079_ (.A(_1620_),
    .B(_1621_),
    .Y(_1636_));
 sky130_fd_sc_hd__and2b_1 _4080_ (.A_N(_1556_),
    .B(_1622_),
    .X(_1637_));
 sky130_fd_sc_hd__nor2_1 _4081_ (.A(_1636_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__xnor2_2 _4082_ (.A(_1635_),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__inv_2 _4083_ (.A(_1625_),
    .Y(_1640_));
 sky130_fd_sc_hd__a31o_1 _4084_ (.A1(_1613_),
    .A2(_1589_),
    .A3(_1640_),
    .B1(_1624_),
    .X(_1641_));
 sky130_fd_sc_hd__xnor2_1 _4085_ (.A(_1639_),
    .B(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__xor2_1 _4086_ (.A(\em0.u1.D[10] ),
    .B(\em0.u1.R[17] ),
    .X(_1643_));
 sky130_fd_sc_hd__xnor2_1 _4087_ (.A(_1600_),
    .B(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__mux2_1 _4088_ (.A0(\em0.u1.R[17] ),
    .A1(_1644_),
    .S(_1609_),
    .X(_1645_));
 sky130_fd_sc_hd__or2_1 _4089_ (.A(_0326_),
    .B(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__o221a_1 _4090_ (.A1(\em0.u1.R[18] ),
    .A2(_1633_),
    .B1(_0893_),
    .B2(_1642_),
    .C1(_1646_),
    .X(_0106_));
 sky130_fd_sc_hd__o21a_1 _4091_ (.A1(_1636_),
    .A2(_1637_),
    .B1(_1635_),
    .X(_1647_));
 sky130_fd_sc_hd__inv_2 _4092_ (.A(_1639_),
    .Y(_1648_));
 sky130_fd_sc_hd__nor2_1 _4093_ (.A(_1648_),
    .B(_1641_),
    .Y(_1649_));
 sky130_fd_sc_hd__xor2_1 _4094_ (.A(\em0.u1.D[11] ),
    .B(\em0.u1.R[18] ),
    .X(_1650_));
 sky130_fd_sc_hd__xnor2_1 _4095_ (.A(_1602_),
    .B(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(\em0.u1.R[18] ),
    .A1(_1651_),
    .S(_1609_),
    .X(_1652_));
 sky130_fd_sc_hd__o22a_1 _4097_ (.A1(\em0.u1.R[19] ),
    .A2(_1633_),
    .B1(_1652_),
    .B2(_0326_),
    .X(_1653_));
 sky130_fd_sc_hd__o31a_1 _4098_ (.A1(_0893_),
    .A2(_1647_),
    .A3(_1649_),
    .B1(_1653_),
    .X(_0107_));
 sky130_fd_sc_hd__nor2_1 _4099_ (.A(_1592_),
    .B(_1593_),
    .Y(_1654_));
 sky130_fd_sc_hd__xnor2_1 _4100_ (.A(_1654_),
    .B(_1604_),
    .Y(_1655_));
 sky130_fd_sc_hd__mux2_1 _4101_ (.A0(\em0.u1.R[19] ),
    .A1(_1655_),
    .S(_1609_),
    .X(_1656_));
 sky130_fd_sc_hd__a22o_1 _4102_ (.A1(net91),
    .A2(_0782_),
    .B1(_1656_),
    .B2(_1710_),
    .X(_0108_));
 sky130_fd_sc_hd__or2b_1 _4103_ (.A(\em0.u1.D[12] ),
    .B_N(\em0.u1.R[19] ),
    .X(_1657_));
 sky130_fd_sc_hd__a21bo_1 _4104_ (.A1(_1657_),
    .A2(_1605_),
    .B1_N(\em0.u1.R[20] ),
    .X(_1658_));
 sky130_fd_sc_hd__nand2_1 _4105_ (.A(_1606_),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__a32o_1 _4106_ (.A1(_1710_),
    .A2(_1609_),
    .A3(_1659_),
    .B1(net67),
    .B2(_0782_),
    .X(_0109_));
 sky130_fd_sc_hd__inv_2 _4107_ (.A(\em0.u1.R[22] ),
    .Y(_1660_));
 sky130_fd_sc_hd__nand2_1 _4108_ (.A(\em0.u1.R[21] ),
    .B(_1606_),
    .Y(_1661_));
 sky130_fd_sc_hd__o21ai_1 _4109_ (.A1(_1660_),
    .A2(_1607_),
    .B1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__a22o_1 _4110_ (.A1(net128),
    .A2(_0782_),
    .B1(_1662_),
    .B2(_1710_),
    .X(_0110_));
 sky130_fd_sc_hd__o221a_1 _4111_ (.A1(\d12.count[8] ),
    .A2(_1715_),
    .B1(_1718_),
    .B2(\d12.count[7] ),
    .C1(_0231_),
    .X(_1663_));
 sky130_fd_sc_hd__a21o_1 _4112_ (.A1(_1872_),
    .A2(\d12.count[5] ),
    .B1(_0238_),
    .X(_1664_));
 sky130_fd_sc_hd__nor4_1 _4113_ (.A(\d12.count[2] ),
    .B(_0229_),
    .C(_0233_),
    .D(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__nand3_1 _4114_ (.A(_0230_),
    .B(_1663_),
    .C(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__a221o_1 _4115_ (.A1(\d12.count[4] ),
    .A2(_1723_),
    .B1(_1777_),
    .B2(\d12.count[3] ),
    .C1(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__a21oi_2 _4116_ (.A1(\d12.count[7] ),
    .A2(_1720_),
    .B1(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__and4_1 _4117_ (.A(\d12.saw_temp[6] ),
    .B(\d12.saw_temp[5] ),
    .C(\d12.saw_temp[2] ),
    .D(\d12.saw_temp[1] ),
    .X(_1669_));
 sky130_fd_sc_hd__and4_1 _4118_ (.A(\d12.saw_temp[4] ),
    .B(\d12.saw_temp[3] ),
    .C(\d12.saw_temp[0] ),
    .D(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__and2_1 _4119_ (.A(\d12.saw_temp[7] ),
    .B(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__o21a_1 _4120_ (.A1(_1671_),
    .A2(_1668_),
    .B1(\d12.saw_temp[0] ),
    .X(_1672_));
 sky130_fd_sc_hd__o21ba_1 _4121_ (.A1(net201),
    .A2(_1668_),
    .B1_N(_1672_),
    .X(_0111_));
 sky130_fd_sc_hd__xor2_1 _4122_ (.A(net154),
    .B(_1672_),
    .X(_0112_));
 sky130_fd_sc_hd__and3_1 _4123_ (.A(\d12.saw_temp[2] ),
    .B(\d12.saw_temp[1] ),
    .C(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__a21oi_1 _4124_ (.A1(\d12.saw_temp[1] ),
    .A2(_1672_),
    .B1(net211),
    .Y(_1674_));
 sky130_fd_sc_hd__nor2_1 _4125_ (.A(_1673_),
    .B(_1674_),
    .Y(_0113_));
 sky130_fd_sc_hd__xor2_1 _4126_ (.A(net149),
    .B(_1673_),
    .X(_0114_));
 sky130_fd_sc_hd__and3_1 _4127_ (.A(\d12.saw_temp[4] ),
    .B(\d12.saw_temp[3] ),
    .C(_1673_),
    .X(_1675_));
 sky130_fd_sc_hd__a21oi_1 _4128_ (.A1(\d12.saw_temp[3] ),
    .A2(_1673_),
    .B1(net176),
    .Y(_1676_));
 sky130_fd_sc_hd__nor2_1 _4129_ (.A(_1675_),
    .B(_1676_),
    .Y(_0115_));
 sky130_fd_sc_hd__xor2_1 _4130_ (.A(net143),
    .B(_1675_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _4131_ (.A(\d12.saw_temp[5] ),
    .B(_1675_),
    .X(_1677_));
 sky130_fd_sc_hd__xor2_1 _4132_ (.A(net101),
    .B(_1677_),
    .X(_0117_));
 sky130_fd_sc_hd__a21oi_1 _4133_ (.A1(_1670_),
    .A2(_1668_),
    .B1(\d12.saw_temp[7] ),
    .Y(_1678_));
 sky130_fd_sc_hd__nor2_1 _4134_ (.A(_1671_),
    .B(_1678_),
    .Y(_0118_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(net190),
    .A1(\em0.u1.Q[0] ),
    .S(\em0.u1.state[3] ),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _4136_ (.A(_1679_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(net179),
    .A1(net92),
    .S(\em0.u1.state[3] ),
    .X(_1680_));
 sky130_fd_sc_hd__clkbuf_1 _4138_ (.A(_1680_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(\em0.mixed_sample[2] ),
    .A1(net78),
    .S(\em0.u1.state[3] ),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_1 _4140_ (.A(_1681_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4141_ (.A0(\em0.mixed_sample[3] ),
    .A1(\em0.u1.Q[3] ),
    .S(\em0.u1.state[3] ),
    .X(_1682_));
 sky130_fd_sc_hd__clkbuf_1 _4142_ (.A(_1682_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4143_ (.A0(\em0.mixed_sample[4] ),
    .A1(net251),
    .S(\em0.u1.state[3] ),
    .X(_1683_));
 sky130_fd_sc_hd__clkbuf_1 _4144_ (.A(_1683_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4145_ (.A0(\em0.mixed_sample[5] ),
    .A1(net208),
    .S(\em0.u1.state[3] ),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _4146_ (.A(_1684_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4147_ (.A0(net187),
    .A1(net88),
    .S(\em0.u1.state[3] ),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _4148_ (.A(_1685_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4149_ (.A0(net188),
    .A1(net63),
    .S(\em0.u1.state[3] ),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_1 _4150_ (.A(_1686_),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _4151_ (.A1(net131),
    .A2(_0782_),
    .B1(_1609_),
    .B2(_1710_),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _4152_ (.A1(_1710_),
    .A2(\em0.u1.Q[0] ),
    .B1(net92),
    .B2(_0782_),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _4153_ (.A1(_1710_),
    .A2(net92),
    .B1(net78),
    .B2(_0782_),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_1 _4154_ (.A1(_1710_),
    .A2(net78),
    .B1(\em0.u1.Q[3] ),
    .B2(_0782_),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _4155_ (.A1(_1710_),
    .A2(net103),
    .B1(net58),
    .B2(_0782_),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _4156_ (.A1(_1710_),
    .A2(net58),
    .B1(\em0.u1.Q[5] ),
    .B2(_0782_),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _4157_ (.A1(_1710_),
    .A2(\em0.u1.Q[5] ),
    .B1(net88),
    .B2(_0782_),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _4158_ (.A1(_1710_),
    .A2(\em0.u1.Q[6] ),
    .B1(net63),
    .B2(_0782_),
    .X(_0134_));
 sky130_fd_sc_hd__xor2_1 _4159_ (.A(_1710_),
    .B(net102),
    .X(_0135_));
 sky130_fd_sc_hd__and3_1 _4160_ (.A(\em0.u1.state[1] ),
    .B(\em0.u1.count[0] ),
    .C(\em0.u1.count[1] ),
    .X(_1687_));
 sky130_fd_sc_hd__a21oi_1 _4161_ (.A1(_1710_),
    .A2(net102),
    .B1(net106),
    .Y(_1688_));
 sky130_fd_sc_hd__nor2_1 _4162_ (.A(_1687_),
    .B(_1688_),
    .Y(_0136_));
 sky130_fd_sc_hd__o22a_1 _4163_ (.A1(_0326_),
    .A2(_1711_),
    .B1(_1687_),
    .B2(net60),
    .X(_0137_));
 sky130_fd_sc_hd__and4_1 _4164_ (.A(\d9.saw_temp[5] ),
    .B(\d9.saw_temp[4] ),
    .C(\d9.saw_temp[1] ),
    .D(\d9.saw_temp[2] ),
    .X(_1689_));
 sky130_fd_sc_hd__and4_1 _4165_ (.A(\d9.saw_temp[6] ),
    .B(\d9.saw_temp[0] ),
    .C(\d9.saw_temp[3] ),
    .D(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__and2_1 _4166_ (.A(\d9.saw_temp[7] ),
    .B(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__a221o_1 _4167_ (.A1(_1735_),
    .A2(\d9.count[1] ),
    .B1(\d9.count[8] ),
    .B2(_1715_),
    .C1(\d9.count[9] ),
    .X(_1692_));
 sky130_fd_sc_hd__a21boi_1 _4168_ (.A1(_1727_),
    .A2(\d9.count[6] ),
    .B1_N(\d9.count[3] ),
    .Y(_1693_));
 sky130_fd_sc_hd__o221a_1 _4169_ (.A1(\d9.count[8] ),
    .A2(_1715_),
    .B1(_1718_),
    .B2(\d9.count[7] ),
    .C1(_2017_),
    .X(_1694_));
 sky130_fd_sc_hd__and4b_1 _4170_ (.A_N(_1692_),
    .B(_2011_),
    .C(_1693_),
    .D(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__a2bb2o_1 _4171_ (.A1_N(\d9.count[2] ),
    .A2_N(_1724_),
    .B1(_1720_),
    .B2(\d9.count[7] ),
    .X(_1696_));
 sky130_fd_sc_hd__a221oi_1 _4172_ (.A1(\d9.count[2] ),
    .A2(_1724_),
    .B1(_1777_),
    .B2(\d9.count[0] ),
    .C1(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__and3_2 _4173_ (.A(_2015_),
    .B(_1695_),
    .C(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__o21a_1 _4174_ (.A1(_1691_),
    .A2(_1698_),
    .B1(\d9.saw_temp[0] ),
    .X(_1699_));
 sky130_fd_sc_hd__nor3_1 _4175_ (.A(net242),
    .B(_1691_),
    .C(_1698_),
    .Y(_1700_));
 sky130_fd_sc_hd__nor2_1 _4176_ (.A(_1699_),
    .B(_1700_),
    .Y(_0138_));
 sky130_fd_sc_hd__xor2_1 _4177_ (.A(net151),
    .B(_1699_),
    .X(_0139_));
 sky130_fd_sc_hd__and3_1 _4178_ (.A(\d9.saw_temp[1] ),
    .B(\d9.saw_temp[2] ),
    .C(_1699_),
    .X(_1701_));
 sky130_fd_sc_hd__a21oi_1 _4179_ (.A1(\d9.saw_temp[1] ),
    .A2(_1699_),
    .B1(net156),
    .Y(_1702_));
 sky130_fd_sc_hd__nor2_1 _4180_ (.A(_1701_),
    .B(_1702_),
    .Y(_0140_));
 sky130_fd_sc_hd__xor2_1 _4181_ (.A(net125),
    .B(_1701_),
    .X(_0141_));
 sky130_fd_sc_hd__and3_1 _4182_ (.A(\d9.saw_temp[4] ),
    .B(\d9.saw_temp[3] ),
    .C(_1701_),
    .X(_1703_));
 sky130_fd_sc_hd__a21oi_1 _4183_ (.A1(\d9.saw_temp[3] ),
    .A2(_1701_),
    .B1(net165),
    .Y(_1704_));
 sky130_fd_sc_hd__nor2_1 _4184_ (.A(_1703_),
    .B(net166),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _4185_ (.A(\d9.saw_temp[5] ),
    .B(_1703_),
    .Y(_1705_));
 sky130_fd_sc_hd__or2_1 _4186_ (.A(\d9.saw_temp[5] ),
    .B(_1703_),
    .X(_1706_));
 sky130_fd_sc_hd__and2_1 _4187_ (.A(_1705_),
    .B(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__clkbuf_1 _4188_ (.A(_1707_),
    .X(_0143_));
 sky130_fd_sc_hd__xnor2_1 _4189_ (.A(net119),
    .B(_1705_),
    .Y(_0144_));
 sky130_fd_sc_hd__a21oi_1 _4190_ (.A1(_1690_),
    .A2(_1698_),
    .B1(net204),
    .Y(_1708_));
 sky130_fd_sc_hd__nor2_1 _4191_ (.A(_1691_),
    .B(_1708_),
    .Y(_0145_));
 sky130_fd_sc_hd__dfrtp_1 _4192_ (.CLK(clknet_leaf_19_clk),
    .D(\p0.nxt_count[0] ),
    .RESET_B(net39),
    .Q(\p0.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4193_ (.CLK(clknet_leaf_18_clk),
    .D(\p0.nxt_count[1] ),
    .RESET_B(net38),
    .Q(\p0.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4194_ (.CLK(clknet_leaf_19_clk),
    .D(\p0.nxt_count[2] ),
    .RESET_B(net39),
    .Q(\p0.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4195_ (.CLK(clknet_leaf_19_clk),
    .D(\p0.nxt_count[3] ),
    .RESET_B(net39),
    .Q(\p0.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4196_ (.CLK(clknet_leaf_22_clk),
    .D(net226),
    .RESET_B(net32),
    .Q(\p0.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4197_ (.CLK(clknet_leaf_22_clk),
    .D(\p0.nxt_count[5] ),
    .RESET_B(net32),
    .Q(\p0.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4198_ (.CLK(clknet_leaf_24_clk),
    .D(\p0.nxt_count[6] ),
    .RESET_B(net32),
    .Q(\p0.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4199_ (.CLK(clknet_leaf_24_clk),
    .D(\p0.nxt_count[7] ),
    .RESET_B(net32),
    .Q(\p0.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4200_ (.CLK(clknet_leaf_13_clk),
    .D(net55),
    .Q(\m0.edgo.delay ));
 sky130_fd_sc_hd__dfxtp_1 _4201_ (.CLK(clknet_leaf_28_clk),
    .D(net54),
    .Q(\m0.edgy.delay ));
 sky130_fd_sc_hd__dfxtp_1 _4202_ (.CLK(clknet_leaf_13_clk),
    .D(net1),
    .Q(\m0.synco.delay ));
 sky130_fd_sc_hd__dfxtp_1 _4203_ (.CLK(clknet_leaf_28_clk),
    .D(net2),
    .Q(\m0.syncy.delay ));
 sky130_fd_sc_hd__dfxtp_1 _4204_ (.CLK(clknet_leaf_13_clk),
    .D(net52),
    .Q(\m0.edgo.in ));
 sky130_fd_sc_hd__dfxtp_1 _4205_ (.CLK(clknet_leaf_28_clk),
    .D(net53),
    .Q(\m0.edgy.in ));
 sky130_fd_sc_hd__dfrtp_1 _4206_ (.CLK(clknet_leaf_28_clk),
    .D(\e0.next_q[0] ),
    .RESET_B(net28),
    .Q(\d1.oct_dwn[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4207_ (.CLK(clknet_leaf_28_clk),
    .D(\e0.next_q[1] ),
    .RESET_B(net28),
    .Q(\d1.oct_dwn[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4208_ (.CLK(clknet_leaf_32_clk),
    .D(\s0.next_q[0] ),
    .RESET_B(net31),
    .Q(\s0.type_switch[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4209_ (.CLK(clknet_leaf_32_clk),
    .D(\s0.next_q[1] ),
    .RESET_B(net31),
    .Q(\s0.type_switch[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4210_ (.CLK(clknet_leaf_37_clk),
    .D(\d1.nxt_count[0] ),
    .RESET_B(net24),
    .Q(\d1.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4211_ (.CLK(clknet_leaf_37_clk),
    .D(\d1.nxt_count[1] ),
    .RESET_B(net24),
    .Q(\d1.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4212_ (.CLK(clknet_leaf_37_clk),
    .D(\d1.nxt_count[2] ),
    .RESET_B(net24),
    .Q(\d1.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4213_ (.CLK(clknet_leaf_37_clk),
    .D(\d1.nxt_count[3] ),
    .RESET_B(net24),
    .Q(\d1.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4214_ (.CLK(clknet_leaf_35_clk),
    .D(\d1.nxt_count[4] ),
    .RESET_B(net24),
    .Q(\d1.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4215_ (.CLK(clknet_leaf_35_clk),
    .D(\d1.nxt_count[5] ),
    .RESET_B(net25),
    .Q(\d1.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4216_ (.CLK(clknet_leaf_35_clk),
    .D(\d1.nxt_count[6] ),
    .RESET_B(net25),
    .Q(\d1.count[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4217_ (.CLK(clknet_leaf_35_clk),
    .D(\d1.nxt_count[7] ),
    .RESET_B(net25),
    .Q(\d1.count[7] ));
 sky130_fd_sc_hd__dfrtp_4 _4218_ (.CLK(clknet_leaf_33_clk),
    .D(net110),
    .RESET_B(net25),
    .Q(\d1.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4219_ (.CLK(clknet_leaf_34_clk),
    .D(\d1.nxt_count[9] ),
    .RESET_B(net25),
    .Q(\d1.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4220_ (.CLK(clknet_leaf_17_clk),
    .D(_0003_),
    .RESET_B(net38),
    .Q(\em0.u1.D[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4221_ (.CLK(clknet_leaf_17_clk),
    .D(_0004_),
    .RESET_B(net38),
    .Q(\em0.u1.D[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4222_ (.CLK(clknet_leaf_17_clk),
    .D(_0005_),
    .RESET_B(net38),
    .Q(\em0.u1.D[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4223_ (.CLK(clknet_leaf_15_clk),
    .D(_0006_),
    .RESET_B(net40),
    .Q(\em0.u1.D[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4224_ (.CLK(clknet_leaf_16_clk),
    .D(_0007_),
    .RESET_B(net40),
    .Q(\em0.u1.D[12] ));
 sky130_fd_sc_hd__dfrtp_2 _4225_ (.CLK(clknet_leaf_26_clk),
    .D(\d2.nxt_count[0] ),
    .RESET_B(net30),
    .Q(\d2.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4226_ (.CLK(clknet_leaf_26_clk),
    .D(\d2.nxt_count[1] ),
    .RESET_B(net30),
    .Q(\d2.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4227_ (.CLK(clknet_leaf_26_clk),
    .D(\d2.nxt_count[2] ),
    .RESET_B(net30),
    .Q(\d2.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4228_ (.CLK(clknet_leaf_28_clk),
    .D(\d2.nxt_count[3] ),
    .RESET_B(net30),
    .Q(\d2.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4229_ (.CLK(clknet_leaf_28_clk),
    .D(\d2.nxt_count[4] ),
    .RESET_B(net30),
    .Q(\d2.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4230_ (.CLK(clknet_leaf_28_clk),
    .D(\d2.nxt_count[5] ),
    .RESET_B(net28),
    .Q(\d2.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4231_ (.CLK(clknet_leaf_26_clk),
    .D(\d2.nxt_count[6] ),
    .RESET_B(net30),
    .Q(\d2.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4232_ (.CLK(clknet_leaf_26_clk),
    .D(\d2.nxt_count[7] ),
    .RESET_B(net30),
    .Q(\d2.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4233_ (.CLK(clknet_leaf_26_clk),
    .D(\d2.nxt_count[8] ),
    .RESET_B(net30),
    .Q(\d2.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4234_ (.CLK(clknet_leaf_26_clk),
    .D(\d2.nxt_count[9] ),
    .RESET_B(net30),
    .Q(\d2.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4235_ (.CLK(clknet_leaf_31_clk),
    .D(_0008_),
    .RESET_B(net31),
    .Q(\d13.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4236_ (.CLK(clknet_leaf_33_clk),
    .D(_0009_),
    .RESET_B(net27),
    .Q(\d13.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4237_ (.CLK(clknet_leaf_32_clk),
    .D(_0010_),
    .RESET_B(net27),
    .Q(\d13.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4238_ (.CLK(clknet_leaf_32_clk),
    .D(_0011_),
    .RESET_B(net27),
    .Q(\d13.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4239_ (.CLK(clknet_leaf_32_clk),
    .D(_0012_),
    .RESET_B(net27),
    .Q(\d13.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4240_ (.CLK(clknet_leaf_32_clk),
    .D(_0013_),
    .RESET_B(net31),
    .Q(\d13.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4241_ (.CLK(clknet_leaf_32_clk),
    .D(_0014_),
    .RESET_B(net31),
    .Q(\d13.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4242_ (.CLK(clknet_leaf_31_clk),
    .D(_0015_),
    .RESET_B(net31),
    .Q(\d13.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4243_ (.CLK(clknet_leaf_27_clk),
    .D(\d3.nxt_count[0] ),
    .RESET_B(net30),
    .Q(\d3.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4244_ (.CLK(clknet_leaf_25_clk),
    .D(\d3.nxt_count[1] ),
    .RESET_B(net30),
    .Q(\d3.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4245_ (.CLK(clknet_leaf_25_clk),
    .D(\d3.nxt_count[2] ),
    .RESET_B(net30),
    .Q(\d3.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4246_ (.CLK(clknet_leaf_25_clk),
    .D(\d3.nxt_count[3] ),
    .RESET_B(net30),
    .Q(\d3.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4247_ (.CLK(clknet_leaf_24_clk),
    .D(\d3.nxt_count[4] ),
    .RESET_B(net30),
    .Q(\d3.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4248_ (.CLK(clknet_leaf_24_clk),
    .D(\d3.nxt_count[5] ),
    .RESET_B(net30),
    .Q(\d3.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4249_ (.CLK(clknet_leaf_24_clk),
    .D(\d3.nxt_count[6] ),
    .RESET_B(net32),
    .Q(\d3.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4250_ (.CLK(clknet_leaf_24_clk),
    .D(\d3.nxt_count[7] ),
    .RESET_B(net32),
    .Q(\d3.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4251_ (.CLK(clknet_leaf_24_clk),
    .D(\d3.nxt_count[8] ),
    .RESET_B(net32),
    .Q(\d3.count[8] ));
 sky130_fd_sc_hd__dfrtp_4 _4252_ (.CLK(clknet_leaf_24_clk),
    .D(\d3.nxt_count[9] ),
    .RESET_B(net32),
    .Q(\d3.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4253_ (.CLK(clknet_leaf_33_clk),
    .D(_0016_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4254_ (.CLK(clknet_leaf_33_clk),
    .D(_0017_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4255_ (.CLK(clknet_leaf_33_clk),
    .D(_0018_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4256_ (.CLK(clknet_leaf_33_clk),
    .D(_0019_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4257_ (.CLK(clknet_leaf_5_clk),
    .D(_0020_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4258_ (.CLK(clknet_leaf_5_clk),
    .D(_0021_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4259_ (.CLK(clknet_leaf_5_clk),
    .D(_0022_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4260_ (.CLK(clknet_leaf_33_clk),
    .D(_0023_),
    .RESET_B(net27),
    .Q(\d2.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4261_ (.CLK(clknet_leaf_28_clk),
    .D(net75),
    .RESET_B(net28),
    .Q(\d4.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4262_ (.CLK(clknet_leaf_28_clk),
    .D(\d4.nxt_count[1] ),
    .RESET_B(net28),
    .Q(\d4.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4263_ (.CLK(clknet_leaf_28_clk),
    .D(\d4.nxt_count[2] ),
    .RESET_B(net28),
    .Q(\d4.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4264_ (.CLK(clknet_leaf_29_clk),
    .D(\d4.nxt_count[3] ),
    .RESET_B(net28),
    .Q(\d4.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4265_ (.CLK(clknet_leaf_29_clk),
    .D(\d4.nxt_count[4] ),
    .RESET_B(net28),
    .Q(\d4.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4266_ (.CLK(clknet_leaf_29_clk),
    .D(\d4.nxt_count[5] ),
    .RESET_B(net28),
    .Q(\d4.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4267_ (.CLK(clknet_leaf_29_clk),
    .D(\d4.nxt_count[6] ),
    .RESET_B(net28),
    .Q(\d4.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4268_ (.CLK(clknet_leaf_29_clk),
    .D(\d4.nxt_count[7] ),
    .RESET_B(net28),
    .Q(\d4.count[7] ));
 sky130_fd_sc_hd__dfrtp_4 _4269_ (.CLK(clknet_leaf_28_clk),
    .D(\d4.nxt_count[8] ),
    .RESET_B(net28),
    .Q(\d4.count[8] ));
 sky130_fd_sc_hd__dfrtp_2 _4270_ (.CLK(clknet_leaf_27_clk),
    .D(net51),
    .RESET_B(net28),
    .Q(\d4.count[9] ));
 sky130_fd_sc_hd__conb_1 _4270__51 (.LO(net51));
 sky130_fd_sc_hd__dfrtp_2 _4271_ (.CLK(clknet_leaf_21_clk),
    .D(_0024_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4272_ (.CLK(clknet_leaf_24_clk),
    .D(_0025_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4273_ (.CLK(clknet_leaf_24_clk),
    .D(_0026_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4274_ (.CLK(clknet_leaf_24_clk),
    .D(_0027_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4275_ (.CLK(clknet_leaf_22_clk),
    .D(_0028_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4276_ (.CLK(clknet_leaf_22_clk),
    .D(_0029_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4277_ (.CLK(clknet_leaf_22_clk),
    .D(_0030_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4278_ (.CLK(clknet_leaf_21_clk),
    .D(_0031_),
    .RESET_B(net32),
    .Q(\d3.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4279_ (.CLK(clknet_leaf_30_clk),
    .D(net83),
    .RESET_B(net28),
    .Q(\d5.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4280_ (.CLK(clknet_leaf_30_clk),
    .D(\d5.nxt_count[1] ),
    .RESET_B(net29),
    .Q(\d5.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4281_ (.CLK(clknet_leaf_30_clk),
    .D(\d5.nxt_count[2] ),
    .RESET_B(net29),
    .Q(\d5.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4282_ (.CLK(clknet_leaf_35_clk),
    .D(\d5.nxt_count[3] ),
    .RESET_B(net29),
    .Q(\d5.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4283_ (.CLK(clknet_leaf_29_clk),
    .D(\d5.nxt_count[4] ),
    .RESET_B(net29),
    .Q(\d5.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4284_ (.CLK(clknet_leaf_29_clk),
    .D(\d5.nxt_count[5] ),
    .RESET_B(net28),
    .Q(\d5.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4285_ (.CLK(clknet_leaf_27_clk),
    .D(\d5.nxt_count[6] ),
    .RESET_B(net28),
    .Q(\d5.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4286_ (.CLK(clknet_leaf_27_clk),
    .D(\d5.nxt_count[7] ),
    .RESET_B(net29),
    .Q(\d5.count[7] ));
 sky130_fd_sc_hd__dfrtp_4 _4287_ (.CLK(clknet_leaf_30_clk),
    .D(\d5.nxt_count[8] ),
    .RESET_B(net29),
    .Q(\d5.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4288_ (.CLK(clknet_leaf_35_clk),
    .D(net50),
    .RESET_B(net25),
    .Q(\d5.count[9] ));
 sky130_fd_sc_hd__conb_1 _4288__50 (.LO(net50));
 sky130_fd_sc_hd__dfrtp_2 _4289_ (.CLK(clknet_leaf_31_clk),
    .D(_0032_),
    .RESET_B(net31),
    .Q(\d4.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4290_ (.CLK(clknet_leaf_31_clk),
    .D(_0033_),
    .RESET_B(net31),
    .Q(\d4.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4291_ (.CLK(clknet_leaf_31_clk),
    .D(_0034_),
    .RESET_B(net31),
    .Q(\d4.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4292_ (.CLK(clknet_leaf_21_clk),
    .D(_0035_),
    .RESET_B(net31),
    .Q(\d4.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4293_ (.CLK(clknet_leaf_21_clk),
    .D(_0036_),
    .RESET_B(net33),
    .Q(\d4.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4294_ (.CLK(clknet_leaf_21_clk),
    .D(_0037_),
    .RESET_B(net31),
    .Q(\d4.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4295_ (.CLK(clknet_leaf_21_clk),
    .D(_0038_),
    .RESET_B(net31),
    .Q(\d4.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4296_ (.CLK(clknet_leaf_31_clk),
    .D(_0039_),
    .RESET_B(net31),
    .Q(\d4.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4297_ (.CLK(clknet_leaf_3_clk),
    .D(\d6.nxt_count[0] ),
    .RESET_B(net26),
    .Q(\d6.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4298_ (.CLK(clknet_leaf_3_clk),
    .D(\d6.nxt_count[1] ),
    .RESET_B(net26),
    .Q(\d6.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4299_ (.CLK(clknet_leaf_3_clk),
    .D(\d6.nxt_count[2] ),
    .RESET_B(net26),
    .Q(\d6.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4300_ (.CLK(clknet_leaf_3_clk),
    .D(\d6.nxt_count[3] ),
    .RESET_B(net26),
    .Q(\d6.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4301_ (.CLK(clknet_leaf_1_clk),
    .D(\d6.nxt_count[4] ),
    .RESET_B(net22),
    .Q(\d6.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4302_ (.CLK(clknet_leaf_1_clk),
    .D(\d6.nxt_count[5] ),
    .RESET_B(net22),
    .Q(\d6.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4303_ (.CLK(clknet_leaf_1_clk),
    .D(\d6.nxt_count[6] ),
    .RESET_B(net22),
    .Q(\d6.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4304_ (.CLK(clknet_leaf_3_clk),
    .D(\d6.nxt_count[7] ),
    .RESET_B(net26),
    .Q(\d6.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4305_ (.CLK(clknet_leaf_3_clk),
    .D(\d6.nxt_count[8] ),
    .RESET_B(net26),
    .Q(\d6.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4306_ (.CLK(clknet_leaf_3_clk),
    .D(net49),
    .RESET_B(net26),
    .Q(\d6.count[9] ));
 sky130_fd_sc_hd__conb_1 _4306__49 (.LO(net49));
 sky130_fd_sc_hd__dfrtp_2 _4307_ (.CLK(clknet_leaf_22_clk),
    .D(_0040_),
    .RESET_B(net33),
    .Q(\d5.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4308_ (.CLK(clknet_leaf_19_clk),
    .D(_0041_),
    .RESET_B(net39),
    .Q(\d5.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4309_ (.CLK(clknet_leaf_19_clk),
    .D(_0042_),
    .RESET_B(net39),
    .Q(\d5.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4310_ (.CLK(clknet_leaf_19_clk),
    .D(_0043_),
    .RESET_B(net39),
    .Q(\d5.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4311_ (.CLK(clknet_leaf_20_clk),
    .D(_0044_),
    .RESET_B(net39),
    .Q(\d5.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4312_ (.CLK(clknet_leaf_20_clk),
    .D(_0045_),
    .RESET_B(net39),
    .Q(\d5.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4313_ (.CLK(clknet_leaf_20_clk),
    .D(_0046_),
    .RESET_B(net39),
    .Q(\d5.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4314_ (.CLK(clknet_leaf_22_clk),
    .D(_0047_),
    .RESET_B(net33),
    .Q(\d5.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4315_ (.CLK(clknet_leaf_33_clk),
    .D(\d7.nxt_count[0] ),
    .RESET_B(net27),
    .Q(\d7.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4316_ (.CLK(clknet_leaf_33_clk),
    .D(\d7.nxt_count[1] ),
    .RESET_B(net27),
    .Q(\d7.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4317_ (.CLK(clknet_leaf_33_clk),
    .D(\d7.nxt_count[2] ),
    .RESET_B(net27),
    .Q(\d7.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4318_ (.CLK(clknet_leaf_33_clk),
    .D(\d7.nxt_count[3] ),
    .RESET_B(net34),
    .Q(\d7.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4319_ (.CLK(clknet_leaf_35_clk),
    .D(\d7.nxt_count[4] ),
    .RESET_B(net25),
    .Q(\d7.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4320_ (.CLK(clknet_leaf_35_clk),
    .D(\d7.nxt_count[5] ),
    .RESET_B(net25),
    .Q(\d7.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4321_ (.CLK(clknet_leaf_30_clk),
    .D(\d7.nxt_count[6] ),
    .RESET_B(net29),
    .Q(\d7.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4322_ (.CLK(clknet_leaf_31_clk),
    .D(\d7.nxt_count[7] ),
    .RESET_B(net31),
    .Q(\d7.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4323_ (.CLK(clknet_leaf_31_clk),
    .D(\d7.nxt_count[8] ),
    .RESET_B(net31),
    .Q(\d7.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4324_ (.CLK(clknet_leaf_31_clk),
    .D(net48),
    .RESET_B(net31),
    .Q(\d7.count[9] ));
 sky130_fd_sc_hd__conb_1 _4324__48 (.LO(net48));
 sky130_fd_sc_hd__dfrtp_4 _4325_ (.CLK(clknet_leaf_6_clk),
    .D(_0048_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4326_ (.CLK(clknet_leaf_6_clk),
    .D(_0049_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4327_ (.CLK(clknet_leaf_6_clk),
    .D(_0050_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4328_ (.CLK(clknet_leaf_7_clk),
    .D(_0051_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4329_ (.CLK(clknet_leaf_7_clk),
    .D(_0052_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4330_ (.CLK(clknet_leaf_7_clk),
    .D(_0053_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4331_ (.CLK(clknet_leaf_6_clk),
    .D(_0054_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4332_ (.CLK(clknet_leaf_6_clk),
    .D(_0055_),
    .RESET_B(net35),
    .Q(\d6.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4333_ (.CLK(clknet_leaf_36_clk),
    .D(net69),
    .RESET_B(net24),
    .Q(\d8.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4334_ (.CLK(clknet_leaf_36_clk),
    .D(\d8.nxt_count[1] ),
    .RESET_B(net24),
    .Q(\d8.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4335_ (.CLK(clknet_leaf_36_clk),
    .D(\d8.nxt_count[2] ),
    .RESET_B(net24),
    .Q(\d8.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4336_ (.CLK(clknet_leaf_36_clk),
    .D(\d8.nxt_count[3] ),
    .RESET_B(net24),
    .Q(\d8.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4337_ (.CLK(clknet_leaf_36_clk),
    .D(\d8.nxt_count[4] ),
    .RESET_B(net24),
    .Q(\d8.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4338_ (.CLK(clknet_leaf_36_clk),
    .D(\d8.nxt_count[5] ),
    .RESET_B(net24),
    .Q(\d8.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4339_ (.CLK(clknet_leaf_36_clk),
    .D(\d8.nxt_count[6] ),
    .RESET_B(net24),
    .Q(\d8.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4340_ (.CLK(clknet_leaf_29_clk),
    .D(\d8.nxt_count[7] ),
    .RESET_B(net28),
    .Q(\d8.count[7] ));
 sky130_fd_sc_hd__dfrtp_4 _4341_ (.CLK(clknet_leaf_29_clk),
    .D(\d8.nxt_count[8] ),
    .RESET_B(net24),
    .Q(\d8.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4342_ (.CLK(clknet_leaf_35_clk),
    .D(net47),
    .RESET_B(net24),
    .Q(\d8.count[9] ));
 sky130_fd_sc_hd__conb_1 _4342__47 (.LO(net47));
 sky130_fd_sc_hd__dfrtp_4 _4343_ (.CLK(clknet_leaf_13_clk),
    .D(_0056_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4344_ (.CLK(clknet_leaf_13_clk),
    .D(_0057_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4345_ (.CLK(clknet_leaf_13_clk),
    .D(_0058_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4346_ (.CLK(clknet_leaf_13_clk),
    .D(_0059_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4347_ (.CLK(clknet_leaf_14_clk),
    .D(_0060_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4348_ (.CLK(clknet_leaf_14_clk),
    .D(_0061_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4349_ (.CLK(clknet_leaf_14_clk),
    .D(_0062_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4350_ (.CLK(clknet_leaf_13_clk),
    .D(_0063_),
    .RESET_B(net40),
    .Q(\d7.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4351_ (.CLK(clknet_leaf_36_clk),
    .D(net77),
    .RESET_B(net24),
    .Q(\d9.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4352_ (.CLK(clknet_leaf_36_clk),
    .D(\d9.nxt_count[1] ),
    .RESET_B(net24),
    .Q(\d9.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4353_ (.CLK(clknet_leaf_36_clk),
    .D(\d9.nxt_count[2] ),
    .RESET_B(net24),
    .Q(\d9.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4354_ (.CLK(clknet_leaf_36_clk),
    .D(\d9.nxt_count[3] ),
    .RESET_B(net24),
    .Q(\d9.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4355_ (.CLK(clknet_leaf_38_clk),
    .D(\d9.nxt_count[4] ),
    .RESET_B(net22),
    .Q(\d9.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4356_ (.CLK(clknet_leaf_38_clk),
    .D(\d9.nxt_count[5] ),
    .RESET_B(net22),
    .Q(\d9.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4357_ (.CLK(clknet_leaf_37_clk),
    .D(\d9.nxt_count[6] ),
    .RESET_B(net22),
    .Q(\d9.count[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4358_ (.CLK(clknet_leaf_37_clk),
    .D(\d9.nxt_count[7] ),
    .RESET_B(net22),
    .Q(\d9.count[7] ));
 sky130_fd_sc_hd__dfrtp_4 _4359_ (.CLK(clknet_leaf_37_clk),
    .D(\d9.nxt_count[8] ),
    .RESET_B(net22),
    .Q(\d9.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4360_ (.CLK(clknet_leaf_37_clk),
    .D(net46),
    .RESET_B(net23),
    .Q(\d9.count[9] ));
 sky130_fd_sc_hd__conb_1 _4360__46 (.LO(net46));
 sky130_fd_sc_hd__dfrtp_2 _4361_ (.CLK(clknet_leaf_7_clk),
    .D(_0064_),
    .RESET_B(net35),
    .Q(\d8.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4362_ (.CLK(clknet_leaf_8_clk),
    .D(_0065_),
    .RESET_B(net36),
    .Q(\d8.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4363_ (.CLK(clknet_leaf_8_clk),
    .D(_0066_),
    .RESET_B(net36),
    .Q(\d8.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4364_ (.CLK(clknet_leaf_8_clk),
    .D(_0067_),
    .RESET_B(net36),
    .Q(\d8.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4365_ (.CLK(clknet_leaf_7_clk),
    .D(_0068_),
    .RESET_B(net36),
    .Q(\d8.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4366_ (.CLK(clknet_leaf_7_clk),
    .D(_0069_),
    .RESET_B(net35),
    .Q(\d8.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4367_ (.CLK(clknet_leaf_7_clk),
    .D(_0070_),
    .RESET_B(net37),
    .Q(\d8.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4368_ (.CLK(clknet_leaf_7_clk),
    .D(_0071_),
    .RESET_B(net37),
    .Q(\d8.saw_temp[7] ));
 sky130_fd_sc_hd__dfstp_1 _4369_ (.CLK(clknet_leaf_17_clk),
    .D(net41),
    .SET_B(net38),
    .Q(\em0.u1.state[0] ));
 sky130_fd_sc_hd__conb_1 _4369__41 (.LO(net41));
 sky130_fd_sc_hd__dfrtp_4 _4370_ (.CLK(clknet_leaf_17_clk),
    .D(_0001_),
    .RESET_B(net38),
    .Q(\em0.u1.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4371_ (.CLK(clknet_leaf_17_clk),
    .D(_0002_),
    .RESET_B(net38),
    .Q(\em0.u1.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4372_ (.CLK(clknet_leaf_17_clk),
    .D(_0000_),
    .RESET_B(net38),
    .Q(\em0.u1.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4373_ (.CLK(clknet_leaf_0_clk),
    .D(\d10.nxt_count[0] ),
    .RESET_B(net23),
    .Q(\d10.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4374_ (.CLK(clknet_leaf_0_clk),
    .D(\d10.nxt_count[1] ),
    .RESET_B(net23),
    .Q(\d10.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4375_ (.CLK(clknet_leaf_0_clk),
    .D(\d10.nxt_count[2] ),
    .RESET_B(net23),
    .Q(\d10.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4376_ (.CLK(clknet_leaf_0_clk),
    .D(\d10.nxt_count[3] ),
    .RESET_B(net23),
    .Q(\d10.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4377_ (.CLK(clknet_leaf_37_clk),
    .D(\d10.nxt_count[4] ),
    .RESET_B(net23),
    .Q(\d10.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4378_ (.CLK(clknet_leaf_37_clk),
    .D(\d10.nxt_count[5] ),
    .RESET_B(net23),
    .Q(\d10.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4379_ (.CLK(clknet_leaf_1_clk),
    .D(\d10.nxt_count[6] ),
    .RESET_B(net23),
    .Q(\d10.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4380_ (.CLK(clknet_leaf_0_clk),
    .D(\d10.nxt_count[7] ),
    .RESET_B(net23),
    .Q(\d10.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4381_ (.CLK(clknet_leaf_0_clk),
    .D(\d10.nxt_count[8] ),
    .RESET_B(net23),
    .Q(\d10.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4382_ (.CLK(clknet_leaf_0_clk),
    .D(net45),
    .RESET_B(net23),
    .Q(\d10.count[9] ));
 sky130_fd_sc_hd__conb_1 _4382__45 (.LO(net45));
 sky130_fd_sc_hd__dfrtp_1 _4383_ (.CLK(clknet_leaf_5_clk),
    .D(_0072_),
    .RESET_B(net26),
    .Q(\d1.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4384_ (.CLK(clknet_leaf_5_clk),
    .D(_0073_),
    .RESET_B(net26),
    .Q(\d1.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4385_ (.CLK(clknet_leaf_4_clk),
    .D(_0074_),
    .RESET_B(net26),
    .Q(\d1.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4386_ (.CLK(clknet_leaf_4_clk),
    .D(_0075_),
    .RESET_B(net26),
    .Q(\d1.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4387_ (.CLK(clknet_leaf_4_clk),
    .D(_0076_),
    .RESET_B(net26),
    .Q(\d1.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4388_ (.CLK(clknet_leaf_4_clk),
    .D(_0077_),
    .RESET_B(net26),
    .Q(\d1.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4389_ (.CLK(clknet_leaf_4_clk),
    .D(_0078_),
    .RESET_B(net27),
    .Q(\d1.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4390_ (.CLK(clknet_leaf_5_clk),
    .D(_0079_),
    .RESET_B(net27),
    .Q(\d1.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4391_ (.CLK(clknet_leaf_1_clk),
    .D(\d11.nxt_count[0] ),
    .RESET_B(net23),
    .Q(\d11.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4392_ (.CLK(clknet_leaf_2_clk),
    .D(\d11.nxt_count[1] ),
    .RESET_B(net23),
    .Q(\d11.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4393_ (.CLK(clknet_leaf_37_clk),
    .D(\d11.nxt_count[2] ),
    .RESET_B(net23),
    .Q(\d11.count[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4394_ (.CLK(clknet_leaf_34_clk),
    .D(\d11.nxt_count[3] ),
    .RESET_B(net25),
    .Q(\d11.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4395_ (.CLK(clknet_leaf_34_clk),
    .D(\d11.nxt_count[4] ),
    .RESET_B(net34),
    .Q(\d11.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4396_ (.CLK(clknet_leaf_34_clk),
    .D(\d11.nxt_count[5] ),
    .RESET_B(net34),
    .Q(\d11.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4397_ (.CLK(clknet_leaf_2_clk),
    .D(\d11.nxt_count[6] ),
    .RESET_B(net26),
    .Q(\d11.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4398_ (.CLK(clknet_leaf_2_clk),
    .D(\d11.nxt_count[7] ),
    .RESET_B(net26),
    .Q(\d11.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4399_ (.CLK(clknet_leaf_2_clk),
    .D(\d11.nxt_count[8] ),
    .RESET_B(net26),
    .Q(\d11.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4400_ (.CLK(clknet_leaf_2_clk),
    .D(net44),
    .RESET_B(net26),
    .Q(\d11.count[9] ));
 sky130_fd_sc_hd__conb_1 _4400__44 (.LO(net44));
 sky130_fd_sc_hd__dfrtp_4 _4401_ (.CLK(clknet_leaf_10_clk),
    .D(_0080_),
    .RESET_B(net36),
    .Q(\d10.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4402_ (.CLK(clknet_leaf_10_clk),
    .D(_0081_),
    .RESET_B(net37),
    .Q(\d10.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4403_ (.CLK(clknet_leaf_10_clk),
    .D(_0082_),
    .RESET_B(net37),
    .Q(\d10.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4404_ (.CLK(clknet_leaf_11_clk),
    .D(_0083_),
    .RESET_B(net37),
    .Q(\d10.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4405_ (.CLK(clknet_leaf_11_clk),
    .D(_0084_),
    .RESET_B(net37),
    .Q(\d10.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4406_ (.CLK(clknet_leaf_11_clk),
    .D(_0085_),
    .RESET_B(net40),
    .Q(\d10.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4407_ (.CLK(clknet_leaf_13_clk),
    .D(_0086_),
    .RESET_B(net40),
    .Q(\d10.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4408_ (.CLK(clknet_leaf_10_clk),
    .D(_0087_),
    .RESET_B(net37),
    .Q(\d10.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4409_ (.CLK(clknet_leaf_38_clk),
    .D(\d12.nxt_count[0] ),
    .RESET_B(net22),
    .Q(\d12.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4410_ (.CLK(clknet_leaf_0_clk),
    .D(\d12.nxt_count[1] ),
    .RESET_B(net22),
    .Q(\d12.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4411_ (.CLK(clknet_leaf_0_clk),
    .D(\d12.nxt_count[2] ),
    .RESET_B(net22),
    .Q(\d12.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4412_ (.CLK(clknet_leaf_0_clk),
    .D(\d12.nxt_count[3] ),
    .RESET_B(net22),
    .Q(\d12.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4413_ (.CLK(clknet_leaf_38_clk),
    .D(\d12.nxt_count[4] ),
    .RESET_B(net22),
    .Q(\d12.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4414_ (.CLK(clknet_leaf_38_clk),
    .D(\d12.nxt_count[5] ),
    .RESET_B(net22),
    .Q(\d12.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4415_ (.CLK(clknet_leaf_38_clk),
    .D(\d12.nxt_count[6] ),
    .RESET_B(net22),
    .Q(\d12.count[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4416_ (.CLK(clknet_leaf_38_clk),
    .D(\d12.nxt_count[7] ),
    .RESET_B(net22),
    .Q(\d12.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4417_ (.CLK(clknet_leaf_38_clk),
    .D(\d12.nxt_count[8] ),
    .RESET_B(net22),
    .Q(\d12.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4418_ (.CLK(clknet_leaf_38_clk),
    .D(net43),
    .RESET_B(net22),
    .Q(\d12.count[9] ));
 sky130_fd_sc_hd__conb_1 _4418__43 (.LO(net43));
 sky130_fd_sc_hd__dfrtp_2 _4419_ (.CLK(clknet_leaf_9_clk),
    .D(_0088_),
    .RESET_B(net36),
    .Q(\d11.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4420_ (.CLK(clknet_leaf_9_clk),
    .D(_0089_),
    .RESET_B(net36),
    .Q(\d11.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4421_ (.CLK(clknet_leaf_9_clk),
    .D(_0090_),
    .RESET_B(net36),
    .Q(\d11.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4422_ (.CLK(clknet_leaf_9_clk),
    .D(_0091_),
    .RESET_B(net36),
    .Q(\d11.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4423_ (.CLK(clknet_leaf_9_clk),
    .D(_0092_),
    .RESET_B(net37),
    .Q(\d11.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4424_ (.CLK(clknet_leaf_9_clk),
    .D(_0093_),
    .RESET_B(net36),
    .Q(\d11.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4425_ (.CLK(clknet_leaf_10_clk),
    .D(_0094_),
    .RESET_B(net37),
    .Q(\d11.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4426_ (.CLK(clknet_leaf_5_clk),
    .D(_0095_),
    .RESET_B(net26),
    .Q(\d11.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4427_ (.CLK(clknet_leaf_20_clk),
    .D(_0096_),
    .RESET_B(net39),
    .Q(\em0.u1.R[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4428_ (.CLK(clknet_leaf_20_clk),
    .D(_0097_),
    .RESET_B(net38),
    .Q(\em0.u1.R[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4429_ (.CLK(clknet_leaf_20_clk),
    .D(_0098_),
    .RESET_B(net38),
    .Q(\em0.u1.R[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4430_ (.CLK(clknet_leaf_20_clk),
    .D(net97),
    .RESET_B(net38),
    .Q(\em0.u1.R[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4431_ (.CLK(clknet_leaf_20_clk),
    .D(_0100_),
    .RESET_B(net38),
    .Q(\em0.u1.R[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4432_ (.CLK(clknet_leaf_17_clk),
    .D(net62),
    .RESET_B(net38),
    .Q(\em0.u1.R[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4433_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0102_),
    .RESET_B(net40),
    .Q(\em0.u1.R[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4434_ (.CLK(clknet_leaf_16_clk),
    .D(net57),
    .RESET_B(net40),
    .Q(\em0.u1.R[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4435_ (.CLK(clknet_leaf_14_clk),
    .D(_0104_),
    .RESET_B(net40),
    .Q(\em0.u1.R[16] ));
 sky130_fd_sc_hd__dfrtp_2 _4436_ (.CLK(clknet_leaf_15_clk),
    .D(_0105_),
    .RESET_B(net40),
    .Q(\em0.u1.R[17] ));
 sky130_fd_sc_hd__dfrtp_2 _4437_ (.CLK(clknet_leaf_15_clk),
    .D(_0106_),
    .RESET_B(net40),
    .Q(\em0.u1.R[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4438_ (.CLK(clknet_leaf_14_clk),
    .D(_0107_),
    .RESET_B(net40),
    .Q(\em0.u1.R[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4439_ (.CLK(clknet_leaf_16_clk),
    .D(_0108_),
    .RESET_B(net16),
    .Q(\em0.u1.R[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4440_ (.CLK(clknet_leaf_16_clk),
    .D(_0109_),
    .RESET_B(net16),
    .Q(\em0.u1.R[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4441_ (.CLK(clknet_leaf_16_clk),
    .D(_0110_),
    .RESET_B(net16),
    .Q(\em0.u1.R[22] ));
 sky130_fd_sc_hd__dfrtp_2 _4442_ (.CLK(clknet_leaf_21_clk),
    .D(net72),
    .RESET_B(net32),
    .Q(\d13.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4443_ (.CLK(clknet_leaf_21_clk),
    .D(\d13.nxt_count[1] ),
    .RESET_B(net32),
    .Q(\d13.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4444_ (.CLK(clknet_leaf_31_clk),
    .D(\d13.nxt_count[2] ),
    .RESET_B(net31),
    .Q(\d13.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4445_ (.CLK(clknet_leaf_31_clk),
    .D(\d13.nxt_count[3] ),
    .RESET_B(net31),
    .Q(\d13.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4446_ (.CLK(clknet_leaf_30_clk),
    .D(\d13.nxt_count[4] ),
    .RESET_B(net29),
    .Q(\d13.count[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4447_ (.CLK(clknet_leaf_30_clk),
    .D(\d13.nxt_count[5] ),
    .RESET_B(net29),
    .Q(\d13.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4448_ (.CLK(clknet_leaf_27_clk),
    .D(\d13.nxt_count[6] ),
    .RESET_B(net29),
    .Q(\d13.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4449_ (.CLK(clknet_leaf_27_clk),
    .D(\d13.nxt_count[7] ),
    .RESET_B(net29),
    .Q(\d13.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4450_ (.CLK(clknet_leaf_27_clk),
    .D(\d13.nxt_count[8] ),
    .RESET_B(net30),
    .Q(\d13.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4451_ (.CLK(clknet_leaf_27_clk),
    .D(net42),
    .RESET_B(net28),
    .Q(\d13.count[9] ));
 sky130_fd_sc_hd__conb_1 _4451__42 (.LO(net42));
 sky130_fd_sc_hd__dfrtp_2 _4452_ (.CLK(clknet_leaf_6_clk),
    .D(_0111_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4453_ (.CLK(clknet_leaf_6_clk),
    .D(_0112_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4454_ (.CLK(clknet_leaf_6_clk),
    .D(_0113_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4455_ (.CLK(clknet_leaf_4_clk),
    .D(_0114_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4456_ (.CLK(clknet_leaf_6_clk),
    .D(_0115_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4457_ (.CLK(clknet_leaf_6_clk),
    .D(_0116_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4458_ (.CLK(clknet_leaf_6_clk),
    .D(_0117_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4459_ (.CLK(clknet_leaf_4_clk),
    .D(_0118_),
    .RESET_B(net35),
    .Q(\d12.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4460_ (.CLK(clknet_leaf_18_clk),
    .D(_0119_),
    .RESET_B(net38),
    .Q(\em0.mixed_sample[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4461_ (.CLK(clknet_leaf_17_clk),
    .D(_0120_),
    .RESET_B(net38),
    .Q(\em0.mixed_sample[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4462_ (.CLK(clknet_leaf_19_clk),
    .D(_0121_),
    .RESET_B(net39),
    .Q(\em0.mixed_sample[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4463_ (.CLK(clknet_leaf_19_clk),
    .D(_0122_),
    .RESET_B(net39),
    .Q(\em0.mixed_sample[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4464_ (.CLK(clknet_leaf_19_clk),
    .D(_0123_),
    .RESET_B(net39),
    .Q(\em0.mixed_sample[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4465_ (.CLK(clknet_leaf_22_clk),
    .D(_0124_),
    .RESET_B(net33),
    .Q(\em0.mixed_sample[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4466_ (.CLK(clknet_leaf_22_clk),
    .D(_0125_),
    .RESET_B(net33),
    .Q(\em0.mixed_sample[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4467_ (.CLK(clknet_leaf_23_clk),
    .D(_0126_),
    .RESET_B(net33),
    .Q(\em0.mixed_sample[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4468_ (.CLK(clknet_leaf_17_clk),
    .D(_0127_),
    .RESET_B(net38),
    .Q(\em0.u1.Q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4469_ (.CLK(clknet_leaf_18_clk),
    .D(net93),
    .RESET_B(net38),
    .Q(\em0.u1.Q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4470_ (.CLK(clknet_leaf_18_clk),
    .D(_0129_),
    .RESET_B(net38),
    .Q(\em0.u1.Q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4471_ (.CLK(clknet_leaf_19_clk),
    .D(net79),
    .RESET_B(net39),
    .Q(\em0.u1.Q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4472_ (.CLK(clknet_leaf_19_clk),
    .D(_0131_),
    .RESET_B(net39),
    .Q(\em0.u1.Q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4473_ (.CLK(clknet_leaf_23_clk),
    .D(net59),
    .RESET_B(net33),
    .Q(\em0.u1.Q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4474_ (.CLK(clknet_leaf_23_clk),
    .D(net89),
    .RESET_B(net33),
    .Q(\em0.u1.Q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4475_ (.CLK(clknet_leaf_23_clk),
    .D(net64),
    .RESET_B(net33),
    .Q(\em0.u1.Q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4476_ (.CLK(clknet_leaf_18_clk),
    .D(_0135_),
    .RESET_B(net16),
    .Q(\em0.u1.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4477_ (.CLK(clknet_leaf_17_clk),
    .D(net107),
    .RESET_B(net39),
    .Q(\em0.u1.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4478_ (.CLK(clknet_leaf_17_clk),
    .D(_0137_),
    .RESET_B(net39),
    .Q(\em0.u1.count[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4479_ (.CLK(clknet_leaf_8_clk),
    .D(_0138_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4480_ (.CLK(clknet_leaf_8_clk),
    .D(_0139_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4481_ (.CLK(clknet_leaf_8_clk),
    .D(_0140_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4482_ (.CLK(clknet_leaf_8_clk),
    .D(_0141_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4483_ (.CLK(clknet_leaf_8_clk),
    .D(_0142_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4484_ (.CLK(clknet_leaf_8_clk),
    .D(_0143_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4485_ (.CLK(clknet_leaf_8_clk),
    .D(_0144_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4486_ (.CLK(clknet_leaf_8_clk),
    .D(_0145_),
    .RESET_B(net36),
    .Q(\d9.saw_temp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4487_ (.CLK(clknet_leaf_25_clk),
    .D(\p0.pwm ),
    .RESET_B(net34),
    .Q(net17));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_6 fanout22 (.A(net34),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_8 fanout23 (.A(net34),
    .X(net23));
 sky130_fd_sc_hd__buf_6 fanout24 (.A(net34),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net34),
    .X(net25));
 sky130_fd_sc_hd__buf_6 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_6 fanout27 (.A(net34),
    .X(net27));
 sky130_fd_sc_hd__buf_6 fanout28 (.A(net30),
    .X(net28));
 sky130_fd_sc_hd__buf_4 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(net34),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 fanout31 (.A(net33),
    .X(net31));
 sky130_fd_sc_hd__buf_6 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_4 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_8 fanout34 (.A(net16),
    .X(net34));
 sky130_fd_sc_hd__buf_6 fanout35 (.A(net37),
    .X(net35));
 sky130_fd_sc_hd__buf_6 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_4 fanout37 (.A(net16),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_6 fanout39 (.A(net16),
    .X(net39));
 sky130_fd_sc_hd__buf_6 fanout40 (.A(net16),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\m0.synco.delay ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\em0.u1.R[12] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\d9.saw_temp[1] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\d4.saw_temp[0] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\d13.saw_temp[1] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\d12.saw_temp[1] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\d7.saw_temp[5] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\d9.saw_temp[2] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\d4.count[4] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\em0.u1.D[11] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\d11.count[6] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\d3.saw_temp[1] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0101_),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\d4.saw_temp[4] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\d5.count[6] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_1903_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\d8.saw_temp[3] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\d9.saw_temp[4] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_1704_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\d8.saw_temp[4] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\d6.saw_temp[4] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\d1.saw_temp[3] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\d2.saw_temp[1] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\em0.u1.Q[7] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\d6.saw_temp[2] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\d1.saw_temp[4] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\d7.saw_temp[4] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\d2.saw_temp[3] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\d11.count[5] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\d12.saw_temp[4] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\d1.saw_temp[1] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\d1.saw_temp[2] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\em0.mixed_sample[1] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\d7.saw_temp[2] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0134_),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\d7.count[4] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\d4.saw_temp[2] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\d10.saw_temp[7] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\d3.count[5] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\d12.count[8] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\d2.count[7] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\em0.mixed_sample[6] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\em0.mixed_sample[7] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\d7.saw_temp[0] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\em0.mixed_sample[0] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\d11.count[0] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\d13.saw_temp[0] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\d7.saw_temp[7] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\d10.count[6] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\d5.count[5] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_1901_),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\d5.saw_temp[0] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\d2.count[5] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\d10.saw_temp[2] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0584_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\d2.count[4] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\em0.u1.R[8] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\d12.saw_temp[0] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\d6.saw_temp[7] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\d3.count[3] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\d9.saw_temp[7] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\d9.count[5] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\d6.saw_temp[0] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\d2.saw_temp[2] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\em0.u1.Q[5] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\d3.count[7] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\d13.saw_temp[4] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\em0.u1.R[21] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\d12.saw_temp[2] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\d4.count[6] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\d1.count[3] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\d10.count[5] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\d13.count[4] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\d8.saw_temp[2] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0544_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\d2.saw_temp[4] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\d13.saw_temp[2] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\m0.edgy.delay ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\d8.count[0] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\d5.saw_temp[2] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0485_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\d10.count[4] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\d3.saw_temp[2] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\p0.count[4] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\p0.nxt_count[4] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\d8.count[6] ),
    .X(net227));
 sky130_fd_sc_hd__buf_1 hold177 (.A(\d5.count[9] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\d5.saw_temp[4] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\d1.count[5] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\d8.nxt_count[0] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\d11.saw_temp[4] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\d3.count[4] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\d10.saw_temp[0] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\d11.count[4] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\d2.saw_temp[0] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\d8.count[4] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\d7.count[5] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\d1.count[6] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\d3.saw_temp[0] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\d9.count[6] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\d6.count[0] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\d3.saw_temp[5] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\d9.saw_temp[0] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\d3.saw_temp[3] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\em0.u1.D[10] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\em0.u1.state[2] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\d4.count[7] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\d11.saw_temp[0] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\d2.count[3] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\d3.count[6] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\d1.count[4] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\m0.syncy.delay ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\d13.count[0] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\em0.u1.Q[4] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\d10.saw_temp[5] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\d13.nxt_count[0] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\d3.count[0] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\d4.count[0] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\d4.nxt_count[0] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\d9.count[0] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\d9.nxt_count[0] ),
    .X(net77));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold27 (.A(\em0.u1.Q[2] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0130_),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\d1.count[0] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\m0.edgy.in ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\p0.count[7] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\d5.count[0] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\d5.nxt_count[0] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\d12.count[0] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\d7.count[0] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\d10.count[0] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\d3.count[8] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\em0.u1.Q[6] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0133_),
    .X(net89));
 sky130_fd_sc_hd__buf_1 hold39 (.A(\p0.count[0] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\m0.edgo.in ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\em0.u1.R[20] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\em0.u1.Q[1] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0128_),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\d7.saw_temp[6] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\em0.u1.R[9] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\em0.u1.R[10] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0099_),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\d2.count[8] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\d11.saw_temp[6] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\d12.count[4] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\em0.u1.R[14] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\d12.saw_temp[6] ),
    .X(net101));
 sky130_fd_sc_hd__buf_1 hold51 (.A(\em0.u1.count[0] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\em0.u1.Q[3] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\d4.saw_temp[3] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\d5.saw_temp[6] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\em0.u1.count[1] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0136_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\d1.saw_temp[6] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\d1.count[8] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\d1.nxt_count[8] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0103_),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\d2.count[0] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\d6.saw_temp[6] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\em0.mixed_sample[7] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\d3.saw_temp[6] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\d13.saw_temp[6] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\em0.u1.D[9] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\d10.saw_temp[6] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\d5.saw_temp[1] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\d9.saw_temp[6] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\d10.saw_temp[3] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\em0.u1.Q[4] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\p0.count[5] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0293_),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\d2.saw_temp[6] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\d10.saw_temp[1] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\d9.saw_temp[3] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\p0.count[2] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0288_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\em0.u1.R[22] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\d8.saw_temp[1] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\d4.saw_temp[6] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0132_),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\em0.u1.Q[0] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\p0.count[3] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\d8.saw_temp[6] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\p0.count[1] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\d11.saw_temp[1] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\d11.saw_temp[3] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\d12.count[6] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\d6.count[4] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\d6.saw_temp[1] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\d6.saw_temp[5] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\em0.u1.count[2] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\d4.count[5] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\d10.saw_temp[5] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\d12.saw_temp[5] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\d10.saw_temp[4] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\d13.saw_temp[3] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\d6.saw_temp[3] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\em0.u1.D[8] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\d6.count[6] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\d12.saw_temp[3] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\d3.saw_temp[4] ),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(modes),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(pb[4]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(pb[5]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(pb[6]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(pb[7]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(pb[8]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(pb[9]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(reset),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(octaves),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(pb[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(pb[10]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(pb[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(pb[12]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(pb[1]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(pb[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(pb[3]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(PWM_o));
 sky130_fd_sc_hd__clkbuf_2 wire18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire19 (.A(_0580_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 wire21 (.A(_1076_),
    .X(net21));
endmodule

