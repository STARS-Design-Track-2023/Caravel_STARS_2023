* NGSPICE file created from stopwatch.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt stopwatch clk nrst out_0[0] out_0[1] out_0[2] out_0[3] out_0[4] out_0[5] out_0[6]
+ out_1[0] out_1[1] out_1[2] out_1[3] out_1[4] out_1[5] out_1[6] out_2[0] out_2[1]
+ out_2[2] out_2[3] out_2[4] out_2[5] out_2[6] out_3[0] out_3[1] out_3[2] out_3[3]
+ out_3[4] out_3[5] out_3[6] pb_0 pb_1 time_done vccd1 vssd1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0985_ _0353_ _0440_ _0327_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0770_ _0264_ _0265_ _0212_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0968_ TIM.cnt\[5\] _0423_ _0360_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0899_ TIM.cnt\[9\] _0327_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0822_ _0071_ MEM.mem1\[6\] _0069_ _0310_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__o211a_1
X_0684_ CTR.time_out\[2\] _0233_ _0237_ net50 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0753_ CTR.time_out\[6\] _0253_ _0254_ net112 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[6\]
+ sky130_fd_sc_hd__a22o_1
X_1098_ clknet_4_0_0_clk MEM.next_mem4\[7\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1021_ clknet_4_5_0_clk net3 net37 vssd1 vssd1 vccd1 vccd1 e2.intermediate sky130_fd_sc_hd__dfrtp_1
X_0805_ _0290_ _0293_ _0125_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0598_ net115 _0165_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__xnor2_1
X_0736_ CTR.time_out\[5\] _0249_ _0250_ net70 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[5\]
+ sky130_fd_sc_hd__a22o_1
X_0667_ _0215_ _0221_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold74 CLKDIV.count\[17\] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 MEM.mem2\[1\] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 MEM.mem5\[7\] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 MEM.mem4\[3\] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 MEM.mem5\[11\] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 _0138_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold96 TIM.cnt\[1\] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0521_ _0072_ _0070_ MEM.mem3\[7\] _0073_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__and4bb_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _0388_ _0390_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0719_ _0189_ _0246_ _0247_ net77 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[3\] sky130_fd_sc_hd__a22o_1
XFILLER_0_50_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 out_2[2] sky130_fd_sc_hd__clkbuf_4
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 out_3[6] sky130_fd_sc_hd__clkbuf_4
Xoutput7 net7 vssd1 vssd1 vccd1 vccd1 out_0[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0504_ _0094_ _0095_ _0096_ _0097_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__or4_2
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0984_ TIM.cnt\[0\] CLKDIV.secpulse vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0967_ TIM.cnt\[4\] _0358_ _0406_ _0428_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__a22o_1
X_0898_ net136 _0362_ _0364_ _0373_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0752_ CTR.time_out\[5\] _0253_ _0254_ net75 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0821_ MEM.mem4\[6\] _0078_ _0079_ MEM.mem3\[6\] _0309_ vssd1 vssd1 vccd1 vccd1 _0310_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0683_ _0200_ _0233_ _0237_ net87 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[1\] sky130_fd_sc_hd__a22o_1
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1097_ clknet_4_1_0_clk MEM.next_mem4\[6\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1020_ clknet_4_5_0_clk net44 net38 vssd1 vssd1 vccd1 vccd1 e2.edge_d sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_0735_ CTR.time_out\[4\] _0249_ _0250_ net107 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[4\]
+ sky130_fd_sc_hd__a22o_1
X_0804_ _0111_ _0292_ _0133_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0597_ _0167_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__clkbuf_1
X_0666_ _0226_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold75 CLKDIV.count\[11\] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 CLKDIV.count\[14\] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 MEM.mem2\[5\] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 MEM.mem2\[10\] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 TIM.cnt\[9\] vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 MEM.mem5\[9\] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 MEM.mem4\[0\] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0520_ _0092_ _0093_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1003_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0718_ CTR.time_out\[2\] _0246_ _0247_ net76 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[2\]
+ sky130_fd_sc_hd__a22o_1
X_0649_ _0069_ _0193_ _0194_ _0195_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput8 net8 vssd1 vssd1 vccd1 vccd1 out_0[4] sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 out_2[3] sky130_fd_sc_hd__buf_2
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 time_done sky130_fd_sc_hd__buf_2
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 out_0[6] sky130_fd_sc_hd__buf_2
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0503_ _0072_ _0073_ MEM.mem5\[10\] _0070_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__a31o_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0983_ _0071_ _0340_ _0076_ _0439_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0897_ _0371_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__nor2_1
X_0966_ _0360_ _0424_ _0425_ _0427_ _0327_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__o32a_1
XFILLER_0_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0751_ CTR.time_out\[4\] _0253_ _0254_ net89 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[4\]
+ sky130_fd_sc_hd__a22o_1
X_0820_ MEM.mem5\[6\] _0075_ _0076_ MEM.mem2\[6\] _0070_ vssd1 vssd1 vccd1 vccd1 _0309_
+ sky130_fd_sc_hd__a221o_1
X_0682_ _0229_ _0233_ _0237_ net57 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1096_ clknet_4_6_0_clk MEM.next_mem4\[5\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0949_ _0350_ _0412_ _0348_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0665_ _0218_ _0220_ _0225_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__or3b_2
X_0803_ _0127_ _0290_ _0291_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0734_ _0189_ _0249_ _0250_ net104 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[3\] sky130_fd_sc_hd__a22o_1
X_0596_ _0165_ _0166_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1079_ clknet_4_6_0_clk MEM.next_mem5\[0\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold65 _0162_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 MEM.mem2\[8\] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 MEM.mem3\[10\] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 TIM.cnt\[10\] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 MEM.mem1\[9\] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net32 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 MEM.mem3\[6\] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 MEM.mem5\[3\] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ _0200_ _0229_ CTR.time_out\[2\] CLKDIV.secpulse vssd1 vssd1 vccd1 vccd1 _0452_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_44_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0648_ _0196_ _0202_ _0191_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0717_ _0200_ _0246_ _0247_ net92 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[1\] sky130_fd_sc_hd__a22o_1
X_0579_ CLKDIV.count\[10\] _0153_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
Xoutput9 net9 vssd1 vssd1 vccd1 vccd1 out_0[5] sky130_fd_sc_hd__clkbuf_4
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 out_2[4] sky130_fd_sc_hd__clkbuf_4
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 out_1[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0502_ _0073_ MEM.raddr\[2\] MEM.mem4\[10\] _0072_ vssd1 vssd1 vccd1 vccd1 _0096_
+ sky130_fd_sc_hd__and4bb_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0982_ _0433_ _0436_ _0242_ _0438_ _0070_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0896_ _0366_ _0368_ _0369_ _0370_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a211oi_1
X_0965_ _0352_ _0426_ _0348_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0750_ _0189_ _0253_ _0254_ net95 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[3\] sky130_fd_sc_hd__a22o_1
X_0681_ _0233_ _0236_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__nor2_4
X_1095_ clknet_4_4_0_clk MEM.next_mem4\[4\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0948_ TIM.cnt\[1\] TIM.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0879_ _0085_ _0236_ _0330_ _0082_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0802_ _0103_ _0111_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__or2_1
X_0664_ net12 _0219_ _0224_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__a21o_1
X_0733_ CTR.time_out\[2\] _0249_ _0250_ net63 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0595_ CLKDIV.count\[16\] _0163_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__or2_1
X_1078_ clknet_4_7_0_clk _0056_ net41 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[5\] sky130_fd_sc_hd__dfrtp_4
Xhold22 MEM.mem4\[2\] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 MEM.mem1\[7\] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 CTR.minutes vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 MEM.mem2\[4\] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 MEM.mem4\[6\] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 TIM.cnt\[5\] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 MEM.mem4\[4\] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 MEM.mem4\[1\] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _0200_ _0229_ CLKDIV.secpulse CTR.time_out\[2\] vssd1 vssd1 vccd1 vccd1 _0451_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0578_ CLKDIV.count\[10\] _0153_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__or2_1
X_0647_ _0183_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0716_ _0229_ _0246_ _0247_ net80 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 out_1[1] sky130_fd_sc_hd__buf_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 out_2[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0501_ _0072_ _0073_ MEM.mem2\[10\] vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__nor3b_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0981_ _0340_ _0437_ _0431_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0964_ TIM.cnt\[4\] _0351_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0895_ _0369_ _0370_ _0366_ _0368_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0680_ _0235_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__buf_8
XFILLER_0_19_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1094_ clknet_4_1_0_clk MEM.next_mem4\[3\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0947_ _0406_ _0410_ _0411_ _0358_ net137 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0878_ TIM.cnt\[7\] TIM.cnt\[6\] _0354_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__or4_1
X_0801_ _0124_ _0122_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0594_ CLKDIV.count\[16\] _0163_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__nand2_1
X_0663_ _0217_ _0223_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__and2_1
X_0732_ _0200_ _0249_ _0250_ net85 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[1\] sky130_fd_sc_hd__a22o_1
XFILLER_0_47_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1077_ clknet_4_13_0_clk _0055_ net38 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[4\] sky130_fd_sc_hd__dfrtp_4
Xhold56 MEM.next_mem2\[4\] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 MEM.mem5\[5\] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 MEM.mem5\[2\] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 MEM.mem1\[10\] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 MEM.mem4\[11\] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 CLKDIV.count\[8\] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 CTR.time_out\[11\] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 MEM.mem2\[9\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1000_ _0389_ _0449_ _0450_ _0390_ _0200_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0715_ _0236_ _0246_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__nor2_4
X_0577_ net113 _0151_ _0154_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__o21a_1
X_0646_ _0183_ _0191_ _0203_ _0208_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__a31oi_4
X_1129_ clknet_4_12_0_clk MEM.next_mem1\[2\] net39 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 out_2[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 out_1[2] sky130_fd_sc_hd__clkbuf_4
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0500_ _0072_ MEM.raddr\[2\] MEM.mem3\[10\] _0073_ vssd1 vssd1 vccd1 vccd1 _0094_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0629_ MEM.mem5\[2\] _0075_ _0076_ MEM.mem2\[2\] _0070_ vssd1 vssd1 vccd1 vccd1 _0192_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0980_ _0230_ _0075_ _0076_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0894_ TIM.cnt\[8\] _0327_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0963_ TIM.cnt\[3\] _0415_ TIM.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1093_ clknet_4_6_0_clk MEM.next_mem4\[2\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0877_ TIM.cnt\[9\] TIM.cnt\[8\] TIM.cnt\[11\] TIM.cnt\[10\] vssd1 vssd1 vccd1 vccd1
+ _0355_ sky130_fd_sc_hd__or4_1
X_0946_ TIM.cnt\[1\] TIM.cnt\[5\] _0084_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0800_ _0273_ _0289_ _0287_ _0285_ vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__a211o_1
X_0731_ _0229_ _0249_ _0250_ net72 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[0\] sky130_fd_sc_hd__a22o_1
X_0593_ net109 _0161_ _0164_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__o21a_1
X_0662_ _0191_ _0212_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1076_ clknet_4_13_0_clk _0054_ net39 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0929_ CTR.time_out\[7\] CTR.time_out\[6\] CTR.time_out\[8\] _0396_ vssd1 vssd1 vccd1
+ vccd1 _0398_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold68 CLKDIV.count\[15\] vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _0152_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 MEM.mem1\[1\] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 MEM.mem3\[2\] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 MEM.mem3\[4\] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 MEM.mem3\[7\] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 MEM.mem2\[11\] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0714_ _0245_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__buf_4
X_0645_ _0069_ _0205_ _0206_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a31o_2
X_0576_ _0024_ _0153_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__nor2_1
X_1128_ clknet_4_12_0_clk MEM.next_mem1\[1\] net39 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1059_ clknet_4_2_0_clk _0037_ net36 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 out_1[3] sky130_fd_sc_hd__clkbuf_4
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 out_3[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0628_ _0069_ _0187_ _0188_ _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__a31o_4
X_0559_ CLKDIV.count\[4\] _0140_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0893_ TIM.cnt\[8\] _0327_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nor2_1
X_0962_ _0423_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1092_ clknet_4_12_0_clk MEM.next_mem4\[1\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0876_ _0327_ _0353_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__nand2_2
X_0945_ _0360_ _0408_ _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0730_ _0236_ _0249_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__nor2_4
X_0661_ _0222_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_0592_ _0024_ _0163_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1075_ clknet_4_14_0_clk _0053_ net39 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[2\] sky130_fd_sc_hd__dfrtp_4
X_0928_ CTR.time_out\[7\] CTR.time_out\[6\] _0396_ CTR.time_out\[8\] vssd1 vssd1 vccd1
+ vccd1 _0397_ sky130_fd_sc_hd__a31o_1
X_0859_ _0328_ _0325_ _0338_ _0339_ vssd1 vssd1 vccd1 vccd1 FSM.next_state\[1\] sky130_fd_sc_hd__a211o_1
Xhold69 MEM.mem5\[8\] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 MEM.mem5\[10\] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 MEM.mem3\[11\] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 MEM.mem1\[6\] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 MEM.mem3\[3\] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 MEM.mem2\[0\] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0713_ MEM.addr\[0\] _0241_ _0230_ _0242_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__and4_1
X_0644_ TIM.cnt\[5\] _0085_ net34 CTR.time_out\[5\] vssd1 vssd1 vccd1 vccd1 _0207_
+ sky130_fd_sc_hd__a22o_1
X_0575_ CLKDIV.count\[9\] _0151_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__and2_1
X_1058_ clknet_4_2_0_clk _0036_ net36 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[10\] sky130_fd_sc_hd__dfrtp_4
X_1127_ clknet_4_12_0_clk MEM.next_mem1\[0\] net39 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 out_1[4] sky130_fd_sc_hd__clkbuf_4
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 out_3[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0558_ _0140_ _0141_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0627_ TIM.cnt\[3\] _0085_ net34 _0189_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__a22o_1
X_0489_ FSM.state\[2\] FSM.state\[1\] _0066_ FSM.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _0083_ sky130_fd_sc_hd__or4b_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0961_ TIM.cnt\[3\] TIM.cnt\[4\] _0415_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__or3_1
X_0892_ _0364_ _0367_ _0368_ _0362_ net134 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1091_ clknet_4_9_0_clk MEM.next_mem4\[0\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0944_ TIM.cnt\[0\] TIM.cnt\[1\] _0407_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0875_ TIM.cnt\[0\] TIM.cnt\[5\] _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0591_ CLKDIV.count\[15\] _0161_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__and2_1
X_0660_ _0215_ _0221_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1074_ clknet_4_15_0_clk _0052_ net39 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0927_ _0236_ _0391_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or2_1
X_0789_ _0224_ _0284_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__nor2_1
X_0858_ _0066_ _0236_ _0322_ _0231_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__a211o_1
Xhold59 MEM.mem2\[2\] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 MEM.mem5\[4\] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 MEM.mem3\[8\] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 MEM.mem4\[8\] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 MEM.mem1\[11\] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0574_ _0151_ net120 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__nor2_1
X_0712_ net98 _0240_ _0244_ CTR.time_out\[11\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[11\]
+ sky130_fd_sc_hd__a22o_1
X_0643_ _0071_ MEM.mem1\[5\] vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__or2_1
X_1126_ clknet_4_3_0_clk MEM.next_mem2\[11\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1057_ clknet_4_2_0_clk _0035_ net36 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 out_1[5] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 out_3[2] sky130_fd_sc_hd__buf_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0557_ net121 _0139_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__nor2_1
X_0626_ CTR.time_out\[3\] vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0488_ FSM.state\[3\] FSM.state\[1\] _0066_ FSM.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _0082_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1109_ clknet_4_1_0_clk MEM.next_mem3\[6\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0609_ net124 _0173_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0960_ _0406_ _0419_ _0422_ _0358_ TIM.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0891_ TIM.cnt\[6\] _0365_ _0366_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout40 net41 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_8
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1090_ clknet_4_3_0_clk MEM.next_mem5\[11\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0874_ TIM.cnt\[4\] _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__or2_1
X_0943_ TIM.cnt\[0\] _0407_ TIM.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0590_ _0161_ net106 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__nor2_1
X_1142_ clknet_4_10_0_clk FSM.next_state\[3\] net40 vssd1 vssd1 vccd1 vccd1 FSM.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_1073_ clknet_4_14_0_clk _0051_ net39 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0926_ _0391_ _0394_ _0395_ _0392_ CTR.time_out\[7\] vssd1 vssd1 vccd1 vccd1 _0033_
+ sky130_fd_sc_hd__a32o_1
X_0857_ _0321_ _0330_ _0336_ _0337_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0788_ _0208_ _0265_ _0283_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a21oi_1
Xhold38 MEM.mem4\[7\] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 MEM.mem3\[9\] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 MEM.mem1\[0\] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 MEM.mem2\[3\] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dlygate4sd3_1
X_0711_ net83 _0240_ _0244_ CTR.time_out\[10\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[10\]
+ sky130_fd_sc_hd__a22o_1
X_0573_ CLKDIV.count\[7\] _0145_ net119 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0642_ MEM.mem4\[5\] _0078_ _0079_ MEM.mem3\[5\] _0204_ vssd1 vssd1 vccd1 vccd1 _0205_
+ sky130_fd_sc_hd__a221o_1
X_1125_ clknet_4_0_0_clk MEM.next_mem2\[10\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1056_ clknet_4_2_0_clk _0034_ net36 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[8\] sky130_fd_sc_hd__dfrtp_4
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 out_3[3] sky130_fd_sc_hd__clkbuf_4
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 out_1[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0909_ _0381_ _0380_ _0379_ _0375_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0625_ _0071_ MEM.mem1\[3\] vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__or2_1
X_0556_ CLKDIV.count\[1\] CLKDIV.count\[0\] CLKDIV.count\[3\] CLKDIV.count\[2\] vssd1
+ vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0487_ _0071_ MEM.mem1\[11\] _0077_ _0080_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__o22a_1
X_1039_ clknet_4_14_0_clk _0007_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1108_ clknet_4_4_0_clk MEM.next_mem3\[5\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0608_ CLKDIV.count\[21\] _0173_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0539_ _0088_ _0102_ _0111_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__or3b_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0890_ _0365_ _0366_ TIM.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout41 net1 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_6
XFILLER_0_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0942_ CLKDIV.secpulse vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
X_0873_ TIM.cnt\[3\] _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1072_ clknet_4_2_0_clk _0050_ net36 vssd1 vssd1 vccd1 vccd1 MEM.addr\[2\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1141_ clknet_4_10_0_clk FSM.next_state\[2\] net40 vssd1 vssd1 vccd1 vccd1 FSM.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_0787_ _0217_ _0279_ _0282_ _0277_ _0262_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__o32a_1
X_0925_ CTR.time_out\[7\] CTR.time_out\[6\] vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__nand2_1
X_0856_ _0067_ _0330_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold28 MEM.mem4\[9\] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 MEM.mem2\[7\] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 MEM.mem3\[0\] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0641_ MEM.mem5\[5\] _0075_ _0076_ MEM.mem2\[5\] _0070_ vssd1 vssd1 vccd1 vccd1 _0204_
+ sky130_fd_sc_hd__a221o_1
X_0710_ net108 _0240_ _0244_ CTR.time_out\[9\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[9\]
+ sky130_fd_sc_hd__a22o_1
X_0572_ CLKDIV.count\[7\] CLKDIV.count\[8\] _0145_ vssd1 vssd1 vccd1 vccd1 _0151_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1124_ clknet_4_3_0_clk MEM.next_mem2\[9\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1055_ clknet_4_1_0_clk _0033_ net35 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 out_2[0] sky130_fd_sc_hd__clkbuf_4
X_0839_ e2.edge_d e2.sync vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__or2b_2
X_0908_ _0375_ _0379_ _0380_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o211ai_2
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 out_3[4] sky130_fd_sc_hd__clkbuf_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ MEM.mem3\[3\] _0079_ _0185_ _0186_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__a211o_1
X_0555_ net126 _0139_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__nor2_1
X_0486_ MEM.mem4\[11\] _0078_ net33 MEM.mem3\[11\] vssd1 vssd1 vccd1 vccd1 _0080_
+ sky130_fd_sc_hd__a22o_1
X_1038_ clknet_4_13_0_clk _0006_ net38 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1107_ clknet_4_4_0_clk MEM.next_mem3\[4\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0607_ _0024_ _0172_ _0173_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__nor3_1
X_0538_ _0126_ _0128_ net26 vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__o21ai_1
X_0469_ _0060_ _0061_ _0062_ _0063_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0941_ _0236_ _0358_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0872_ TIM.cnt\[1\] TIM.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1071_ clknet_4_2_0_clk _0049_ net36 vssd1 vssd1 vccd1 vccd1 MEM.addr\[1\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1140_ clknet_4_8_0_clk FSM.next_state\[1\] net40 vssd1 vssd1 vccd1 vccd1 FSM.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0924_ CTR.time_out\[7\] CTR.time_out\[6\] vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or2_1
X_0786_ _0208_ _0280_ _0281_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0855_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
Xhold18 MEM.mem3\[5\] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 MEM.mem4\[5\] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0571_ _0150_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
X_0640_ _0196_ _0202_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1123_ clknet_4_0_0_clk MEM.next_mem2\[8\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1054_ clknet_4_1_0_clk _0032_ net35 vssd1 vssd1 vccd1 vccd1 CTR.time_out\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0907_ TIM.cnt\[10\] _0327_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__nand2_2
X_0769_ _0210_ _0211_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nor2_1
X_0838_ _0299_ _0320_ _0316_ _0319_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__o2bb2a_2
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 out_2[1] sky130_fd_sc_hd__clkbuf_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0554_ CLKDIV.count\[1\] CLKDIV.count\[0\] CLKDIV.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _0139_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0623_ MEM.mem5\[3\] _0075_ _0076_ MEM.mem2\[3\] vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__a22o_1
X_0485_ _0072_ _0070_ _0073_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__nor3b_2
X_1106_ clknet_4_4_0_clk MEM.next_mem3\[3\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1037_ clknet_4_13_0_clk _0005_ net38 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0606_ CLKDIV.count\[19\] CLKDIV.count\[20\] _0168_ vssd1 vssd1 vccd1 vccd1 _0173_
+ sky130_fd_sc_hd__and3_1
X_0537_ _0113_ _0122_ _0129_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__o21bai_4
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0468_ CLKDIV.count\[17\] CLKDIV.count\[16\] CLKDIV.count\[18\] CLKDIV.count\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__or4b_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ net130 _0403_ _0405_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0871_ _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1070_ clknet_4_2_0_clk _0048_ net36 vssd1 vssd1 vccd1 vccd1 MEM.addr\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0923_ _0393_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__clkbuf_1
X_0854_ _0066_ _0086_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__or2b_2
X_0785_ _0191_ _0203_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold19 MEM.mem5\[0\] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0570_ _0065_ _0148_ _0149_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1122_ clknet_4_1_0_clk MEM.next_mem2\[7\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1053_ clknet_4_12_0_clk _0031_ net39 vssd1 vssd1 vccd1 vccd1 CTR.minutes sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0837_ _0308_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
X_0906_ TIM.cnt\[10\] _0327_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0768_ _0210_ _0211_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__and2_1
X_0699_ MEM.addr\[0\] _0241_ _0230_ _0242_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__and4b_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0553_ CLKDIV.count\[1\] net114 net125 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__a21oi_1
X_0484_ _0073_ _0070_ _0072_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__nor3b_4
X_0622_ _0072_ _0184_ MEM.mem4\[3\] _0070_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__a31o_1
X_1105_ clknet_4_6_0_clk MEM.next_mem3\[2\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1036_ clknet_4_7_0_clk _0004_ net38 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0467_ CLKDIV.count\[21\] CLKDIV.count\[22\] CLKDIV.count\[23\] CLKDIV.count\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__or4bb_1
X_0605_ CLKDIV.count\[19\] _0168_ net131 vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0536_ _0088_ _0101_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1019_ clknet_4_5_0_clk net43 net37 vssd1 vssd1 vccd1 vccd1 e2.sync sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0519_ _0088_ _0102_ _0112_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__nand3_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0870_ TIM.cnt\[1\] TIM.cnt\[3\] TIM.cnt\[2\] TIM.cnt\[4\] TIM.cnt\[5\] vssd1 vssd1
+ vccd1 vccd1 _0348_ sky130_fd_sc_hd__a41o_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ _0200_ _0229_ CLKDIV.secpulse vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0922_ _0391_ _0392_ CTR.time_out\[6\] vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__mux2_1
X_0853_ _0334_ vssd1 vssd1 vccd1 vccd1 FSM.next_state\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0784_ _0191_ _0203_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__nand2_1
Xinput1 nrst vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1052_ clknet_4_10_0_clk _0030_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[11\] sky130_fd_sc_hd__dfrtp_2
X_1121_ clknet_4_1_0_clk MEM.next_mem2\[6\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0767_ _0196_ net12 _0262_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__a21o_1
X_0836_ _0297_ _0316_ _0313_ _0308_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__a211o_1
X_0905_ _0374_ _0376_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0698_ _0066_ _0231_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0621_ _0073_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0552_ _0137_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__clkbuf_1
X_0483_ MEM.mem5\[11\] _0075_ _0076_ MEM.mem2\[11\] _0070_ vssd1 vssd1 vccd1 vccd1
+ _0077_ sky130_fd_sc_hd__a221o_1
X_1035_ clknet_4_7_0_clk _0003_ net38 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1104_ clknet_4_6_0_clk MEM.next_mem3\[1\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0819_ _0300_ _0307_ _0131_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0604_ net102 _0168_ _0171_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0466_ CLKDIV.count\[8\] CLKDIV.count\[11\] CLKDIV.count\[10\] CLKDIV.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__or4bb_1
X_0535_ _0088_ _0127_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1018_ clknet_4_1_0_clk net2 net35 vssd1 vssd1 vccd1 vccd1 e1.intermediate sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0518_ _0103_ _0111_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__nand2_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0998_ _0229_ CLKDIV.secpulse _0200_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ _0236_ _0391_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__nor2_1
X_0783_ _0276_ _0220_ _0223_ _0278_ _0209_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0852_ _0322_ _0325_ _0332_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or4b_1
Xinput2 pb_0 vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1120_ clknet_4_6_0_clk MEM.next_mem2\[5\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1051_ clknet_4_10_0_clk _0029_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0904_ _0364_ _0377_ _0378_ _0362_ net127 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0766_ _0183_ _0191_ _0208_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__o21ai_1
X_0697_ MEM.addr\[1\] vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
X_0835_ _0319_ _0298_ _0312_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0551_ _0058_ _0136_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__and2_1
X_0620_ _0069_ _0180_ _0181_ _0182_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__a31o_2
XFILLER_0_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0482_ _0072_ _0073_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__nor2_4
X_1034_ clknet_4_13_0_clk _0002_ net38 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1103_ clknet_4_6_0_clk MEM.next_mem3\[0\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_0749_ CTR.time_out\[2\] _0253_ _0254_ net86 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[2\]
+ sky130_fd_sc_hd__a22o_1
X_0818_ _0302_ _0306_ net26 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0603_ net102 _0168_ _0065_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__o21ai_1
X_0534_ _0103_ _0113_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__nor2_1
X_0465_ CLKDIV.count\[13\] CLKDIV.count\[14\] CLKDIV.count\[15\] CLKDIV.count\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1017_ clknet_4_8_0_clk net45 net40 vssd1 vssd1 vccd1 vccd1 e1.edge_d sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0517_ TIM.cnt\[8\] _0085_ _0108_ _0109_ _0110_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a221o_2
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout35 net36 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_6
XFILLER_0_51_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0997_ _0389_ _0447_ _0448_ _0390_ _0229_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0920_ CTR.minutes _0336_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__and2_1
X_0782_ _0210_ _0216_ _0277_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0851_ _0067_ _0321_ _0330_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__or3_1
Xinput3 pb_1 vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1050_ clknet_4_10_0_clk _0028_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0834_ _0319_ _0317_ _0315_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__o21a_1
X_0903_ _0374_ _0375_ _0376_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__or3b_1
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0765_ _0259_ _0260_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__and2_1
X_0696_ _0239_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0550_ CLKDIV.count\[1\] CLKDIV.count\[0\] vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0481_ _0074_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__buf_4
X_1102_ clknet_4_3_0_clk MEM.next_mem4\[11\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1033_ clknet_4_7_0_clk _0001_ net38 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0817_ _0129_ _0305_ _0113_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a21oi_1
X_0748_ _0200_ _0253_ _0254_ net103 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[1\] sky130_fd_sc_hd__a22o_1
X_0679_ FSM.state\[1\] _0234_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0602_ _0170_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__clkbuf_1
X_0464_ CLKDIV.count\[3\] CLKDIV.count\[2\] _0057_ _0058_ vssd1 vssd1 vccd1 vccd1
+ _0059_ sky130_fd_sc_hd__or4_1
X_0533_ net31 _0123_ _0125_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1016_ clknet_4_1_0_clk net42 net35 vssd1 vssd1 vccd1 vccd1 e1.sync sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0516_ CTR.time_out\[8\] _0086_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__and2_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout36 net41 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_6
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0996_ _0229_ CLKDIV.secpulse vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0850_ net32 _0327_ _0234_ _0329_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a221o_1
X_0781_ _0191_ _0216_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0979_ _0070_ _0075_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0833_ _0297_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__inv_2
X_0902_ _0374_ _0375_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0764_ _0202_ _0225_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__xnor2_2
X_0695_ MEM.addr\[0\] MEM.addr\[1\] MEM.addr\[2\] _0232_ _0238_ vssd1 vssd1 vccd1
+ vccd1 _0239_ sky130_fd_sc_hd__o41a_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap33 _0079_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0480_ _0072_ _0073_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__and2_1
X_1032_ clknet_4_5_0_clk _0023_ net38 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[9\] sky130_fd_sc_hd__dfrtp_1
X_1101_ clknet_4_0_0_clk MEM.next_mem4\[10\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_0816_ _0121_ _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__nand2_1
X_0747_ _0229_ _0253_ _0254_ net60 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0678_ FSM.state\[2\] FSM.state\[3\] vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0601_ _0168_ _0169_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0463_ CLKDIV.count\[1\] CLKDIV.count\[0\] vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__or2_1
X_0532_ _0102_ _0124_ _0088_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1015_ _0461_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0515_ _0067_ _0068_ _0071_ MEM.mem1\[8\] vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__o2bb2a_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout37 net41 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_6
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0995_ _0229_ CLKDIV.secpulse vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0780_ _0191_ _0212_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0978_ _0072_ _0431_ _0434_ _0435_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0832_ _0318_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_0763_ _0258_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
X_0901_ _0370_ _0372_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0694_ FSM.state\[2\] FSM.state\[3\] FSM.state\[1\] vssd1 vssd1 vccd1 vccd1 _0238_
+ sky130_fd_sc_hd__or3_4
XFILLER_0_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap34 _0086_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_4
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_1031_ clknet_4_5_0_clk _0022_ net41 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[8\] sky130_fd_sc_hd__dfrtp_1
X_1100_ clknet_4_3_0_clk MEM.next_mem4\[9\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_0746_ _0236_ _0253_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__nor2_4
XFILLER_0_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0815_ _0088_ _0111_ _0303_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0677_ _0230_ _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__nor2_8
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0600_ CLKDIV.count\[17\] CLKDIV.count\[16\] _0163_ CLKDIV.count\[18\] vssd1 vssd1
+ vccd1 vccd1 _0169_ sky130_fd_sc_hd__a31o_1
X_0531_ _0111_ _0121_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0462_ CLKDIV.count\[5\] CLKDIV.count\[4\] CLKDIV.count\[6\] CLKDIV.count\[7\] vssd1
+ vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1014_ _0460_ _0458_ CTR.time_out\[5\] vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0729_ _0248_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0514_ _0104_ _0105_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__or4_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout38 net41 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_6
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0994_ MEM.addr\[2\] _0443_ _0446_ _0242_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0977_ _0075_ _0076_ _0232_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__nor3_1
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ TIM.cnt\[9\] _0327_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0831_ _0297_ _0312_ _0298_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__or3b_2
X_0693_ CTR.time_out\[11\] _0233_ _0237_ net78 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[11\]
+ sky130_fd_sc_hd__a22o_1
X_0762_ TIM.cnt\[0\] _0085_ net34 _0229_ _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__a221o_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1030_ clknet_4_5_0_clk _0021_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0814_ _0103_ _0111_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__nor2_1
X_0745_ _0252_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__buf_4
X_0676_ _0066_ _0231_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0530_ _0113_ _0122_ _0103_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1013_ _0335_ _0457_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nor2_1
X_0659_ net12 _0219_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0728_ MEM.addr\[0\] MEM.addr\[1\] _0230_ _0242_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__and4b_1
XFILLER_0_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0513_ _0072_ _0073_ MEM.mem5\[8\] MEM.raddr\[2\] vssd1 vssd1 vccd1 vccd1 _0107_
+ sky130_fd_sc_hd__a31o_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 net41 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_6
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0993_ MEM.addr\[2\] _0251_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0976_ MEM.addr\[1\] _0433_ _0076_ _0075_ _0340_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0830_ _0297_ _0317_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__nand2_1
XFILLER_0_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0692_ CTR.time_out\[10\] _0233_ _0237_ net64 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[10\]
+ sky130_fd_sc_hd__a22o_1
X_0761_ _0071_ MEM.mem1\[0\] _0069_ _0256_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0959_ _0084_ _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0813_ _0088_ _0113_ _0301_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0744_ _0251_ _0230_ _0242_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__and3b_1
X_0675_ FSM.state\[3\] FSM.state\[1\] FSM.state\[2\] vssd1 vssd1 vccd1 vccd1 _0231_
+ sky130_fd_sc_hd__nor3b_4
X_1089_ clknet_4_0_0_clk MEM.next_mem5\[10\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1012_ CTR.time_out\[4\] _0458_ _0459_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0727_ CTR.time_out\[11\] _0246_ _0247_ net66 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[11\]
+ sky130_fd_sc_hd__a22o_1
X_0589_ CLKDIV.count\[13\] _0159_ net105 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0658_ _0208_ _0213_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0512_ _0073_ MEM.raddr\[2\] MEM.mem4\[8\] _0072_ vssd1 vssd1 vccd1 vccd1 _0106_
+ sky130_fd_sc_hd__and4bb_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0992_ MEM.addr\[0\] _0241_ _0242_ _0445_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0975_ _0070_ _0075_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0760_ MEM.mem4\[0\] _0078_ net33 MEM.mem3\[0\] _0255_ vssd1 vssd1 vccd1 vccd1 _0256_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0691_ CTR.time_out\[9\] _0233_ _0237_ net51 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[9\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0889_ TIM.cnt\[7\] _0327_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__nand2_1
X_0958_ _0351_ _0420_ _0348_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0812_ _0112_ _0291_ _0121_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__a21oi_1
X_0743_ MEM.addr\[0\] MEM.addr\[1\] vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0674_ MEM.addr\[2\] vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__inv_2
X_1088_ clknet_4_3_0_clk MEM.next_mem5\[9\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1011_ CTR.time_out\[4\] _0335_ _0387_ _0456_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or4_1
X_0726_ CTR.time_out\[10\] _0246_ _0247_ net84 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[10\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0588_ CLKDIV.count\[13\] CLKDIV.count\[14\] _0159_ vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__and3_1
X_0657_ _0209_ _0214_ _0218_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0511_ _0072_ _0073_ MEM.mem2\[8\] vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0709_ net73 _0240_ _0244_ CTR.time_out\[8\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[8\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ _0443_ _0444_ MEM.addr\[1\] vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0974_ _0070_ MEM.addr\[0\] _0340_ _0075_ _0432_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__a41o_1
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_0690_ CTR.time_out\[8\] _0233_ _0237_ net49 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[8\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0888_ TIM.cnt\[7\] _0327_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__or2_1
X_0957_ TIM.cnt\[3\] _0350_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0673_ CTR.time_out\[0\] vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__buf_4
X_0811_ _0129_ _0122_ _0113_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__and3b_1
X_0742_ CTR.time_out\[11\] _0249_ _0250_ net53 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[11\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1087_ clknet_4_0_0_clk MEM.next_mem5\[8\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1010_ _0389_ _0457_ _0454_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__a21o_1
X_0656_ _0183_ _0191_ _0208_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__o21a_1
X_0725_ CTR.time_out\[9\] _0246_ _0247_ net68 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[9\]
+ sky130_fd_sc_hd__a22o_1
X_0587_ net111 _0159_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1139_ clknet_4_9_0_clk FSM.next_state\[0\] net40 vssd1 vssd1 vccd1 vccd1 FSM.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0510_ _0072_ MEM.raddr\[2\] MEM.mem3\[8\] _0073_ vssd1 vssd1 vccd1 vccd1 _0104_
+ sky130_fd_sc_hd__and4bb_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 e1.intermediate vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0639_ _0198_ _0199_ _0201_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__a21oi_4
X_0708_ net58 _0240_ _0244_ CTR.time_out\[7\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0990_ net135 _0443_ _0444_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0973_ _0231_ _0431_ _0073_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0956_ TIM.cnt\[3\] _0415_ _0418_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0887_ _0236_ _0362_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0810_ _0297_ _0298_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__nor2_1
X_0672_ _0220_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__inv_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0741_ CTR.time_out\[10\] _0249_ _0250_ net81 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[10\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1086_ clknet_4_0_0_clk MEM.next_mem5\[7\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_0939_ CTR.time_out\[11\] _0403_ _0238_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0586_ _0024_ _0159_ _0160_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__nor3b_1
X_0655_ _0191_ _0216_ _0217_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__o21ai_2
X_0724_ CTR.time_out\[8\] _0246_ _0247_ net56 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[8\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1138_ clknet_4_8_0_clk MEM.next_mem1\[11\] net40 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1069_ clknet_4_9_0_clk _0047_ net39 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 e2.intermediate vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0707_ net91 _0240_ _0244_ CTR.time_out\[6\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[6\]
+ sky130_fd_sc_hd__a22o_1
X_0569_ CLKDIV.count\[7\] _0145_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__nand2_1
X_0638_ TIM.cnt\[1\] _0085_ net34 _0200_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ FSM.state\[3\] FSM.state\[1\] vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0886_ _0363_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__clkbuf_1
X_0955_ TIM.cnt\[3\] _0415_ _0360_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0740_ CTR.time_out\[9\] _0249_ _0250_ net69 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[9\]
+ sky130_fd_sc_hd__a22o_1
X_0671_ _0215_ net12 _0220_ _0218_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__a31o_1
X_1085_ clknet_4_1_0_clk MEM.next_mem5\[6\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_0938_ CTR.time_out\[10\] _0401_ _0404_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__o21a_1
X_0869_ TIM.cnt\[6\] _0234_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0723_ CTR.time_out\[7\] _0246_ _0247_ net54 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[7\]
+ sky130_fd_sc_hd__a22o_1
X_0585_ CLKDIV.count\[11\] CLKDIV.count\[10\] _0153_ CLKDIV.count\[12\] vssd1 vssd1
+ vccd1 vccd1 _0160_ sky130_fd_sc_hd__a31o_1
X_0654_ _0208_ _0183_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1137_ clknet_4_10_0_clk MEM.next_mem1\[10\] net40 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1068_ clknet_4_2_0_clk _0046_ net35 vssd1 vssd1 vccd1 vccd1 MEM.raddr\[2\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 e2.sync vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
X_0706_ net94 _0240_ _0244_ CTR.time_out\[5\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0568_ CLKDIV.count\[7\] _0145_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__or2_1
X_0637_ CTR.time_out\[1\] vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_4
X_0499_ TIM.cnt\[9\] _0085_ _0086_ CTR.time_out\[9\] vssd1 vssd1 vccd1 vccd1 _0093_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0971_ net117 _0238_ _0356_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0885_ _0347_ TIM.cnt\[6\] _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__mux2_1
X_0954_ _0354_ _0406_ _0417_ _0358_ net132 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0670_ _0228_ vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_1084_ clknet_4_4_0_clk MEM.next_mem5\[5\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_0799_ _0273_ _0289_ _0285_ _0261_ vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__a211o_1
X_0937_ _0236_ _0403_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nor2_1
X_0868_ _0346_ vssd1 vssd1 vccd1 vccd1 FSM.next_state\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0653_ _0196_ _0202_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0722_ CTR.time_out\[6\] _0246_ _0247_ net62 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[6\]
+ sky130_fd_sc_hd__a22o_1
X_0584_ _0158_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__buf_1
XFILLER_0_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1067_ clknet_4_2_0_clk _0045_ net36 vssd1 vssd1 vccd1 vccd1 MEM.raddr\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1136_ clknet_4_8_0_clk MEM.next_mem1\[9\] net40 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 e1.sync vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dlygate4sd3_1
X_0705_ net96 _0240_ _0244_ CTR.time_out\[4\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[4\]
+ sky130_fd_sc_hd__a22o_1
X_0636_ _0071_ MEM.mem1\[1\] _0069_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__o21a_1
X_0567_ _0147_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__clkbuf_1
X_0498_ _0089_ _0090_ _0091_ _0069_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1119_ clknet_4_4_0_clk net97 net37 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0619_ TIM.cnt\[4\] _0085_ net34 CTR.time_out\[4\] vssd1 vssd1 vccd1 vccd1 _0182_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_0970_ _0406_ _0429_ _0430_ _0358_ net129 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0884_ _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__buf_2
X_0953_ _0084_ _0413_ _0416_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1083_ clknet_4_4_0_clk MEM.next_mem5\[4\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_0936_ CTR.time_out\[10\] CTR.time_out\[9\] _0398_ vssd1 vssd1 vccd1 vccd1 _0403_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0798_ _0259_ _0260_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0867_ _0327_ _0331_ _0345_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0583_ CLKDIV.count\[11\] CLKDIV.count\[10\] CLKDIV.count\[12\] _0153_ vssd1 vssd1
+ vccd1 vccd1 _0158_ sky130_fd_sc_hd__and4_1
X_0652_ _0209_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0721_ CTR.time_out\[5\] _0246_ _0247_ net59 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1066_ clknet_4_2_0_clk _0044_ net36 vssd1 vssd1 vccd1 vccd1 MEM.raddr\[0\] sky130_fd_sc_hd__dfstp_1
X_1135_ clknet_4_8_0_clk MEM.next_mem1\[8\] net40 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_0919_ net118 _0388_ _0390_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 MEM.mem1\[5\] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0566_ _0145_ _0146_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__and2b_1
X_0635_ MEM.mem4\[1\] _0078_ net33 MEM.mem3\[1\] _0197_ vssd1 vssd1 vccd1 vccd1 _0198_
+ sky130_fd_sc_hd__a221o_1
X_0704_ net90 _0240_ _0244_ _0189_ vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[3\] sky130_fd_sc_hd__a22o_1
X_0497_ _0071_ MEM.mem1\[9\] vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1049_ clknet_4_10_0_clk _0027_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[8\] sky130_fd_sc_hd__dfrtp_1
X_1118_ clknet_4_4_0_clk MEM.next_mem2\[3\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0549_ net114 _0024_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__nor2_1
X_0618_ _0071_ MEM.mem1\[4\] vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0952_ _0327_ _0414_ _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0883_ _0359_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1082_ clknet_4_4_0_clk MEM.next_mem5\[3\] net37 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_0935_ CTR.time_out\[9\] _0398_ _0402_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0866_ _0082_ _0321_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0797_ _0260_ _0273_ _0258_ vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0720_ CTR.time_out\[4\] _0246_ _0247_ net65 vssd1 vssd1 vccd1 vccd1 MEM.next_mem3\[4\]
+ sky130_fd_sc_hd__a22o_1
X_0582_ net116 _0156_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__xnor2_1
X_0651_ _0210_ _0211_ _0213_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1134_ clknet_4_8_0_clk MEM.next_mem1\[7\] net40 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1065_ clknet_4_11_0_clk _0043_ net40 vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0918_ _0236_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__nor2_1
X_0849_ _0330_ _0326_ _0066_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_11_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6 MEM.mem1\[3\] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlygate4sd3_1
X_0703_ net100 _0240_ _0244_ CTR.time_out\[2\] vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0565_ CLKDIV.count\[5\] CLKDIV.count\[4\] _0140_ CLKDIV.count\[6\] vssd1 vssd1 vccd1
+ vccd1 _0146_ sky130_fd_sc_hd__a31o_1
X_0634_ MEM.mem5\[1\] _0075_ _0076_ MEM.mem2\[1\] _0070_ vssd1 vssd1 vccd1 vccd1 _0197_
+ sky130_fd_sc_hd__a221o_1
X_0496_ MEM.mem4\[9\] _0078_ net33 MEM.mem3\[9\] vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1117_ clknet_4_7_0_clk net101 net38 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1048_ clknet_4_10_0_clk _0026_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0548_ _0133_ _0126_ net26 _0128_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__a31o_1
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0479_ MEM.raddr\[0\] vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__clkbuf_8
X_0617_ MEM.mem4\[4\] _0078_ _0079_ MEM.mem3\[4\] _0179_ vssd1 vssd1 vccd1 vccd1 _0180_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0882_ _0084_ _0353_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or2_2
X_0951_ TIM.cnt\[2\] _0409_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1081_ clknet_4_6_0_clk MEM.next_mem5\[2\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0934_ _0236_ _0401_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__nor2_1
X_0865_ _0344_ vssd1 vssd1 vccd1 vccd1 FSM.next_state\[2\] sky130_fd_sc_hd__clkbuf_1
X_0796_ _0275_ _0288_ _0285_ vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__a21o_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0581_ _0157_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__clkbuf_1
X_0650_ _0191_ _0212_ _0183_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_1133_ clknet_4_8_0_clk MEM.next_mem1\[6\] net40 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1064_ clknet_4_11_0_clk _0042_ net41 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0917_ _0335_ _0387_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__nor2_2
X_0779_ _0259_ _0273_ _0260_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0848_ e1.edge_d e1.sync vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7 MEM.mem1\[4\] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dlygate4sd3_1
X_0702_ net93 _0240_ _0244_ _0200_ vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[1\] sky130_fd_sc_hd__a22o_1
X_0633_ _0069_ _0193_ _0194_ _0195_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_4_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0564_ CLKDIV.count\[5\] CLKDIV.count\[4\] CLKDIV.count\[6\] _0140_ vssd1 vssd1 vccd1
+ vccd1 _0145_ sky130_fd_sc_hd__and4_1
X_0495_ MEM.mem5\[9\] _0075_ _0076_ MEM.mem2\[9\] _0070_ vssd1 vssd1 vccd1 vccd1 _0089_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1116_ clknet_4_7_0_clk MEM.next_mem2\[1\] net41 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1047_ clknet_4_10_0_clk _0025_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0616_ MEM.mem5\[4\] _0075_ _0076_ MEM.mem2\[4\] _0070_ vssd1 vssd1 vccd1 vccd1 _0179_
+ sky130_fd_sc_hd__a221o_1
X_0547_ net31 _0130_ net29 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__a21o_1
X_0478_ MEM.raddr\[1\] vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0881_ _0084_ _0238_ _0349_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__a31o_1
X_0950_ TIM.cnt\[2\] _0409_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ clknet_4_7_0_clk MEM.next_mem5\[1\] net41 vssd1 vssd1 vccd1 vccd1 MEM.mem5\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0795_ _0286_ _0273_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__or2b_1
X_0933_ CTR.time_out\[9\] _0398_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__and2_1
X_0864_ _0340_ _0322_ _0337_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0580_ _0065_ _0155_ _0156_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1132_ clknet_4_12_0_clk MEM.next_mem1\[5\] net39 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1063_ clknet_4_11_0_clk _0041_ net41 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0916_ _0200_ _0229_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0778_ _0261_ _0273_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__nand2_1
X_0847_ _0066_ _0328_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold8 MEM.mem1\[8\] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dlygate4sd3_1
X_0563_ net122 _0142_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0701_ net99 _0240_ _0244_ _0229_ vssd1 vssd1 vccd1 vccd1 MEM.next_mem2\[0\] sky130_fd_sc_hd__a22o_1
X_0632_ TIM.cnt\[2\] _0085_ net34 CTR.time_out\[2\] vssd1 vssd1 vccd1 vccd1 _0195_
+ sky130_fd_sc_hd__a22o_1
X_0494_ _0069_ _0081_ _0087_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__a21oi_4
X_1046_ clknet_4_15_0_clk _0015_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1115_ clknet_4_6_0_clk MEM.next_mem2\[0\] net38 vssd1 vssd1 vccd1 vccd1 MEM.mem2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0615_ _0178_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0546_ _0135_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0477_ _0070_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1029_ clknet_4_5_0_clk _0020_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ _0111_ _0121_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__or2_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0880_ CLKDIV.secpulse _0354_ _0357_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ _0400_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__clkbuf_1
X_0863_ net34 _0341_ _0342_ _0324_ _0328_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0794_ _0259_ _0287_ vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__nand2_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1062_ clknet_4_11_0_clk _0040_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
X_1131_ clknet_4_12_0_clk MEM.next_mem1\[4\] net39 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0915_ _0189_ CTR.time_out\[2\] CTR.time_out\[5\] CTR.time_out\[4\] vssd1 vssd1 vccd1
+ vccd1 _0387_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0777_ _0263_ _0271_ _0272_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__a21oi_4
X_0846_ e1.edge_d e1.sync vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold9 MEM.mem1\[2\] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0700_ _0243_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__buf_4
X_0562_ _0144_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__clkbuf_1
X_0631_ _0071_ MEM.mem1\[2\] vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__or2_1
X_0493_ TIM.cnt\[11\] _0085_ _0086_ CTR.time_out\[11\] vssd1 vssd1 vccd1 vccd1 _0087_
+ sky130_fd_sc_hd__a22o_1
X_1114_ clknet_4_3_0_clk MEM.next_mem3\[11\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1045_ clknet_4_15_0_clk _0014_ net41 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0829_ _0313_ _0316_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0614_ _0065_ _0176_ _0177_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0545_ _0133_ _0128_ _0134_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0476_ MEM.raddr\[2\] vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__buf_6
X_1028_ clknet_4_5_0_clk _0019_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0528_ TIM.cnt\[7\] _0085_ _0118_ _0119_ _0120_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__a221o_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0931_ _0238_ _0397_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__and3_1
X_0862_ _0328_ _0323_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__nand2_1
X_0793_ _0260_ _0273_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1130_ clknet_4_9_0_clk MEM.next_mem1\[3\] net39 vssd1 vssd1 vccd1 vccd1 MEM.mem1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1061_ clknet_4_11_0_clk _0039_ net40 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0914_ _0385_ _0386_ net133 _0362_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__a2bb2o_1
X_0845_ _0066_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__nor2_4
X_0776_ _0223_ _0267_ _0217_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0561_ _0142_ _0143_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__and2_1
X_0630_ MEM.mem4\[2\] _0078_ net33 MEM.mem3\[2\] _0192_ vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__a221o_1
X_0492_ FSM.state\[2\] FSM.state\[3\] FSM.state\[1\] vssd1 vssd1 vccd1 vccd1 _0086_
+ sky130_fd_sc_hd__nor3b_4
X_1044_ clknet_4_15_0_clk _0013_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_1113_ clknet_4_0_0_clk MEM.next_mem3\[10\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0828_ _0298_ _0312_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__nand2_1
X_0759_ MEM.mem5\[0\] _0075_ _0076_ MEM.mem2\[0\] _0070_ vssd1 vssd1 vccd1 vccd1 _0255_
+ sky130_fd_sc_hd__a221o_1
X_0613_ CLKDIV.count\[21\] CLKDIV.count\[22\] _0173_ CLKDIV.count\[23\] vssd1 vssd1
+ vccd1 vccd1 _0177_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0544_ _0131_ _0130_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0475_ _0067_ _0068_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__nand2_8
X_1027_ clknet_4_5_0_clk _0018_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 CLKDIV.count\[20\] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ CTR.time_out\[7\] _0086_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0792_ _0273_ _0286_ vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__nand2_1
X_0930_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
X_0861_ _0066_ _0328_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1060_ clknet_4_11_0_clk _0038_ net41 vssd1 vssd1 vccd1 vccd1 TIM.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0775_ _0209_ _0269_ _0270_ _0218_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a211o_1
X_0913_ _0381_ _0382_ _0384_ _0362_ _0236_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__a311o_1
X_0844_ FSM.state\[2\] FSM.state\[1\] FSM.state\[3\] vssd1 vssd1 vccd1 vccd1 _0326_
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0560_ CLKDIV.count\[4\] _0140_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__or2_1
X_0491_ _0082_ _0084_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__nand2_8
XFILLER_0_29_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1043_ clknet_4_15_0_clk _0012_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1112_ clknet_4_3_0_clk MEM.next_mem3\[9\] net36 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ _0299_ _0314_ _0315_ vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__o21a_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0758_ CTR.time_out\[11\] _0253_ _0254_ net71 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[11\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0689_ CTR.time_out\[7\] _0233_ _0237_ net52 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0612_ CLKDIV.count\[22\] CLKDIV.count\[23\] _0174_ vssd1 vssd1 vccd1 vccd1 _0176_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0543_ net31 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__inv_2
X_0474_ FSM.state\[3\] FSM.state\[1\] _0066_ FSM.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _0068_ sky130_fd_sc_hd__or4bb_4
X_1026_ clknet_4_5_0_clk _0017_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold80 CLKDIV.count\[3\] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 TIM.cnt\[2\] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0526_ _0067_ _0068_ _0071_ MEM.mem1\[7\] vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1009_ _0189_ CTR.time_out\[4\] _0452_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__nand3_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0509_ TIM.cnt\[10\] _0085_ _0098_ _0099_ _0100_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__a221o_2
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0791_ _0258_ _0260_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__xnor2_1
X_0860_ _0066_ _0231_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__and2_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0989_ MEM.addr\[0\] _0232_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0912_ _0381_ _0382_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__a21oi_1
X_0774_ _0209_ _0267_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0843_ _0066_ net34 _0324_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0490_ _0083_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1042_ clknet_4_15_0_clk _0010_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_1111_ clknet_4_0_0_clk MEM.next_mem3\[8\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0826_ _0297_ _0298_ _0308_ _0312_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__or4b_1
XFILLER_0_10_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0757_ CTR.time_out\[10\] _0253_ _0254_ net88 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[10\]
+ sky130_fd_sc_hd__a22o_1
X_0688_ CTR.time_out\[6\] _0233_ _0237_ net55 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[6\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0611_ net123 _0174_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__xor2_1
X_0542_ net31 _0130_ net29 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__a21o_1
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0473_ FSM.state\[3\] _0066_ FSM.state\[1\] FSM.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _0067_ sky130_fd_sc_hd__or4bb_4
X_1025_ clknet_4_5_0_clk _0016_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_0809_ _0121_ _0134_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold81 CLKDIV.count\[5\] vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 CLKDIV.count\[13\] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 TIM.cnt\[11\] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0525_ _0114_ _0115_ _0116_ _0117_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__or4_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _0389_ _0455_ _0456_ _0454_ _0189_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__a32o_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0508_ _0092_ _0093_ _0101_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__a21o_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0790_ _0274_ _0275_ _0285_ vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__a21o_1
XFILLER_0_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0988_ _0242_ _0236_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0911_ TIM.cnt\[11\] _0084_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__xor2_1
X_0842_ _0238_ _0323_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__nor2_1
X_0773_ _0212_ net17 _0266_ _0268_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1110_ clknet_4_0_0_clk MEM.next_mem3\[7\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem3\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1041_ clknet_4_14_0_clk _0009_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0825_ _0308_ _0313_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0756_ CTR.time_out\[9\] _0253_ _0254_ net61 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[9\]
+ sky130_fd_sc_hd__a22o_1
X_0687_ CTR.time_out\[5\] _0233_ _0237_ net46 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0610_ _0174_ _0175_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__nor2_1
X_0541_ _0132_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0472_ FSM.state\[0\] vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__buf_4
X_1024_ clknet_4_5_0_clk _0011_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[1\] sky130_fd_sc_hd__dfrtp_1
X_0808_ _0129_ _0290_ _0296_ _0131_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0739_ CTR.time_out\[8\] _0249_ _0250_ net67 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[8\]
+ sky130_fd_sc_hd__a22o_1
Xhold82 CLKDIV.count\[22\] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 MEM.next_mem2\[2\] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 TIM.cnt\[7\] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 MEM.mem5\[6\] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ _0072_ _0073_ MEM.mem5\[7\] _0070_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__a31o_1
X_1007_ _0189_ _0452_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__nand2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput4 net4 vssd1 vssd1 vccd1 vccd1 out_0[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0507_ TIM.cnt\[10\] _0085_ _0098_ _0099_ _0100_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__a221oi_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0987_ _0442_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0772_ _0264_ _0265_ _0267_ _0220_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__o31a_1
X_0910_ _0364_ _0382_ _0383_ _0362_ net128 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__a32o_1
X_0841_ _0066_ _0321_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1040_ clknet_4_14_0_clk _0008_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0824_ _0298_ _0312_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0755_ CTR.time_out\[8\] _0253_ _0254_ net110 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[8\]
+ sky130_fd_sc_hd__a22o_1
X_0686_ CTR.time_out\[4\] _0233_ _0237_ net48 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[4\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0471_ _0065_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
X_0540_ _0126_ _0131_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1023_ clknet_4_7_0_clk _0000_ net37 vssd1 vssd1 vccd1 vccd1 CLKDIV.count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0807_ _0128_ _0294_ _0295_ net26 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__o211ai_1
X_0738_ CTR.time_out\[7\] _0249_ _0250_ net79 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[7\]
+ sky130_fd_sc_hd__a22o_1
X_0669_ _0215_ _0224_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold83 CLKDIV.count\[21\] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 CLKDIV.count\[19\] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 CLKDIV.count\[9\] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 MEM.addr\[0\] vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold50 MEM.mem2\[6\] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0523_ _0073_ _0070_ MEM.mem4\[7\] _0072_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__and4bb_1
X_1006_ _0189_ _0452_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput5 net5 vssd1 vssd1 vccd1 vccd1 out_0[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0506_ CTR.time_out\[10\] _0086_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__and2_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0986_ _0441_ TIM.cnt\[0\] _0359_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0771_ _0203_ _0216_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__and2b_1
X_0840_ _0082_ _0321_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0969_ _0352_ _0349_ _0327_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0823_ TIM.cnt\[6\] _0085_ _0086_ CTR.time_out\[6\] _0311_ vssd1 vssd1 vccd1 vccd1
+ _0312_ sky130_fd_sc_hd__a221o_1
X_0754_ CTR.time_out\[7\] _0253_ _0254_ net82 vssd1 vssd1 vccd1 vccd1 MEM.next_mem5\[7\]
+ sky130_fd_sc_hd__a22o_1
X_0685_ _0189_ _0233_ _0237_ net47 vssd1 vssd1 vccd1 vccd1 MEM.next_mem1\[3\] sky130_fd_sc_hd__a22o_1
X_1099_ clknet_4_0_0_clk MEM.next_mem4\[8\] net35 vssd1 vssd1 vccd1 vccd1 MEM.mem4\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_0470_ _0059_ _0064_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__or2_2
X_1022_ clknet_4_15_0_clk _0024_ net39 vssd1 vssd1 vccd1 vccd1 CLKDIV.secpulse sky130_fd_sc_hd__dfrtp_4
X_0668_ _0227_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
X_0806_ _0111_ _0128_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0737_ CTR.time_out\[6\] _0249_ _0250_ net74 vssd1 vssd1 vccd1 vccd1 MEM.next_mem4\[6\]
+ sky130_fd_sc_hd__a22o_1
X_0599_ CLKDIV.count\[17\] CLKDIV.count\[16\] CLKDIV.count\[18\] _0163_ vssd1 vssd1
+ vccd1 vccd1 _0168_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold40 MEM.mem4\[10\] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold73 CLKDIV.count\[0\] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 CLKDIV.count\[2\] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 MEM.mem5\[1\] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 TIM.cnt\[8\] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 MEM.mem3\[1\] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0522_ _0072_ _0073_ MEM.mem2\[7\] vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__nor3b_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ _0389_ _0451_ _0453_ _0454_ CTR.time_out\[2\] vssd1 vssd1 vccd1 vccd1 _0053_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 out_3[5] sky130_fd_sc_hd__clkbuf_4
Xoutput6 net6 vssd1 vssd1 vccd1 vccd1 out_0[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0505_ _0067_ _0068_ _0071_ MEM.mem1\[10\] vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__o2bb2a_1
.ends

