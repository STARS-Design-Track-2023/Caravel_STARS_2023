// This is the unpowered netlist.
module Eighty_Twos (clk,
    cs,
    nrst,
    store_en,
    gpi,
    gpo);
 input clk;
 input cs;
 input nrst;
 output store_en;
 input [33:0] gpi;
 output [33:0] gpo;

 wire \ALU.flags_to_alu[0] ;
 wire \ALU.flags_to_alu[1] ;
 wire \ALU.flags_to_alu[2] ;
 wire \ALU.flags_to_alu[3] ;
 wire \ALU.flags_to_alu[4] ;
 wire \ALU.flags_to_alu[5] ;
 wire \ALU.flags_to_alu[6] ;
 wire \ALU.flags_to_alu[7] ;
 wire \ALU.immediate[0] ;
 wire \ALU.immediate[10] ;
 wire \ALU.immediate[11] ;
 wire \ALU.immediate[12] ;
 wire \ALU.immediate[13] ;
 wire \ALU.immediate[14] ;
 wire \ALU.immediate[15] ;
 wire \ALU.immediate[1] ;
 wire \ALU.immediate[2] ;
 wire \ALU.immediate[3] ;
 wire \ALU.immediate[4] ;
 wire \ALU.immediate[5] ;
 wire \ALU.immediate[6] ;
 wire \ALU.immediate[7] ;
 wire \ALU.immediate[8] ;
 wire \ALU.immediate[9] ;
 wire \ByteBuffer.counter[0] ;
 wire \ByteBuffer.counter[1] ;
 wire \ByteBuffer.instr[16] ;
 wire \ByteBuffer.instr[17] ;
 wire \ByteBuffer.instr[18] ;
 wire \ByteBuffer.instr[19] ;
 wire \ByteBuffer.instr[20] ;
 wire \ByteBuffer.instr[21] ;
 wire \ByteBuffer.instr[22] ;
 wire \ByteBuffer.instr[23] ;
 wire \ByteBuffer.next_counter[0] ;
 wire \ByteBuffer.next_counter[1] ;
 wire \ByteDecoder.num_bytes[1] ;
 wire \ByteDecoder.num_bytes[2] ;
 wire \ByteDecoder.num_bytes[3] ;
 wire \ByteDecoder.state[0] ;
 wire \ByteDecoder.state[1] ;
 wire \FSM.next_state[0] ;
 wire \FSM.next_state[1] ;
 wire \MemControl.state[0] ;
 wire \MemControl.state[1] ;
 wire \MemControl.state[2] ;
 wire \PC.i_mem_addr[0] ;
 wire \PC.i_mem_addr[10] ;
 wire \PC.i_mem_addr[11] ;
 wire \PC.i_mem_addr[12] ;
 wire \PC.i_mem_addr[13] ;
 wire \PC.i_mem_addr[14] ;
 wire \PC.i_mem_addr[15] ;
 wire \PC.i_mem_addr[1] ;
 wire \PC.i_mem_addr[2] ;
 wire \PC.i_mem_addr[3] ;
 wire \PC.i_mem_addr[4] ;
 wire \PC.i_mem_addr[5] ;
 wire \PC.i_mem_addr[6] ;
 wire \PC.i_mem_addr[7] ;
 wire \PC.i_mem_addr[8] ;
 wire \PC.i_mem_addr[9] ;
 wire \RegFile.A[0] ;
 wire \RegFile.A[1] ;
 wire \RegFile.A[2] ;
 wire \RegFile.A[3] ;
 wire \RegFile.A[4] ;
 wire \RegFile.A[5] ;
 wire \RegFile.A[6] ;
 wire \RegFile.A[7] ;
 wire \RegFile.B[0] ;
 wire \RegFile.B[1] ;
 wire \RegFile.B[2] ;
 wire \RegFile.B[3] ;
 wire \RegFile.B[4] ;
 wire \RegFile.B[5] ;
 wire \RegFile.B[6] ;
 wire \RegFile.B[7] ;
 wire \RegFile.C[0] ;
 wire \RegFile.C[1] ;
 wire \RegFile.C[2] ;
 wire \RegFile.C[3] ;
 wire \RegFile.C[4] ;
 wire \RegFile.C[5] ;
 wire \RegFile.C[6] ;
 wire \RegFile.C[7] ;
 wire \RegFile.D[0] ;
 wire \RegFile.D[1] ;
 wire \RegFile.D[2] ;
 wire \RegFile.D[3] ;
 wire \RegFile.D[4] ;
 wire \RegFile.D[5] ;
 wire \RegFile.D[6] ;
 wire \RegFile.D[7] ;
 wire \RegFile.E[0] ;
 wire \RegFile.E[1] ;
 wire \RegFile.E[2] ;
 wire \RegFile.E[3] ;
 wire \RegFile.E[4] ;
 wire \RegFile.E[5] ;
 wire \RegFile.E[6] ;
 wire \RegFile.E[7] ;
 wire \RegFile.H[0] ;
 wire \RegFile.H[1] ;
 wire \RegFile.H[2] ;
 wire \RegFile.H[3] ;
 wire \RegFile.H[4] ;
 wire \RegFile.H[5] ;
 wire \RegFile.H[6] ;
 wire \RegFile.H[7] ;
 wire \RegFile.L[0] ;
 wire \RegFile.L[1] ;
 wire \RegFile.L[2] ;
 wire \RegFile.L[3] ;
 wire \RegFile.L[4] ;
 wire \RegFile.L[5] ;
 wire \RegFile.L[6] ;
 wire \RegFile.L[7] ;
 wire _0000_;
 wire _0001_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire clknet_0__0514_;
 wire clknet_0__0515_;
 wire clknet_0__0516_;
 wire clknet_0__0517_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf__0514_;
 wire clknet_1_0__leaf__0515_;
 wire clknet_1_0__leaf__0516_;
 wire clknet_1_0__leaf__0517_;
 wire clknet_1_1__leaf__0514_;
 wire clknet_1_1__leaf__0515_;
 wire clknet_1_1__leaf__0516_;
 wire clknet_1_1__leaf__0517_;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0204_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_91 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__inv_2 _1275_ (.A(\ByteBuffer.instr[19] ),
    .Y(_0618_));
 sky130_fd_sc_hd__clkbuf_8 _1276_ (.A(\ByteBuffer.instr[16] ),
    .X(_0619_));
 sky130_fd_sc_hd__inv_2 _1277_ (.A(\ByteBuffer.instr[17] ),
    .Y(_0620_));
 sky130_fd_sc_hd__or2_2 _1278_ (.A(_0619_),
    .B(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__buf_6 _1279_ (.A(\ByteBuffer.instr[17] ),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_2 _1280_ (.A(_0619_),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__clkbuf_8 _1281_ (.A(\ByteBuffer.instr[18] ),
    .X(_0624_));
 sky130_fd_sc_hd__or2_1 _1282_ (.A(\ByteBuffer.instr[23] ),
    .B(\ByteBuffer.instr[22] ),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_4 _1283_ (.A(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__nand2_1 _1284_ (.A(\ByteDecoder.state[1] ),
    .B(\ByteDecoder.state[0] ),
    .Y(_0627_));
 sky130_fd_sc_hd__or3_4 _1285_ (.A(_0624_),
    .B(_0626_),
    .C(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__nor2_8 _1286_ (.A(_0623_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__buf_8 _1287_ (.A(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__o21a_2 _1288_ (.A1(_0618_),
    .A2(_0621_),
    .B1(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__nand2b_4 _1289_ (.A_N(\ByteBuffer.instr[23] ),
    .B(\ByteBuffer.instr[22] ),
    .Y(_0632_));
 sky130_fd_sc_hd__a21boi_1 _1290_ (.A1(_0619_),
    .A2(_0622_),
    .B1_N(_0624_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(\ByteBuffer.instr[20] ),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__xor2_4 _1292_ (.A(\ByteBuffer.instr[17] ),
    .B(_0624_),
    .X(_0635_));
 sky130_fd_sc_hd__nand3b_2 _1293_ (.A_N(_0624_),
    .B(_0622_),
    .C(\ByteBuffer.instr[21] ),
    .Y(_0636_));
 sky130_fd_sc_hd__and3b_1 _1294_ (.A_N(_0626_),
    .B(_0635_),
    .C(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__a2bb2o_4 _1295_ (.A1_N(_0622_),
    .A2_N(_0632_),
    .B1(_0634_),
    .B2(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__and2b_1 _1296_ (.A_N(_0624_),
    .B(\ByteBuffer.instr[17] ),
    .X(_0639_));
 sky130_fd_sc_hd__a21bo_1 _1297_ (.A1(\ByteBuffer.instr[20] ),
    .A2(_0639_),
    .B1_N(_0632_),
    .X(_0640_));
 sky130_fd_sc_hd__a21bo_1 _1298_ (.A1(_0619_),
    .A2(_0622_),
    .B1_N(_0624_),
    .X(_0641_));
 sky130_fd_sc_hd__and4bb_4 _1299_ (.A_N(\ByteBuffer.instr[17] ),
    .B_N(_0624_),
    .C(\ByteBuffer.instr[19] ),
    .D(_0619_),
    .X(_0642_));
 sky130_fd_sc_hd__or4bb_1 _1300_ (.A(\ByteBuffer.instr[21] ),
    .B(_0624_),
    .C_N(\ByteBuffer.instr[17] ),
    .D_N(\ByteBuffer.instr[20] ),
    .X(_0643_));
 sky130_fd_sc_hd__o221ai_4 _1301_ (.A1(_0618_),
    .A2(_0641_),
    .B1(_0635_),
    .B2(_0642_),
    .C1(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__buf_8 _1302_ (.A(\ByteBuffer.instr[23] ),
    .X(_0645_));
 sky130_fd_sc_hd__a221oi_2 _1303_ (.A1(_0619_),
    .A2(_0640_),
    .B1(_0644_),
    .B2(_0632_),
    .C1(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__inv_2 _1304_ (.A(_0624_),
    .Y(_0647_));
 sky130_fd_sc_hd__and2_2 _1305_ (.A(\ByteBuffer.instr[23] ),
    .B(\ByteBuffer.instr[22] ),
    .X(_0648_));
 sky130_fd_sc_hd__and3_1 _1306_ (.A(_0620_),
    .B(_0647_),
    .C(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__clkbuf_4 _1307_ (.A(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__or3_1 _1308_ (.A(_0638_),
    .B(net54),
    .C(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__buf_4 _1309_ (.A(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or2_1 _1310_ (.A(_0623_),
    .B(_0628_),
    .X(_0653_));
 sky130_fd_sc_hd__clkbuf_8 _1311_ (.A(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__buf_8 _1312_ (.A(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _1313_ (.A(_0619_),
    .B(_0622_),
    .Y(_0656_));
 sky130_fd_sc_hd__nor2_1 _1314_ (.A(\ByteBuffer.instr[21] ),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__and2_1 _1315_ (.A(\ByteDecoder.state[1] ),
    .B(\ByteDecoder.state[0] ),
    .X(_0658_));
 sky130_fd_sc_hd__buf_4 _1316_ (.A(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__and2_1 _1317_ (.A(\ByteBuffer.instr[20] ),
    .B(\ByteBuffer.instr[21] ),
    .X(_0660_));
 sky130_fd_sc_hd__and3b_1 _1318_ (.A_N(_0619_),
    .B(_0622_),
    .C(_0624_),
    .X(_0661_));
 sky130_fd_sc_hd__and4_1 _1319_ (.A(\ByteBuffer.instr[22] ),
    .B(_0618_),
    .C(_0660_),
    .D(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__nor2_1 _1320_ (.A(_0645_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__o311a_4 _1321_ (.A1(_0626_),
    .A2(_0657_),
    .A3(_0635_),
    .B1(_0659_),
    .C1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__o211a_1 _1322_ (.A1(_0622_),
    .A2(_0618_),
    .B1(_0647_),
    .C1(_0619_),
    .X(_0665_));
 sky130_fd_sc_hd__or2_2 _1323_ (.A(_0633_),
    .B(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__or4bb_1 _1324_ (.A(_0622_),
    .B(_0624_),
    .C_N(\ByteBuffer.instr[19] ),
    .D_N(_0619_),
    .X(_0667_));
 sky130_fd_sc_hd__nand2b_1 _1325_ (.A_N(\ByteBuffer.instr[20] ),
    .B(\ByteBuffer.instr[21] ),
    .Y(_0668_));
 sky130_fd_sc_hd__nor2_1 _1326_ (.A(_0667_),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__inv_2 _1327_ (.A(_0645_),
    .Y(_0670_));
 sky130_fd_sc_hd__or3_1 _1328_ (.A(_0670_),
    .B(_0661_),
    .C(_0639_),
    .X(_0671_));
 sky130_fd_sc_hd__xnor2_4 _1329_ (.A(_0645_),
    .B(\ByteBuffer.instr[22] ),
    .Y(_0672_));
 sky130_fd_sc_hd__o211a_1 _1330_ (.A1(_0669_),
    .A2(_0671_),
    .B1(_0672_),
    .C1(_0659_),
    .X(_0673_));
 sky130_fd_sc_hd__o21ai_4 _1331_ (.A1(_0666_),
    .A2(_0626_),
    .B1(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__nor2_8 _1332_ (.A(_0664_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__nor2_4 _1333_ (.A(_0655_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__a221o_2 _1334_ (.A1(_0619_),
    .A2(_0640_),
    .B1(_0644_),
    .B2(_0632_),
    .C1(_0645_),
    .X(_0677_));
 sky130_fd_sc_hd__nand2_8 _1335_ (.A(_0645_),
    .B(\ByteBuffer.instr[22] ),
    .Y(_0678_));
 sky130_fd_sc_hd__or3_4 _1336_ (.A(_0622_),
    .B(_0624_),
    .C(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__a21oi_4 _1337_ (.A1(_0677_),
    .A2(_0679_),
    .B1(_0638_),
    .Y(_0680_));
 sky130_fd_sc_hd__a22o_4 _1338_ (.A1(_0619_),
    .A2(_0640_),
    .B1(_0644_),
    .B2(_0632_),
    .X(_0681_));
 sky130_fd_sc_hd__and2_1 _1339_ (.A(_0638_),
    .B(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_8 _1340_ (.A(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__o2bb2a_2 _1341_ (.A1_N(_0637_),
    .A2_N(_0634_),
    .B1(_0632_),
    .B2(_0622_),
    .X(_0684_));
 sky130_fd_sc_hd__a21oi_4 _1342_ (.A1(_0677_),
    .A2(_0679_),
    .B1(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__and3_1 _1343_ (.A(_0684_),
    .B(_0677_),
    .C(_0679_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_8 _1344_ (.A(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__a221o_1 _1345_ (.A1(\RegFile.D[6] ),
    .A2(_0683_),
    .B1(net51),
    .B2(\RegFile.B[6] ),
    .C1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__a21o_1 _1346_ (.A1(\RegFile.H[6] ),
    .A2(net52),
    .B1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__o211a_1 _1347_ (.A1(\RegFile.A[6] ),
    .A2(_0652_),
    .B1(_0676_),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__inv_2 _1348_ (.A(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__o21a_2 _1349_ (.A1(_0666_),
    .A2(_0626_),
    .B1(_0673_),
    .X(_0692_));
 sky130_fd_sc_hd__nor2_8 _1350_ (.A(_0664_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__or2_2 _1351_ (.A(_0670_),
    .B(_0619_),
    .X(_0694_));
 sky130_fd_sc_hd__inv_2 _1352_ (.A(\ByteBuffer.instr[21] ),
    .Y(_0695_));
 sky130_fd_sc_hd__or3b_2 _1353_ (.A(_0619_),
    .B(_0624_),
    .C_N(_0622_),
    .X(_0696_));
 sky130_fd_sc_hd__inv_2 _1354_ (.A(\ByteBuffer.instr[20] ),
    .Y(_0697_));
 sky130_fd_sc_hd__o2111ai_4 _1355_ (.A1(_0695_),
    .A2(_0696_),
    .B1(_0672_),
    .C1(_0642_),
    .D1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a21o_4 _1356_ (.A1(_0694_),
    .A2(_0698_),
    .B1(_0648_),
    .X(_0699_));
 sky130_fd_sc_hd__inv_2 _1357_ (.A(\ByteBuffer.instr[22] ),
    .Y(_0700_));
 sky130_fd_sc_hd__nand2_1 _1358_ (.A(_0645_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__o22a_2 _1359_ (.A1(\ByteBuffer.instr[21] ),
    .A2(_0667_),
    .B1(_0668_),
    .B2(_0696_),
    .X(_0702_));
 sky130_fd_sc_hd__o22a_4 _1360_ (.A1(_0622_),
    .A2(_0701_),
    .B1(_0702_),
    .B2(_0626_),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_8 _1361_ (.A(_0699_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__nor2_8 _1362_ (.A(_0699_),
    .B(_0703_),
    .Y(_0705_));
 sky130_fd_sc_hd__o22ai_4 _1363_ (.A1(_0622_),
    .A2(_0701_),
    .B1(_0702_),
    .B2(_0626_),
    .Y(_0706_));
 sky130_fd_sc_hd__nor2_8 _1364_ (.A(_0699_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21oi_4 _1365_ (.A1(_0694_),
    .A2(_0698_),
    .B1(_0648_),
    .Y(_0708_));
 sky130_fd_sc_hd__nor2_4 _1366_ (.A(_0708_),
    .B(_0703_),
    .Y(_0709_));
 sky130_fd_sc_hd__a22o_1 _1367_ (.A1(\RegFile.H[6] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[6] ),
    .X(_0710_));
 sky130_fd_sc_hd__nor2_8 _1368_ (.A(_0708_),
    .B(net53),
    .Y(_0711_));
 sky130_fd_sc_hd__a211o_1 _1369_ (.A1(\RegFile.B[6] ),
    .A2(_0705_),
    .B1(_0710_),
    .C1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__o211a_1 _1370_ (.A1(\RegFile.A[6] ),
    .A2(_0704_),
    .B1(_0712_),
    .C1(_0630_),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _1371_ (.A1(\ALU.immediate[14] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__nor2_1 _1372_ (.A(_0691_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__and2_1 _1373_ (.A(_0690_),
    .B(_0714_),
    .X(_0716_));
 sky130_fd_sc_hd__nor2_1 _1374_ (.A(_0690_),
    .B(_0714_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor2_1 _1375_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a221o_1 _1376_ (.A1(\RegFile.D[3] ),
    .A2(_0683_),
    .B1(net51),
    .B2(\RegFile.B[3] ),
    .C1(_0687_),
    .X(_0719_));
 sky130_fd_sc_hd__a21o_1 _1377_ (.A1(\RegFile.H[3] ),
    .A2(net52),
    .B1(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__o211a_2 _1378_ (.A1(\RegFile.A[3] ),
    .A2(_0652_),
    .B1(_0676_),
    .C1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__a22o_1 _1379_ (.A1(\RegFile.H[3] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[3] ),
    .X(_0722_));
 sky130_fd_sc_hd__a211o_1 _1380_ (.A1(\RegFile.B[3] ),
    .A2(_0705_),
    .B1(_0722_),
    .C1(_0711_),
    .X(_0723_));
 sky130_fd_sc_hd__o211a_1 _1381_ (.A1(\RegFile.A[3] ),
    .A2(_0704_),
    .B1(_0723_),
    .C1(_0630_),
    .X(_0724_));
 sky130_fd_sc_hd__a22o_2 _1382_ (.A1(\ALU.immediate[11] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__xnor2_2 _1383_ (.A(_0721_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__a221o_1 _1384_ (.A1(\RegFile.D[2] ),
    .A2(_0683_),
    .B1(net51),
    .B2(\RegFile.B[2] ),
    .C1(_0687_),
    .X(_0727_));
 sky130_fd_sc_hd__a21o_1 _1385_ (.A1(\RegFile.H[2] ),
    .A2(net52),
    .B1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__o211a_1 _1386_ (.A1(\RegFile.A[2] ),
    .A2(_0652_),
    .B1(_0676_),
    .C1(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _1387_ (.A1(\RegFile.H[2] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[2] ),
    .X(_0730_));
 sky130_fd_sc_hd__a211o_1 _1388_ (.A1(\RegFile.B[2] ),
    .A2(_0705_),
    .B1(_0730_),
    .C1(_0711_),
    .X(_0731_));
 sky130_fd_sc_hd__o211a_1 _1389_ (.A1(\RegFile.A[2] ),
    .A2(_0704_),
    .B1(_0731_),
    .C1(_0630_),
    .X(_0732_));
 sky130_fd_sc_hd__a22o_1 _1390_ (.A1(\ALU.immediate[10] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(_0729_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__or2_1 _1392_ (.A(_0729_),
    .B(_0733_),
    .X(_0735_));
 sky130_fd_sc_hd__and2_2 _1393_ (.A(_0734_),
    .B(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__inv_2 _1394_ (.A(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__a221o_1 _1395_ (.A1(\RegFile.D[1] ),
    .A2(_0683_),
    .B1(net51),
    .B2(\RegFile.B[1] ),
    .C1(_0687_),
    .X(_0738_));
 sky130_fd_sc_hd__a21o_1 _1396_ (.A1(\RegFile.H[1] ),
    .A2(net52),
    .B1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__o211ai_4 _1397_ (.A1(\RegFile.A[1] ),
    .A2(_0652_),
    .B1(_0676_),
    .C1(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__nor2_1 _1398_ (.A(\RegFile.A[1] ),
    .B(_0704_),
    .Y(_0741_));
 sky130_fd_sc_hd__a22o_1 _1399_ (.A1(\RegFile.H[1] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[1] ),
    .X(_0742_));
 sky130_fd_sc_hd__a211o_1 _1400_ (.A1(\RegFile.B[1] ),
    .A2(_0705_),
    .B1(_0742_),
    .C1(_0711_),
    .X(_0743_));
 sky130_fd_sc_hd__and3b_1 _1401_ (.A_N(_0741_),
    .B(_0743_),
    .C(_0630_),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _1402_ (.A1(\ALU.immediate[9] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(_0740_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__a221o_1 _1404_ (.A1(\RegFile.H[0] ),
    .A2(net52),
    .B1(_0683_),
    .B2(\RegFile.D[0] ),
    .C1(_0687_),
    .X(_0747_));
 sky130_fd_sc_hd__a21o_1 _1405_ (.A1(\RegFile.B[0] ),
    .A2(net51),
    .B1(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__o211a_1 _1406_ (.A1(\RegFile.A[0] ),
    .A2(_0652_),
    .B1(_0676_),
    .C1(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _1407_ (.A1(\RegFile.H[0] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[0] ),
    .X(_0750_));
 sky130_fd_sc_hd__a211o_1 _1408_ (.A1(\RegFile.B[0] ),
    .A2(_0705_),
    .B1(_0750_),
    .C1(_0711_),
    .X(_0751_));
 sky130_fd_sc_hd__o211a_1 _1409_ (.A1(\RegFile.A[0] ),
    .A2(_0704_),
    .B1(_0751_),
    .C1(_0630_),
    .X(_0752_));
 sky130_fd_sc_hd__a22o_1 _1410_ (.A1(\ALU.immediate[8] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__nand2_1 _1411_ (.A(_0749_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__or2_1 _1412_ (.A(_0749_),
    .B(_0753_),
    .X(_0755_));
 sky130_fd_sc_hd__nand2_2 _1413_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__or3_2 _1414_ (.A(\ByteBuffer.instr[22] ),
    .B(_0642_),
    .C(_0635_),
    .X(_0757_));
 sky130_fd_sc_hd__a21bo_1 _1415_ (.A1(_0619_),
    .A2(_0622_),
    .B1_N(\ByteBuffer.instr[21] ),
    .X(_0758_));
 sky130_fd_sc_hd__a21o_1 _1416_ (.A1(_0700_),
    .A2(_0758_),
    .B1(_0647_),
    .X(_0759_));
 sky130_fd_sc_hd__and3_4 _1417_ (.A(_0670_),
    .B(_0757_),
    .C(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__and4_4 _1418_ (.A(_0684_),
    .B(_0677_),
    .C(_0679_),
    .D(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__a31oi_4 _1419_ (.A1(_0670_),
    .A2(_0757_),
    .A3(_0759_),
    .B1(_0650_),
    .Y(_0762_));
 sky130_fd_sc_hd__o211a_2 _1420_ (.A1(net54),
    .A2(_0650_),
    .B1(_0762_),
    .C1(_0638_),
    .X(_0763_));
 sky130_fd_sc_hd__a22o_1 _1421_ (.A1(\RegFile.E[5] ),
    .A2(_0761_),
    .B1(_0763_),
    .B2(\RegFile.H[5] ),
    .X(_0764_));
 sky130_fd_sc_hd__o211a_2 _1422_ (.A1(net54),
    .A2(_0650_),
    .B1(_0762_),
    .C1(_0684_),
    .X(_0765_));
 sky130_fd_sc_hd__a31o_1 _1423_ (.A1(_0670_),
    .A2(_0757_),
    .A3(_0759_),
    .B1(_0650_),
    .X(_0766_));
 sky130_fd_sc_hd__o211a_2 _1424_ (.A1(net54),
    .A2(_0650_),
    .B1(_0766_),
    .C1(_0684_),
    .X(_0767_));
 sky130_fd_sc_hd__and4_1 _1425_ (.A(\RegFile.C[5] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0768_));
 sky130_fd_sc_hd__a221o_1 _1426_ (.A1(\ALU.flags_to_alu[5] ),
    .A2(_0765_),
    .B1(_0767_),
    .B2(\RegFile.D[5] ),
    .C1(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__and3_2 _1427_ (.A(_0638_),
    .B(_0681_),
    .C(_0762_),
    .X(_0770_));
 sky130_fd_sc_hd__o211a_4 _1428_ (.A1(net54),
    .A2(_0650_),
    .B1(_0766_),
    .C1(_0638_),
    .X(_0771_));
 sky130_fd_sc_hd__nor4_1 _1429_ (.A(_0638_),
    .B(net54),
    .C(_0650_),
    .D(_0760_),
    .Y(_0772_));
 sky130_fd_sc_hd__a221o_1 _1430_ (.A1(\RegFile.L[5] ),
    .A2(_0770_),
    .B1(_0771_),
    .B2(\RegFile.B[5] ),
    .C1(net50),
    .X(_0773_));
 sky130_fd_sc_hd__or2_2 _1431_ (.A(_0760_),
    .B(_0652_),
    .X(_0774_));
 sky130_fd_sc_hd__o32a_2 _1432_ (.A1(_0764_),
    .A2(_0769_),
    .A3(_0773_),
    .B1(_0774_),
    .B2(\RegFile.A[5] ),
    .X(_0775_));
 sky130_fd_sc_hd__a221o_1 _1433_ (.A1(\RegFile.E[5] ),
    .A2(_0683_),
    .B1(_0685_),
    .B2(\RegFile.C[5] ),
    .C1(_0654_),
    .X(_0776_));
 sky130_fd_sc_hd__a22o_1 _1434_ (.A1(\RegFile.L[5] ),
    .A2(_0680_),
    .B1(_0687_),
    .B2(\ALU.flags_to_alu[5] ),
    .X(_0777_));
 sky130_fd_sc_hd__or2_2 _1435_ (.A(_0776_),
    .B(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__or2_1 _1436_ (.A(_0664_),
    .B(_0674_),
    .X(_0779_));
 sky130_fd_sc_hd__clkbuf_8 _1437_ (.A(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o211ai_4 _1438_ (.A1(_0629_),
    .A2(_0775_),
    .B1(_0778_),
    .C1(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_1 _1439_ (.A(\ALU.immediate[5] ),
    .B(_0675_),
    .Y(_0782_));
 sky130_fd_sc_hd__o2bb2a_1 _1440_ (.A1_N(_0672_),
    .A2_N(_0642_),
    .B1(_0624_),
    .B2(_0670_),
    .X(_0783_));
 sky130_fd_sc_hd__and3_4 _1441_ (.A(_0783_),
    .B(_0708_),
    .C(net53),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_2 _1442_ (.A1(_0645_),
    .A2(_0647_),
    .B1(_0642_),
    .B2(_0672_),
    .X(_0785_));
 sky130_fd_sc_hd__and3_2 _1443_ (.A(_0785_),
    .B(_0708_),
    .C(_0703_),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _1444_ (.A1(\RegFile.H[5] ),
    .A2(_0784_),
    .B1(_0786_),
    .B2(\RegFile.D[5] ),
    .X(_0787_));
 sky130_fd_sc_hd__and3_2 _1445_ (.A(_0783_),
    .B(_0708_),
    .C(_0703_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_4 _1446_ (.A(_0678_),
    .B(_0785_),
    .Y(_0789_));
 sky130_fd_sc_hd__or2_1 _1447_ (.A(\RegFile.E[5] ),
    .B(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__a22o_1 _1448_ (.A1(\ALU.flags_to_alu[5] ),
    .A2(_0788_),
    .B1(_0790_),
    .B2(_0711_),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_2 _1449_ (.A(_0648_),
    .B(_0783_),
    .Y(_0792_));
 sky130_fd_sc_hd__and3_2 _1450_ (.A(_0792_),
    .B(_0699_),
    .C(net53),
    .X(_0793_));
 sky130_fd_sc_hd__and3_2 _1451_ (.A(_0785_),
    .B(_0708_),
    .C(_0706_),
    .X(_0794_));
 sky130_fd_sc_hd__and4_1 _1452_ (.A(\RegFile.L[5] ),
    .B(_0789_),
    .C(_0699_),
    .D(net53),
    .X(_0795_));
 sky130_fd_sc_hd__a221o_1 _1453_ (.A1(\RegFile.C[5] ),
    .A2(_0793_),
    .B1(_0794_),
    .B2(\RegFile.B[5] ),
    .C1(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__or3_1 _1454_ (.A(\RegFile.A[5] ),
    .B(_0792_),
    .C(_0704_),
    .X(_0797_));
 sky130_fd_sc_hd__o31a_1 _1455_ (.A1(_0787_),
    .A2(_0791_),
    .A3(_0796_),
    .B1(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__a22o_1 _1456_ (.A1(\RegFile.C[5] ),
    .A2(_0705_),
    .B1(_0707_),
    .B2(\RegFile.L[5] ),
    .X(_0799_));
 sky130_fd_sc_hd__a31o_1 _1457_ (.A1(\RegFile.E[5] ),
    .A2(_0699_),
    .A3(net53),
    .B1(_0654_),
    .X(_0800_));
 sky130_fd_sc_hd__a211o_1 _1458_ (.A1(\ALU.flags_to_alu[5] ),
    .A2(_0711_),
    .B1(_0799_),
    .C1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__o211ai_4 _1459_ (.A1(_0630_),
    .A2(_0798_),
    .B1(_0801_),
    .C1(_0693_),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _1460_ (.A(_0782_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_1 _1461_ (.A(_0781_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__and2_1 _1462_ (.A(_0781_),
    .B(_0803_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_2 _1463_ (.A(_0804_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__and4_1 _1464_ (.A(\RegFile.C[2] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0807_));
 sky130_fd_sc_hd__and4_1 _1465_ (.A(\RegFile.L[2] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0762_),
    .X(_0808_));
 sky130_fd_sc_hd__a2111o_1 _1466_ (.A1(\RegFile.D[2] ),
    .A2(_0767_),
    .B1(_0807_),
    .C1(_0808_),
    .D1(net49),
    .X(_0809_));
 sky130_fd_sc_hd__a22o_1 _1467_ (.A1(\ALU.flags_to_alu[2] ),
    .A2(_0765_),
    .B1(_0763_),
    .B2(\RegFile.H[2] ),
    .X(_0810_));
 sky130_fd_sc_hd__a22o_1 _1468_ (.A1(\RegFile.E[2] ),
    .A2(_0761_),
    .B1(_0771_),
    .B2(\RegFile.B[2] ),
    .X(_0811_));
 sky130_fd_sc_hd__o32a_1 _1469_ (.A1(_0809_),
    .A2(_0810_),
    .A3(_0811_),
    .B1(_0774_),
    .B2(\RegFile.A[2] ),
    .X(_0812_));
 sky130_fd_sc_hd__a221o_1 _1470_ (.A1(\ALU.flags_to_alu[2] ),
    .A2(_0687_),
    .B1(_0683_),
    .B2(\RegFile.E[2] ),
    .C1(_0654_),
    .X(_0813_));
 sky130_fd_sc_hd__a22o_1 _1471_ (.A1(\RegFile.L[2] ),
    .A2(_0680_),
    .B1(_0685_),
    .B2(\RegFile.C[2] ),
    .X(_0814_));
 sky130_fd_sc_hd__o22a_4 _1472_ (.A1(_0629_),
    .A2(_0812_),
    .B1(_0813_),
    .B2(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nand2_8 _1473_ (.A(_0780_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__and3_2 _1474_ (.A(_0789_),
    .B(_0699_),
    .C(net53),
    .X(_0817_));
 sky130_fd_sc_hd__and4_1 _1475_ (.A(\RegFile.B[2] ),
    .B(_0785_),
    .C(_0708_),
    .D(_0706_),
    .X(_0818_));
 sky130_fd_sc_hd__a221o_1 _1476_ (.A1(\ALU.flags_to_alu[2] ),
    .A2(_0788_),
    .B1(_0817_),
    .B2(\RegFile.L[2] ),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__or2_1 _1477_ (.A(\RegFile.E[2] ),
    .B(_0789_),
    .X(_0820_));
 sky130_fd_sc_hd__a22o_1 _1478_ (.A1(\RegFile.H[2] ),
    .A2(_0784_),
    .B1(_0820_),
    .B2(_0711_),
    .X(_0821_));
 sky130_fd_sc_hd__a22o_1 _1479_ (.A1(\RegFile.C[2] ),
    .A2(_0793_),
    .B1(_0786_),
    .B2(\RegFile.D[2] ),
    .X(_0822_));
 sky130_fd_sc_hd__or3_1 _1480_ (.A(_0819_),
    .B(_0821_),
    .C(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__or3_1 _1481_ (.A(\RegFile.A[2] ),
    .B(_0792_),
    .C(_0704_),
    .X(_0824_));
 sky130_fd_sc_hd__o21a_1 _1482_ (.A1(\RegFile.E[2] ),
    .A2(_0703_),
    .B1(_0699_),
    .X(_0825_));
 sky130_fd_sc_hd__a221o_1 _1483_ (.A1(\RegFile.C[2] ),
    .A2(_0705_),
    .B1(_0707_),
    .B2(\RegFile.L[2] ),
    .C1(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__o211a_1 _1484_ (.A1(\ALU.flags_to_alu[2] ),
    .A2(_0704_),
    .B1(_0826_),
    .C1(_0629_),
    .X(_0827_));
 sky130_fd_sc_hd__or2_2 _1485_ (.A(_0664_),
    .B(_0692_),
    .X(_0828_));
 sky130_fd_sc_hd__a311o_1 _1486_ (.A1(_0654_),
    .A2(_0823_),
    .A3(_0824_),
    .B1(_0827_),
    .C1(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__inv_2 _1487_ (.A(_0664_),
    .Y(_0830_));
 sky130_fd_sc_hd__o211a_4 _1488_ (.A1(\ALU.immediate[2] ),
    .A2(_0674_),
    .B1(_0829_),
    .C1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__nor2_1 _1489_ (.A(_0816_),
    .B(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__and4_1 _1490_ (.A(\RegFile.B[3] ),
    .B(_0785_),
    .C(_0708_),
    .D(_0706_),
    .X(_0833_));
 sky130_fd_sc_hd__a221o_1 _1491_ (.A1(\ALU.flags_to_alu[3] ),
    .A2(_0788_),
    .B1(_0817_),
    .B2(\RegFile.L[3] ),
    .C1(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__or2_1 _1492_ (.A(\RegFile.E[3] ),
    .B(_0789_),
    .X(_0835_));
 sky130_fd_sc_hd__a22o_1 _1493_ (.A1(\RegFile.H[3] ),
    .A2(_0784_),
    .B1(_0835_),
    .B2(_0711_),
    .X(_0836_));
 sky130_fd_sc_hd__a22o_1 _1494_ (.A1(\RegFile.C[3] ),
    .A2(_0793_),
    .B1(_0786_),
    .B2(\RegFile.D[3] ),
    .X(_0837_));
 sky130_fd_sc_hd__or3_1 _1495_ (.A(_0834_),
    .B(_0836_),
    .C(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__or3_1 _1496_ (.A(\RegFile.A[3] ),
    .B(_0792_),
    .C(_0704_),
    .X(_0839_));
 sky130_fd_sc_hd__o21a_1 _1497_ (.A1(\RegFile.E[3] ),
    .A2(_0703_),
    .B1(_0699_),
    .X(_0840_));
 sky130_fd_sc_hd__a221o_1 _1498_ (.A1(\RegFile.C[3] ),
    .A2(_0705_),
    .B1(_0707_),
    .B2(\RegFile.L[3] ),
    .C1(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__o211a_1 _1499_ (.A1(\ALU.flags_to_alu[3] ),
    .A2(_0704_),
    .B1(_0841_),
    .C1(_0629_),
    .X(_0842_));
 sky130_fd_sc_hd__a311o_1 _1500_ (.A1(_0655_),
    .A2(_0838_),
    .A3(_0839_),
    .B1(_0842_),
    .C1(_0828_),
    .X(_0843_));
 sky130_fd_sc_hd__o211a_2 _1501_ (.A1(\ALU.immediate[3] ),
    .A2(_0674_),
    .B1(_0843_),
    .C1(_0830_),
    .X(_0844_));
 sky130_fd_sc_hd__and4_1 _1502_ (.A(\RegFile.C[3] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0845_));
 sky130_fd_sc_hd__and4_1 _1503_ (.A(\RegFile.L[3] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0762_),
    .X(_0846_));
 sky130_fd_sc_hd__a2111o_1 _1504_ (.A1(\RegFile.E[3] ),
    .A2(_0761_),
    .B1(_0845_),
    .C1(_0846_),
    .D1(net49),
    .X(_0847_));
 sky130_fd_sc_hd__a22o_1 _1505_ (.A1(\RegFile.D[3] ),
    .A2(_0767_),
    .B1(_0771_),
    .B2(\RegFile.B[3] ),
    .X(_0848_));
 sky130_fd_sc_hd__a22o_1 _1506_ (.A1(\ALU.flags_to_alu[3] ),
    .A2(_0765_),
    .B1(_0763_),
    .B2(\RegFile.H[3] ),
    .X(_0849_));
 sky130_fd_sc_hd__o32a_1 _1507_ (.A1(_0847_),
    .A2(_0848_),
    .A3(_0849_),
    .B1(_0774_),
    .B2(\RegFile.A[3] ),
    .X(_0850_));
 sky130_fd_sc_hd__a221o_1 _1508_ (.A1(\ALU.flags_to_alu[3] ),
    .A2(_0687_),
    .B1(_0683_),
    .B2(\RegFile.E[3] ),
    .C1(_0654_),
    .X(_0851_));
 sky130_fd_sc_hd__a22o_1 _1509_ (.A1(\RegFile.L[3] ),
    .A2(_0680_),
    .B1(_0685_),
    .B2(\RegFile.C[3] ),
    .X(_0852_));
 sky130_fd_sc_hd__o22a_1 _1510_ (.A1(_0629_),
    .A2(_0850_),
    .B1(_0851_),
    .B2(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__and2_1 _1511_ (.A(_0780_),
    .B(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_4 _1512_ (.A(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__and2b_1 _1513_ (.A_N(_0844_),
    .B(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__and4_1 _1514_ (.A(\RegFile.L[1] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0762_),
    .X(_0857_));
 sky130_fd_sc_hd__and4_1 _1515_ (.A(\RegFile.C[1] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0858_));
 sky130_fd_sc_hd__a2111o_1 _1516_ (.A1(\RegFile.D[1] ),
    .A2(_0767_),
    .B1(_0857_),
    .C1(_0858_),
    .D1(net49),
    .X(_0859_));
 sky130_fd_sc_hd__a22o_1 _1517_ (.A1(\RegFile.B[1] ),
    .A2(_0771_),
    .B1(_0763_),
    .B2(\RegFile.H[1] ),
    .X(_0860_));
 sky130_fd_sc_hd__a22o_1 _1518_ (.A1(\ALU.flags_to_alu[1] ),
    .A2(_0765_),
    .B1(_0761_),
    .B2(\RegFile.E[1] ),
    .X(_0861_));
 sky130_fd_sc_hd__nor3_1 _1519_ (.A(_0859_),
    .B(_0860_),
    .C(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__nor2_1 _1520_ (.A(\RegFile.A[1] ),
    .B(_0774_),
    .Y(_0863_));
 sky130_fd_sc_hd__a221o_1 _1521_ (.A1(\RegFile.E[1] ),
    .A2(_0683_),
    .B1(_0685_),
    .B2(\RegFile.C[1] ),
    .C1(_0687_),
    .X(_0864_));
 sky130_fd_sc_hd__a21oi_1 _1522_ (.A1(\RegFile.L[1] ),
    .A2(_0680_),
    .B1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__o21ai_1 _1523_ (.A1(\ALU.flags_to_alu[1] ),
    .A2(_0652_),
    .B1(_0629_),
    .Y(_0866_));
 sky130_fd_sc_hd__o32a_4 _1524_ (.A1(_0629_),
    .A2(_0862_),
    .A3(_0863_),
    .B1(_0865_),
    .B2(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__or2_1 _1525_ (.A(_0675_),
    .B(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__nand2_1 _1526_ (.A(\ALU.immediate[1] ),
    .B(_0675_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_1 _1527_ (.A(\RegFile.C[1] ),
    .B(_0793_),
    .Y(_0870_));
 sky130_fd_sc_hd__a22oi_1 _1528_ (.A1(\RegFile.H[1] ),
    .A2(_0784_),
    .B1(_0788_),
    .B2(\ALU.flags_to_alu[1] ),
    .Y(_0871_));
 sky130_fd_sc_hd__and4_1 _1529_ (.A(\RegFile.B[1] ),
    .B(_0785_),
    .C(_0708_),
    .D(_0706_),
    .X(_0872_));
 sky130_fd_sc_hd__and4_1 _1530_ (.A(\RegFile.D[1] ),
    .B(_0785_),
    .C(_0708_),
    .D(_0703_),
    .X(_0873_));
 sky130_fd_sc_hd__o211a_1 _1531_ (.A1(\RegFile.E[1] ),
    .A2(_0789_),
    .B1(_0699_),
    .C1(_0703_),
    .X(_0874_));
 sky130_fd_sc_hd__a2111oi_1 _1532_ (.A1(\RegFile.L[1] ),
    .A2(_0817_),
    .B1(_0872_),
    .C1(_0873_),
    .D1(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__a32o_1 _1533_ (.A1(_0870_),
    .A2(_0871_),
    .A3(_0875_),
    .B1(_0741_),
    .B2(_0789_),
    .X(_0876_));
 sky130_fd_sc_hd__and3_1 _1534_ (.A(\RegFile.E[1] ),
    .B(_0699_),
    .C(_0706_),
    .X(_0877_));
 sky130_fd_sc_hd__a221o_1 _1535_ (.A1(\RegFile.C[1] ),
    .A2(_0705_),
    .B1(_0707_),
    .B2(\RegFile.L[1] ),
    .C1(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__a211oi_1 _1536_ (.A1(\ALU.flags_to_alu[1] ),
    .A2(_0711_),
    .B1(_0878_),
    .C1(_0654_),
    .Y(_0879_));
 sky130_fd_sc_hd__a211o_2 _1537_ (.A1(_0654_),
    .A2(_0876_),
    .B1(_0879_),
    .C1(_0828_),
    .X(_0880_));
 sky130_fd_sc_hd__nand2_1 _1538_ (.A(_0869_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__or2_1 _1539_ (.A(_0868_),
    .B(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__or3_2 _1540_ (.A(_0675_),
    .B(_0867_),
    .C(_0880_),
    .X(_0883_));
 sky130_fd_sc_hd__o211ai_1 _1541_ (.A1(_0675_),
    .A2(_0867_),
    .B1(_0869_),
    .C1(_0880_),
    .Y(_0884_));
 sky130_fd_sc_hd__o21ai_4 _1542_ (.A1(\ALU.immediate[0] ),
    .A2(_0664_),
    .B1(_0692_),
    .Y(_0885_));
 sky130_fd_sc_hd__a22o_1 _1543_ (.A1(\RegFile.D[0] ),
    .A2(_0786_),
    .B1(_0794_),
    .B2(\RegFile.B[0] ),
    .X(_0886_));
 sky130_fd_sc_hd__and4_1 _1544_ (.A(\RegFile.C[0] ),
    .B(_0792_),
    .C(_0699_),
    .D(net53),
    .X(_0887_));
 sky130_fd_sc_hd__a221o_1 _1545_ (.A1(\RegFile.H[0] ),
    .A2(_0784_),
    .B1(_0788_),
    .B2(\ALU.flags_to_alu[0] ),
    .C1(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__or2_1 _1546_ (.A(\RegFile.E[0] ),
    .B(_0789_),
    .X(_0889_));
 sky130_fd_sc_hd__a22o_1 _1547_ (.A1(\RegFile.L[0] ),
    .A2(_0817_),
    .B1(_0889_),
    .B2(_0711_),
    .X(_0890_));
 sky130_fd_sc_hd__or3_1 _1548_ (.A(\RegFile.A[0] ),
    .B(_0792_),
    .C(_0704_),
    .X(_0891_));
 sky130_fd_sc_hd__o31a_1 _1549_ (.A1(_0886_),
    .A2(_0888_),
    .A3(_0890_),
    .B1(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__a22o_1 _1550_ (.A1(\RegFile.C[0] ),
    .A2(_0705_),
    .B1(_0709_),
    .B2(\RegFile.E[0] ),
    .X(_0893_));
 sky130_fd_sc_hd__a221o_1 _1551_ (.A1(\ALU.flags_to_alu[0] ),
    .A2(_0711_),
    .B1(_0707_),
    .B2(\RegFile.L[0] ),
    .C1(_0654_),
    .X(_0894_));
 sky130_fd_sc_hd__o21a_1 _1552_ (.A1(_0893_),
    .A2(_0894_),
    .B1(_0693_),
    .X(_0895_));
 sky130_fd_sc_hd__o21ai_4 _1553_ (.A1(_0629_),
    .A2(_0892_),
    .B1(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__and4_1 _1554_ (.A(\RegFile.C[0] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0897_));
 sky130_fd_sc_hd__a221o_1 _1555_ (.A1(\RegFile.L[0] ),
    .A2(_0770_),
    .B1(_0771_),
    .B2(\RegFile.B[0] ),
    .C1(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__o2111a_1 _1556_ (.A1(net54),
    .A2(_0650_),
    .B1(_0762_),
    .C1(_0638_),
    .D1(\RegFile.H[0] ),
    .X(_0899_));
 sky130_fd_sc_hd__o2111a_1 _1557_ (.A1(net54),
    .A2(_0650_),
    .B1(_0766_),
    .C1(_0684_),
    .D1(\RegFile.D[0] ),
    .X(_0900_));
 sky130_fd_sc_hd__o2111a_1 _1558_ (.A1(_0646_),
    .A2(_0650_),
    .B1(_0762_),
    .C1(_0684_),
    .D1(\ALU.flags_to_alu[0] ),
    .X(_0901_));
 sky130_fd_sc_hd__a2111o_1 _1559_ (.A1(\RegFile.E[0] ),
    .A2(_0761_),
    .B1(_0899_),
    .C1(_0900_),
    .D1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__a2111o_1 _1560_ (.A1(\RegFile.A[0] ),
    .A2(_0772_),
    .B1(_0898_),
    .C1(_0902_),
    .D1(_0629_),
    .X(_0903_));
 sky130_fd_sc_hd__a221o_1 _1561_ (.A1(\RegFile.E[0] ),
    .A2(_0683_),
    .B1(_0685_),
    .B2(\RegFile.C[0] ),
    .C1(_0654_),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _1562_ (.A1(\RegFile.L[0] ),
    .A2(_0680_),
    .B1(_0687_),
    .B2(\ALU.flags_to_alu[0] ),
    .X(_0905_));
 sky130_fd_sc_hd__or2_1 _1563_ (.A(_0904_),
    .B(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__and3_1 _1564_ (.A(_0780_),
    .B(_0903_),
    .C(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__buf_2 _1565_ (.A(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__a21oi_1 _1566_ (.A1(_0885_),
    .A2(_0896_),
    .B1(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21o_1 _1567_ (.A1(_0883_),
    .A2(_0884_),
    .B1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__xnor2_1 _1568_ (.A(_0816_),
    .B(_0831_),
    .Y(_0911_));
 sky130_fd_sc_hd__a21oi_2 _1569_ (.A1(_0882_),
    .A2(_0910_),
    .B1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__or2b_1 _1570_ (.A(_0855_),
    .B_N(_0844_),
    .X(_0913_));
 sky130_fd_sc_hd__a22o_1 _1571_ (.A1(\RegFile.E[4] ),
    .A2(_0761_),
    .B1(_0763_),
    .B2(\RegFile.H[4] ),
    .X(_0914_));
 sky130_fd_sc_hd__and4_1 _1572_ (.A(\RegFile.C[4] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0915_));
 sky130_fd_sc_hd__a221o_1 _1573_ (.A1(\ALU.flags_to_alu[4] ),
    .A2(_0765_),
    .B1(_0767_),
    .B2(\RegFile.D[4] ),
    .C1(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__a221o_1 _1574_ (.A1(\RegFile.L[4] ),
    .A2(_0770_),
    .B1(_0771_),
    .B2(\RegFile.B[4] ),
    .C1(net50),
    .X(_0917_));
 sky130_fd_sc_hd__o32a_1 _1575_ (.A1(_0914_),
    .A2(_0916_),
    .A3(_0917_),
    .B1(_0774_),
    .B2(\RegFile.A[4] ),
    .X(_0918_));
 sky130_fd_sc_hd__a221o_1 _1576_ (.A1(\ALU.flags_to_alu[4] ),
    .A2(_0687_),
    .B1(_0683_),
    .B2(\RegFile.E[4] ),
    .C1(_0654_),
    .X(_0919_));
 sky130_fd_sc_hd__a22o_1 _1577_ (.A1(\RegFile.L[4] ),
    .A2(net52),
    .B1(net51),
    .B2(\RegFile.C[4] ),
    .X(_0920_));
 sky130_fd_sc_hd__o22a_2 _1578_ (.A1(_0629_),
    .A2(_0918_),
    .B1(_0919_),
    .B2(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__nand2_2 _1579_ (.A(_0780_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__or3_1 _1580_ (.A(\RegFile.A[4] ),
    .B(_0792_),
    .C(_0704_),
    .X(_0923_));
 sky130_fd_sc_hd__a22o_1 _1581_ (.A1(\RegFile.H[4] ),
    .A2(_0784_),
    .B1(_0786_),
    .B2(\RegFile.D[4] ),
    .X(_0924_));
 sky130_fd_sc_hd__a22o_1 _1582_ (.A1(\RegFile.C[4] ),
    .A2(_0793_),
    .B1(_0794_),
    .B2(\RegFile.B[4] ),
    .X(_0925_));
 sky130_fd_sc_hd__or2_1 _1583_ (.A(\RegFile.E[4] ),
    .B(_0789_),
    .X(_0926_));
 sky130_fd_sc_hd__a22o_1 _1584_ (.A1(\ALU.flags_to_alu[4] ),
    .A2(_0788_),
    .B1(_0926_),
    .B2(_0711_),
    .X(_0927_));
 sky130_fd_sc_hd__a2111o_1 _1585_ (.A1(\RegFile.L[4] ),
    .A2(_0817_),
    .B1(_0924_),
    .C1(_0925_),
    .D1(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__a21o_1 _1586_ (.A1(_0923_),
    .A2(_0928_),
    .B1(_0629_),
    .X(_0929_));
 sky130_fd_sc_hd__and3_1 _1587_ (.A(\ALU.flags_to_alu[4] ),
    .B(_0699_),
    .C(_0703_),
    .X(_0930_));
 sky130_fd_sc_hd__a22o_1 _1588_ (.A1(\RegFile.C[4] ),
    .A2(_0705_),
    .B1(_0707_),
    .B2(\RegFile.L[4] ),
    .X(_0931_));
 sky130_fd_sc_hd__a31o_1 _1589_ (.A1(\RegFile.E[4] ),
    .A2(_0699_),
    .A3(net53),
    .B1(_0654_),
    .X(_0932_));
 sky130_fd_sc_hd__o31a_1 _1590_ (.A1(_0930_),
    .A2(_0931_),
    .A3(_0932_),
    .B1(_0693_),
    .X(_0933_));
 sky130_fd_sc_hd__a22o_1 _1591_ (.A1(\ALU.immediate[4] ),
    .A2(_0675_),
    .B1(_0929_),
    .B2(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__nor2_1 _1592_ (.A(_0922_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__and2_1 _1593_ (.A(_0922_),
    .B(_0934_),
    .X(_0936_));
 sky130_fd_sc_hd__nor2_2 _1594_ (.A(_0935_),
    .B(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__o311a_1 _1595_ (.A1(_0832_),
    .A2(_0856_),
    .A3(_0912_),
    .B1(_0913_),
    .C1(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__a22o_1 _1596_ (.A1(\RegFile.E[7] ),
    .A2(_0761_),
    .B1(_0771_),
    .B2(\RegFile.B[7] ),
    .X(_0939_));
 sky130_fd_sc_hd__and4_1 _1597_ (.A(\RegFile.C[7] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0940_));
 sky130_fd_sc_hd__a221o_1 _1598_ (.A1(\ALU.flags_to_alu[7] ),
    .A2(_0765_),
    .B1(_0767_),
    .B2(\RegFile.D[7] ),
    .C1(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__a221o_1 _1599_ (.A1(\RegFile.L[7] ),
    .A2(_0770_),
    .B1(_0763_),
    .B2(\RegFile.H[7] ),
    .C1(net50),
    .X(_0942_));
 sky130_fd_sc_hd__o32a_1 _1600_ (.A1(_0939_),
    .A2(_0941_),
    .A3(_0942_),
    .B1(_0774_),
    .B2(\RegFile.A[7] ),
    .X(_0943_));
 sky130_fd_sc_hd__a221o_1 _1601_ (.A1(\ALU.flags_to_alu[7] ),
    .A2(_0687_),
    .B1(_0683_),
    .B2(\RegFile.E[7] ),
    .C1(_0654_),
    .X(_0944_));
 sky130_fd_sc_hd__a22o_1 _1602_ (.A1(\RegFile.L[7] ),
    .A2(net52),
    .B1(net51),
    .B2(\RegFile.C[7] ),
    .X(_0945_));
 sky130_fd_sc_hd__o22a_2 _1603_ (.A1(_0629_),
    .A2(_0943_),
    .B1(_0944_),
    .B2(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__nand2_4 _1604_ (.A(_0780_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__or3_1 _1605_ (.A(\RegFile.A[7] ),
    .B(_0792_),
    .C(_0704_),
    .X(_0948_));
 sky130_fd_sc_hd__and2_1 _1606_ (.A(\ALU.flags_to_alu[7] ),
    .B(_0788_),
    .X(_0949_));
 sky130_fd_sc_hd__a22o_1 _1607_ (.A1(\RegFile.C[7] ),
    .A2(_0793_),
    .B1(_0786_),
    .B2(\RegFile.D[7] ),
    .X(_0950_));
 sky130_fd_sc_hd__or2_1 _1608_ (.A(\RegFile.E[7] ),
    .B(_0789_),
    .X(_0951_));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(\RegFile.B[7] ),
    .A2(_0794_),
    .B1(_0951_),
    .B2(_0711_),
    .X(_0952_));
 sky130_fd_sc_hd__a22o_1 _1610_ (.A1(\RegFile.H[7] ),
    .A2(_0784_),
    .B1(_0817_),
    .B2(\RegFile.L[7] ),
    .X(_0953_));
 sky130_fd_sc_hd__or4_1 _1611_ (.A(_0949_),
    .B(_0950_),
    .C(_0952_),
    .D(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__a21o_1 _1612_ (.A1(_0948_),
    .A2(_0954_),
    .B1(_0629_),
    .X(_0955_));
 sky130_fd_sc_hd__and3_1 _1613_ (.A(\RegFile.C[7] ),
    .B(_0708_),
    .C(net53),
    .X(_0956_));
 sky130_fd_sc_hd__a221o_1 _1614_ (.A1(\ALU.flags_to_alu[7] ),
    .A2(_0711_),
    .B1(_0707_),
    .B2(\RegFile.L[7] ),
    .C1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__a211o_1 _1615_ (.A1(\RegFile.E[7] ),
    .A2(_0709_),
    .B1(_0957_),
    .C1(_0654_),
    .X(_0958_));
 sky130_fd_sc_hd__a32o_2 _1616_ (.A1(_0955_),
    .A2(_0693_),
    .A3(_0958_),
    .B1(_0675_),
    .B2(\ALU.immediate[7] ),
    .X(_0959_));
 sky130_fd_sc_hd__xnor2_4 _1617_ (.A(_0947_),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__a22oi_1 _1618_ (.A1(\RegFile.E[6] ),
    .A2(_0761_),
    .B1(_0771_),
    .B2(\RegFile.B[6] ),
    .Y(_0961_));
 sky130_fd_sc_hd__and4_1 _1619_ (.A(\RegFile.C[6] ),
    .B(_0638_),
    .C(_0681_),
    .D(_0760_),
    .X(_0962_));
 sky130_fd_sc_hd__a221oi_1 _1620_ (.A1(\ALU.flags_to_alu[6] ),
    .A2(_0765_),
    .B1(_0767_),
    .B2(\RegFile.D[6] ),
    .C1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__a221oi_1 _1621_ (.A1(\RegFile.L[6] ),
    .A2(_0770_),
    .B1(_0763_),
    .B2(\RegFile.H[6] ),
    .C1(net50),
    .Y(_0964_));
 sky130_fd_sc_hd__inv_2 _1622_ (.A(\RegFile.A[6] ),
    .Y(_0965_));
 sky130_fd_sc_hd__a32o_1 _1623_ (.A1(_0961_),
    .A2(_0963_),
    .A3(_0964_),
    .B1(net49),
    .B2(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__a221o_1 _1624_ (.A1(\ALU.flags_to_alu[6] ),
    .A2(_0687_),
    .B1(_0683_),
    .B2(\RegFile.E[6] ),
    .C1(_0654_),
    .X(_0967_));
 sky130_fd_sc_hd__a22o_1 _1625_ (.A1(\RegFile.L[6] ),
    .A2(_0680_),
    .B1(_0685_),
    .B2(\RegFile.C[6] ),
    .X(_0968_));
 sky130_fd_sc_hd__o2bb2a_2 _1626_ (.A1_N(_0654_),
    .A2_N(_0966_),
    .B1(_0967_),
    .B2(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__nand2_2 _1627_ (.A(_0780_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__or3_1 _1628_ (.A(\RegFile.A[6] ),
    .B(_0792_),
    .C(_0704_),
    .X(_0971_));
 sky130_fd_sc_hd__and2_1 _1629_ (.A(\ALU.flags_to_alu[6] ),
    .B(_0788_),
    .X(_0972_));
 sky130_fd_sc_hd__a22o_1 _1630_ (.A1(\RegFile.C[6] ),
    .A2(_0793_),
    .B1(_0786_),
    .B2(\RegFile.D[6] ),
    .X(_0973_));
 sky130_fd_sc_hd__or2_1 _1631_ (.A(\RegFile.E[6] ),
    .B(_0789_),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _1632_ (.A1(\RegFile.B[6] ),
    .A2(_0794_),
    .B1(_0974_),
    .B2(_0711_),
    .X(_0975_));
 sky130_fd_sc_hd__a22o_1 _1633_ (.A1(\RegFile.H[6] ),
    .A2(_0784_),
    .B1(_0817_),
    .B2(\RegFile.L[6] ),
    .X(_0976_));
 sky130_fd_sc_hd__or4_1 _1634_ (.A(_0972_),
    .B(_0973_),
    .C(_0975_),
    .D(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__a21o_1 _1635_ (.A1(_0971_),
    .A2(_0977_),
    .B1(_0629_),
    .X(_0978_));
 sky130_fd_sc_hd__a22o_1 _1636_ (.A1(\RegFile.C[6] ),
    .A2(_0705_),
    .B1(_0707_),
    .B2(\RegFile.L[6] ),
    .X(_0979_));
 sky130_fd_sc_hd__a221o_1 _1637_ (.A1(\ALU.flags_to_alu[6] ),
    .A2(_0711_),
    .B1(_0709_),
    .B2(\RegFile.E[6] ),
    .C1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__or2_1 _1638_ (.A(_0655_),
    .B(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__a32o_4 _1639_ (.A1(_0693_),
    .A2(_0978_),
    .A3(_0981_),
    .B1(_0675_),
    .B2(\ALU.immediate[6] ),
    .X(_0982_));
 sky130_fd_sc_hd__xnor2_2 _1640_ (.A(_0970_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__nor2_1 _1641_ (.A(_0960_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__o21ba_1 _1642_ (.A1(_0804_),
    .A2(_0935_),
    .B1_N(_0805_),
    .X(_0985_));
 sky130_fd_sc_hd__and2_1 _1643_ (.A(_0947_),
    .B(_0959_),
    .X(_0986_));
 sky130_fd_sc_hd__or2_1 _1644_ (.A(_0947_),
    .B(_0959_),
    .X(_0987_));
 sky130_fd_sc_hd__o31a_1 _1645_ (.A1(_0986_),
    .A2(_0970_),
    .A3(_0982_),
    .B1(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__a21bo_1 _1646_ (.A1(_0984_),
    .A2(_0985_),
    .B1_N(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__a31o_1 _1647_ (.A1(_0806_),
    .A2(_0938_),
    .A3(_0984_),
    .B1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__nor2_1 _1648_ (.A(_0740_),
    .B(_0745_),
    .Y(_0991_));
 sky130_fd_sc_hd__inv_2 _1649_ (.A(_0749_),
    .Y(_0992_));
 sky130_fd_sc_hd__nor2_1 _1650_ (.A(_0992_),
    .B(_0753_),
    .Y(_0993_));
 sky130_fd_sc_hd__a211o_1 _1651_ (.A1(_0756_),
    .A2(_0990_),
    .B1(_0991_),
    .C1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__inv_2 _1652_ (.A(_0729_),
    .Y(_0995_));
 sky130_fd_sc_hd__nor2_1 _1653_ (.A(_0995_),
    .B(_0733_),
    .Y(_0996_));
 sky130_fd_sc_hd__a31o_1 _1654_ (.A1(_0737_),
    .A2(_0746_),
    .A3(_0994_),
    .B1(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__inv_2 _1655_ (.A(_0721_),
    .Y(_0998_));
 sky130_fd_sc_hd__nor2_1 _1656_ (.A(_0998_),
    .B(_0725_),
    .Y(_0999_));
 sky130_fd_sc_hd__a21oi_1 _1657_ (.A1(_0726_),
    .A2(_0997_),
    .B1(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__a221o_1 _1658_ (.A1(\RegFile.D[5] ),
    .A2(_0683_),
    .B1(net51),
    .B2(\RegFile.B[5] ),
    .C1(_0687_),
    .X(_1001_));
 sky130_fd_sc_hd__a21o_1 _1659_ (.A1(\RegFile.H[5] ),
    .A2(net52),
    .B1(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__o211a_1 _1660_ (.A1(\RegFile.A[5] ),
    .A2(_0652_),
    .B1(_0676_),
    .C1(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__a22o_1 _1661_ (.A1(\RegFile.H[5] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[5] ),
    .X(_1004_));
 sky130_fd_sc_hd__a211o_1 _1662_ (.A1(\RegFile.B[5] ),
    .A2(_0705_),
    .B1(_1004_),
    .C1(_0711_),
    .X(_1005_));
 sky130_fd_sc_hd__o211a_1 _1663_ (.A1(\RegFile.A[5] ),
    .A2(_0704_),
    .B1(_1005_),
    .C1(_0630_),
    .X(_1006_));
 sky130_fd_sc_hd__a22o_1 _1664_ (.A1(\ALU.immediate[13] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__nand2_1 _1665_ (.A(_1003_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__inv_2 _1666_ (.A(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__nor2_1 _1667_ (.A(_1003_),
    .B(_1007_),
    .Y(_1010_));
 sky130_fd_sc_hd__nor2_1 _1668_ (.A(_1009_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__a221o_1 _1669_ (.A1(\RegFile.D[4] ),
    .A2(_0683_),
    .B1(net51),
    .B2(\RegFile.B[4] ),
    .C1(_0687_),
    .X(_1012_));
 sky130_fd_sc_hd__a21o_1 _1670_ (.A1(\RegFile.H[4] ),
    .A2(net52),
    .B1(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__o211ai_2 _1671_ (.A1(\RegFile.A[4] ),
    .A2(_0652_),
    .B1(_0676_),
    .C1(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__a22o_1 _1672_ (.A1(\RegFile.H[4] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[4] ),
    .X(_1015_));
 sky130_fd_sc_hd__a211o_1 _1673_ (.A1(\RegFile.B[4] ),
    .A2(_0705_),
    .B1(_1015_),
    .C1(_0711_),
    .X(_1016_));
 sky130_fd_sc_hd__o211a_1 _1674_ (.A1(\RegFile.A[4] ),
    .A2(_0704_),
    .B1(_1016_),
    .C1(_0630_),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_1 _1675_ (.A1(\ALU.immediate[12] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(_1014_),
    .B(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__inv_2 _1677_ (.A(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__nand2_1 _1678_ (.A(_1014_),
    .B(_1018_),
    .Y(_1021_));
 sky130_fd_sc_hd__nand2_1 _1679_ (.A(_1020_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__inv_2 _1680_ (.A(_1003_),
    .Y(_1023_));
 sky130_fd_sc_hd__o22a_1 _1681_ (.A1(_1023_),
    .A2(_1007_),
    .B1(_1011_),
    .B2(_1020_),
    .X(_1024_));
 sky130_fd_sc_hd__o31a_1 _1682_ (.A1(_1000_),
    .A2(_1011_),
    .A3(_1022_),
    .B1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__nor2_1 _1683_ (.A(_0718_),
    .B(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__a221o_1 _1684_ (.A1(\RegFile.D[7] ),
    .A2(_0683_),
    .B1(net51),
    .B2(\RegFile.B[7] ),
    .C1(_0687_),
    .X(_1027_));
 sky130_fd_sc_hd__a21o_1 _1685_ (.A1(\RegFile.H[7] ),
    .A2(net52),
    .B1(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__o211a_1 _1686_ (.A1(\RegFile.A[7] ),
    .A2(_0652_),
    .B1(_1028_),
    .C1(_0676_),
    .X(_1029_));
 sky130_fd_sc_hd__a22o_1 _1687_ (.A1(\RegFile.H[7] ),
    .A2(_0707_),
    .B1(_0709_),
    .B2(\RegFile.D[7] ),
    .X(_1030_));
 sky130_fd_sc_hd__a211o_1 _1688_ (.A1(\RegFile.B[7] ),
    .A2(_0705_),
    .B1(_1030_),
    .C1(_0711_),
    .X(_1031_));
 sky130_fd_sc_hd__o211a_1 _1689_ (.A1(\RegFile.A[7] ),
    .A2(_0704_),
    .B1(_1031_),
    .C1(_0630_),
    .X(_1032_));
 sky130_fd_sc_hd__a22o_1 _1690_ (.A1(\ALU.immediate[15] ),
    .A2(_0675_),
    .B1(_0693_),
    .B2(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__nand2_1 _1691_ (.A(_1029_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__nor2_1 _1692_ (.A(_1029_),
    .B(_1033_),
    .Y(_1035_));
 sky130_fd_sc_hd__inv_2 _1693_ (.A(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__nand2_1 _1694_ (.A(_1034_),
    .B(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__o21a_1 _1695_ (.A1(_0715_),
    .A2(_1026_),
    .B1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__and3_1 _1696_ (.A(\ByteBuffer.instr[20] ),
    .B(_0622_),
    .C(_0624_),
    .X(_1039_));
 sky130_fd_sc_hd__a221o_1 _1697_ (.A1(_0619_),
    .A2(_0620_),
    .B1(_0647_),
    .B2(\ByteBuffer.instr[19] ),
    .C1(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__o211a_1 _1698_ (.A1(_0622_),
    .A2(_0624_),
    .B1(_0621_),
    .C1(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__a221o_1 _1699_ (.A1(\ByteBuffer.instr[20] ),
    .A2(_0645_),
    .B1(_0672_),
    .B2(_1041_),
    .C1(_0648_),
    .X(_1042_));
 sky130_fd_sc_hd__o21ai_4 _1700_ (.A1(_0678_),
    .A2(_1039_),
    .B1(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__and3b_2 _1701_ (.A_N(_0656_),
    .B(_0700_),
    .C(_0624_),
    .X(_1044_));
 sky130_fd_sc_hd__a21o_1 _1702_ (.A1(_0622_),
    .A2(_0624_),
    .B1(_0678_),
    .X(_1045_));
 sky130_fd_sc_hd__o211a_1 _1703_ (.A1(_0645_),
    .A2(_1044_),
    .B1(_1045_),
    .C1(\ByteBuffer.instr[21] ),
    .X(_1046_));
 sky130_fd_sc_hd__a21oi_4 _1704_ (.A1(_0670_),
    .A2(_1044_),
    .B1(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__o211ai_4 _1705_ (.A1(_0645_),
    .A2(_1044_),
    .B1(_1045_),
    .C1(\ByteBuffer.instr[19] ),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_8 _1706_ (.A(_1047_),
    .B(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__nor2_2 _1707_ (.A(net48),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__o31ai_2 _1708_ (.A1(_1037_),
    .A2(_0715_),
    .A3(_1026_),
    .B1(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__inv_2 _1709_ (.A(_0726_),
    .Y(_1052_));
 sky130_fd_sc_hd__inv_2 _1710_ (.A(_0991_),
    .Y(_1053_));
 sky130_fd_sc_hd__nand2_1 _1711_ (.A(_0746_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__inv_2 _1712_ (.A(_0756_),
    .Y(_1055_));
 sky130_fd_sc_hd__nor2_1 _1713_ (.A(_0855_),
    .B(_0844_),
    .Y(_1056_));
 sky130_fd_sc_hd__xor2_4 _1714_ (.A(_0816_),
    .B(_0831_),
    .X(_1057_));
 sky130_fd_sc_hd__o211a_1 _1715_ (.A1(_0675_),
    .A2(_0867_),
    .B1(_0869_),
    .C1(_0880_),
    .X(_1058_));
 sky130_fd_sc_hd__a21bo_1 _1716_ (.A1(_0885_),
    .A2(_0896_),
    .B1_N(_0908_),
    .X(_1059_));
 sky130_fd_sc_hd__o21a_2 _1717_ (.A1(_1058_),
    .A2(_1059_),
    .B1(_0883_),
    .X(_1060_));
 sky130_fd_sc_hd__nand2_1 _1718_ (.A(_0855_),
    .B(_0844_),
    .Y(_1061_));
 sky130_fd_sc_hd__or2b_1 _1719_ (.A(_0816_),
    .B_N(_0831_),
    .X(_1062_));
 sky130_fd_sc_hd__o211a_1 _1720_ (.A1(_1057_),
    .A2(_1060_),
    .B1(_1061_),
    .C1(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__nor2_1 _1721_ (.A(_1056_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__nor2_1 _1722_ (.A(_0806_),
    .B(_0937_),
    .Y(_1065_));
 sky130_fd_sc_hd__and2_1 _1723_ (.A(_0780_),
    .B(_0946_),
    .X(_1066_));
 sky130_fd_sc_hd__nand2_1 _1724_ (.A(_1066_),
    .B(_0959_),
    .Y(_1067_));
 sky130_fd_sc_hd__and2_1 _1725_ (.A(_0780_),
    .B(_0969_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_2 _1726_ (.A(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__nand2_1 _1727_ (.A(_1069_),
    .B(_0982_),
    .Y(_1070_));
 sky130_fd_sc_hd__a21o_1 _1728_ (.A1(_0782_),
    .A2(_0802_),
    .B1(_0781_),
    .X(_1071_));
 sky130_fd_sc_hd__nand4_2 _1729_ (.A(_0780_),
    .B(_0921_),
    .C(_0929_),
    .D(_0933_),
    .Y(_1072_));
 sky130_fd_sc_hd__and3_1 _1730_ (.A(_0781_),
    .B(_0782_),
    .C(_0802_),
    .X(_1073_));
 sky130_fd_sc_hd__a21o_1 _1731_ (.A1(_1071_),
    .A2(_1072_),
    .B1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__nor2_1 _1732_ (.A(_1066_),
    .B(_0959_),
    .Y(_1075_));
 sky130_fd_sc_hd__nor2_1 _1733_ (.A(_1069_),
    .B(_0982_),
    .Y(_1076_));
 sky130_fd_sc_hd__a211o_1 _1734_ (.A1(_1070_),
    .A2(_1074_),
    .B1(_1075_),
    .C1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_1 _1735_ (.A(_1067_),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__a41o_1 _1736_ (.A1(_0960_),
    .A2(_0983_),
    .A3(_1064_),
    .A4(_1065_),
    .B1(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__a21bo_1 _1737_ (.A1(_1055_),
    .A2(_1079_),
    .B1_N(_0754_),
    .X(_1080_));
 sky130_fd_sc_hd__and2b_1 _1738_ (.A_N(_0740_),
    .B(_0745_),
    .X(_1081_));
 sky130_fd_sc_hd__a21o_1 _1739_ (.A1(_1054_),
    .A2(_1080_),
    .B1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__a22o_1 _1740_ (.A1(_0721_),
    .A2(_0725_),
    .B1(_0729_),
    .B2(_0733_),
    .X(_1083_));
 sky130_fd_sc_hd__o21a_1 _1741_ (.A1(_0721_),
    .A2(_0725_),
    .B1(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__a31o_1 _1742_ (.A1(_1052_),
    .A2(_0736_),
    .A3(_1082_),
    .B1(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__or2b_1 _1743_ (.A(_1014_),
    .B_N(_1018_),
    .X(_1086_));
 sky130_fd_sc_hd__a21oi_1 _1744_ (.A1(_1008_),
    .A2(_1086_),
    .B1(_1010_),
    .Y(_1087_));
 sky130_fd_sc_hd__a31o_1 _1745_ (.A1(_1011_),
    .A2(_1022_),
    .A3(_1085_),
    .B1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__a21oi_1 _1746_ (.A1(_0718_),
    .A2(_1088_),
    .B1(_0716_),
    .Y(_1089_));
 sky130_fd_sc_hd__xnor2_1 _1747_ (.A(_1037_),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__and2_1 _1748_ (.A(_1047_),
    .B(_1048_),
    .X(_1091_));
 sky130_fd_sc_hd__buf_6 _1749_ (.A(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__nand2_4 _1750_ (.A(net48),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__o22ai_4 _1751_ (.A1(_1038_),
    .A2(_1051_),
    .B1(_1090_),
    .B2(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__nand2_1 _1752_ (.A(_0970_),
    .B(_0982_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _1753_ (.A(_0960_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__or2_1 _1754_ (.A(_0960_),
    .B(_1095_),
    .X(_1097_));
 sky130_fd_sc_hd__and2_1 _1755_ (.A(_1096_),
    .B(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__or2_1 _1756_ (.A(_0970_),
    .B(_0982_),
    .X(_1099_));
 sky130_fd_sc_hd__and2_1 _1757_ (.A(_1099_),
    .B(_1095_),
    .X(_1100_));
 sky130_fd_sc_hd__nor2_1 _1758_ (.A(_1100_),
    .B(_0805_),
    .Y(_1101_));
 sky130_fd_sc_hd__and2_1 _1759_ (.A(_1100_),
    .B(_0805_),
    .X(_1102_));
 sky130_fd_sc_hd__nor2_1 _1760_ (.A(_1101_),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__and2b_1 _1761_ (.A_N(_0855_),
    .B(_0844_),
    .X(_1104_));
 sky130_fd_sc_hd__or2_1 _1762_ (.A(_0937_),
    .B(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__nand2_1 _1763_ (.A(_0816_),
    .B(_0831_),
    .Y(_1106_));
 sky130_fd_sc_hd__nand2_1 _1764_ (.A(_0868_),
    .B(_0881_),
    .Y(_1107_));
 sky130_fd_sc_hd__a21o_1 _1765_ (.A1(_0885_),
    .A2(_0896_),
    .B1(_0908_),
    .X(_1108_));
 sky130_fd_sc_hd__inv_2 _1766_ (.A(\ALU.flags_to_alu[0] ),
    .Y(_1109_));
 sky130_fd_sc_hd__a31o_1 _1767_ (.A1(_0908_),
    .A2(_0885_),
    .A3(_0896_),
    .B1(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__a2bb2o_1 _1768_ (.A1_N(_0868_),
    .A2_N(_0881_),
    .B1(_1108_),
    .B2(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__a21o_1 _1769_ (.A1(_1107_),
    .A2(_1111_),
    .B1(_0832_),
    .X(_1112_));
 sky130_fd_sc_hd__nor2_2 _1770_ (.A(_1104_),
    .B(_0856_),
    .Y(_1113_));
 sky130_fd_sc_hd__a21bo_1 _1771_ (.A1(_1106_),
    .A2(_1112_),
    .B1_N(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__xnor2_1 _1772_ (.A(_0937_),
    .B(_0913_),
    .Y(_1115_));
 sky130_fd_sc_hd__nand2_1 _1773_ (.A(_1114_),
    .B(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__xnor2_1 _1774_ (.A(_0806_),
    .B(_0936_),
    .Y(_1117_));
 sky130_fd_sc_hd__a21oi_1 _1775_ (.A1(_1105_),
    .A2(_1116_),
    .B1(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__o21bai_1 _1776_ (.A1(_0806_),
    .A2(_0936_),
    .B1_N(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__and2_1 _1777_ (.A(_1103_),
    .B(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__or3_1 _1778_ (.A(_1098_),
    .B(_1101_),
    .C(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__o211a_2 _1779_ (.A1(_0645_),
    .A2(_1044_),
    .B1(_1045_),
    .C1(\ByteBuffer.instr[19] ),
    .X(_1122_));
 sky130_fd_sc_hd__nand2_2 _1780_ (.A(_1047_),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__nor2_2 _1781_ (.A(_1043_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__o21ai_1 _1782_ (.A1(_1101_),
    .A2(_1120_),
    .B1(_1098_),
    .Y(_1125_));
 sky130_fd_sc_hd__and3_1 _1783_ (.A(_1121_),
    .B(_1124_),
    .C(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__or3_2 _1784_ (.A(_0937_),
    .B(_1056_),
    .C(_1063_),
    .X(_1127_));
 sky130_fd_sc_hd__o21a_1 _1785_ (.A1(_0806_),
    .A2(_1127_),
    .B1(_1074_),
    .X(_1128_));
 sky130_fd_sc_hd__o21ai_1 _1786_ (.A1(_1100_),
    .A2(_1128_),
    .B1(_1070_),
    .Y(_1129_));
 sky130_fd_sc_hd__xnor2_1 _1787_ (.A(_0960_),
    .B(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__xnor2_1 _1788_ (.A(_0983_),
    .B(_1128_),
    .Y(_1131_));
 sky130_fd_sc_hd__inv_2 _1789_ (.A(_0806_),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_1 _1790_ (.A(_1072_),
    .B(_1127_),
    .Y(_1133_));
 sky130_fd_sc_hd__xnor2_2 _1791_ (.A(_1132_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__or3_1 _1792_ (.A(_0935_),
    .B(_0936_),
    .C(_1064_),
    .X(_1135_));
 sky130_fd_sc_hd__nand2_2 _1793_ (.A(_1127_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__xnor2_2 _1794_ (.A(_1057_),
    .B(_1060_),
    .Y(_1137_));
 sky130_fd_sc_hd__and2_1 _1795_ (.A(_0883_),
    .B(_0884_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_2 _1796_ (.A(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__nand3b_1 _1797_ (.A_N(_0908_),
    .B(_0885_),
    .C(_0896_),
    .Y(_1140_));
 sky130_fd_sc_hd__and3_1 _1798_ (.A(\ALU.flags_to_alu[0] ),
    .B(_1059_),
    .C(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__nand2_1 _1799_ (.A(_1139_),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__nor2_1 _1800_ (.A(_1137_),
    .B(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__o21ai_1 _1801_ (.A1(_1057_),
    .A2(_1060_),
    .B1(_1062_),
    .Y(_1144_));
 sky130_fd_sc_hd__xnor2_1 _1802_ (.A(_1144_),
    .B(_1113_),
    .Y(_1145_));
 sky130_fd_sc_hd__nand2_1 _1803_ (.A(_1143_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__nor3_2 _1804_ (.A(_1134_),
    .B(_1136_),
    .C(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(_1131_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__nor2_1 _1806_ (.A(_1130_),
    .B(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__o21a_1 _1807_ (.A1(_0678_),
    .A2(_1039_),
    .B1(_1042_),
    .X(_1150_));
 sky130_fd_sc_hd__buf_6 _1808_ (.A(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__a2111oi_1 _1809_ (.A1(_1130_),
    .A2(_1148_),
    .B1(_1149_),
    .C1(_1151_),
    .D1(_1123_),
    .Y(_1152_));
 sky130_fd_sc_hd__inv_2 _1810_ (.A(_0982_),
    .Y(_1153_));
 sky130_fd_sc_hd__nor2_1 _1811_ (.A(_0935_),
    .B(_0938_),
    .Y(_1154_));
 sky130_fd_sc_hd__o21ba_1 _1812_ (.A1(_1132_),
    .A2(_1154_),
    .B1_N(_0804_),
    .X(_1155_));
 sky130_fd_sc_hd__nor2_1 _1813_ (.A(_0983_),
    .B(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__a21o_1 _1814_ (.A1(_1069_),
    .A2(_1153_),
    .B1(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__xnor2_1 _1815_ (.A(_0960_),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__and3_1 _1816_ (.A(\ByteBuffer.instr[21] ),
    .B(_0645_),
    .C(_1045_),
    .X(_1159_));
 sky130_fd_sc_hd__and2_2 _1817_ (.A(_1122_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__o21a_1 _1818_ (.A1(_1092_),
    .A2(_1160_),
    .B1(_1151_),
    .X(_1161_));
 sky130_fd_sc_hd__and2_1 _1819_ (.A(_1043_),
    .B(_1160_),
    .X(_1162_));
 sky130_fd_sc_hd__or3b_2 _1820_ (.A(\ByteBuffer.instr[21] ),
    .B(_0645_),
    .C_N(_1044_),
    .X(_1163_));
 sky130_fd_sc_hd__nor2_2 _1821_ (.A(_1122_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__nor2_2 _1822_ (.A(_1048_),
    .B(_1163_),
    .Y(_1165_));
 sky130_fd_sc_hd__nor2_4 _1823_ (.A(_1151_),
    .B(_1049_),
    .Y(_1166_));
 sky130_fd_sc_hd__a31o_1 _1824_ (.A1(\ALU.flags_to_alu[0] ),
    .A2(_1151_),
    .A3(_1165_),
    .B1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__or3b_4 _1825_ (.A(_1043_),
    .B(_1122_),
    .C_N(_1159_),
    .X(_1168_));
 sky130_fd_sc_hd__nor2_1 _1826_ (.A(_1075_),
    .B(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__a211o_1 _1827_ (.A1(_1069_),
    .A2(_1164_),
    .B1(_1167_),
    .C1(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__or3b_1 _1828_ (.A(_1151_),
    .B(_1122_),
    .C_N(_1159_),
    .X(_1171_));
 sky130_fd_sc_hd__buf_2 _1829_ (.A(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__and3_1 _1830_ (.A(\ByteBuffer.instr[21] ),
    .B(_0670_),
    .C(_1044_),
    .X(_1173_));
 sky130_fd_sc_hd__nand2_1 _1831_ (.A(_1151_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_2 _1832_ (.A(_1043_),
    .B(_1173_),
    .Y(_1175_));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(_1174_),
    .A1(_1175_),
    .S(_0947_),
    .X(_1176_));
 sky130_fd_sc_hd__o21ai_1 _1834_ (.A1(_1172_),
    .A2(_1067_),
    .B1(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__a31o_1 _1835_ (.A1(_0908_),
    .A2(_1043_),
    .A3(_1165_),
    .B1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__a211o_1 _1836_ (.A1(_0960_),
    .A2(_1162_),
    .B1(_1170_),
    .C1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__a21o_1 _1837_ (.A1(_1158_),
    .A2(_1161_),
    .B1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__nand2_1 _1838_ (.A(_1130_),
    .B(_1166_),
    .Y(_1181_));
 sky130_fd_sc_hd__o31a_2 _1839_ (.A1(_1126_),
    .A2(_1152_),
    .A3(_1180_),
    .B1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__nand2_1 _1840_ (.A(_0655_),
    .B(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__a21bo_2 _1841_ (.A1(_0631_),
    .A2(_1094_),
    .B1_N(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__nor2_1 _1842_ (.A(_0642_),
    .B(_0666_),
    .Y(_1185_));
 sky130_fd_sc_hd__a21o_1 _1843_ (.A1(\ByteBuffer.instr[20] ),
    .A2(_0665_),
    .B1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__nand2_1 _1844_ (.A(_0700_),
    .B(_0641_),
    .Y(_1187_));
 sky130_fd_sc_hd__a221o_2 _1845_ (.A1(_0700_),
    .A2(_1186_),
    .B1(_1187_),
    .B2(\ByteBuffer.instr[19] ),
    .C1(_0645_),
    .X(_1188_));
 sky130_fd_sc_hd__nor2_1 _1846_ (.A(_0668_),
    .B(_0696_),
    .Y(_1189_));
 sky130_fd_sc_hd__a2bb2o_1 _1847_ (.A1_N(_1189_),
    .A2_N(_0666_),
    .B1(_0665_),
    .B2(\ByteBuffer.instr[21] ),
    .X(_1190_));
 sky130_fd_sc_hd__a221o_2 _1848_ (.A1(\ByteBuffer.instr[20] ),
    .A2(_1187_),
    .B1(_1190_),
    .B2(_0700_),
    .C1(_0645_),
    .X(_1191_));
 sky130_fd_sc_hd__nand2_4 _1849_ (.A(_1188_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__a221o_2 _1850_ (.A1(_0700_),
    .A2(_1185_),
    .B1(_1187_),
    .B2(\ByteBuffer.instr[21] ),
    .C1(_0645_),
    .X(_1193_));
 sky130_fd_sc_hd__a211o_1 _1851_ (.A1(_0622_),
    .A2(\ByteBuffer.instr[19] ),
    .B1(_0624_),
    .C1(_0619_),
    .X(_1194_));
 sky130_fd_sc_hd__or3b_1 _1852_ (.A(_0647_),
    .B(_0656_),
    .C_N(_0660_),
    .X(_1195_));
 sky130_fd_sc_hd__a21oi_1 _1853_ (.A1(_1194_),
    .A2(_1195_),
    .B1(_0626_),
    .Y(_1196_));
 sky130_fd_sc_hd__a21o_1 _1854_ (.A1(_0645_),
    .A2(_0700_),
    .B1(_0661_),
    .X(_1197_));
 sky130_fd_sc_hd__nand2_1 _1855_ (.A(\ByteBuffer.instr[19] ),
    .B(_0660_),
    .Y(_1198_));
 sky130_fd_sc_hd__a31o_1 _1856_ (.A1(_0632_),
    .A2(_1197_),
    .A3(_1198_),
    .B1(_0663_),
    .X(_1199_));
 sky130_fd_sc_hd__or3b_1 _1857_ (.A(_1196_),
    .B(_0627_),
    .C_N(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_4 _1858_ (.A(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__o21bai_4 _1859_ (.A1(_0630_),
    .A2(_1193_),
    .B1_N(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__nor2_4 _1860_ (.A(_1192_),
    .B(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__mux2_1 _1861_ (.A0(\RegFile.A[7] ),
    .A1(_1184_),
    .S(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _1862_ (.A(_1204_),
    .X(_0157_));
 sky130_fd_sc_hd__o21ai_1 _1863_ (.A1(_1103_),
    .A2(_1119_),
    .B1(_1124_),
    .Y(_1205_));
 sky130_fd_sc_hd__a2bb2o_1 _1864_ (.A1_N(_1120_),
    .A2_N(_1205_),
    .B1(_1131_),
    .B2(_1166_),
    .X(_1206_));
 sky130_fd_sc_hd__nor2_2 _1865_ (.A(_1151_),
    .B(_1123_),
    .Y(_1207_));
 sky130_fd_sc_hd__or2_1 _1866_ (.A(_1131_),
    .B(_1147_),
    .X(_1208_));
 sky130_fd_sc_hd__and3_1 _1867_ (.A(_1148_),
    .B(_1207_),
    .C(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__nand2_2 _1868_ (.A(_1043_),
    .B(_1160_),
    .Y(_1210_));
 sky130_fd_sc_hd__and2_1 _1869_ (.A(_0983_),
    .B(_1155_),
    .X(_1211_));
 sky130_fd_sc_hd__or2_1 _1870_ (.A(_1156_),
    .B(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__o21ai_4 _1871_ (.A1(_1092_),
    .A2(_1160_),
    .B1(_1151_),
    .Y(_1213_));
 sky130_fd_sc_hd__or2_2 _1872_ (.A(_1122_),
    .B(_1163_),
    .X(_1214_));
 sky130_fd_sc_hd__nand2_1 _1873_ (.A(_1066_),
    .B(_1165_),
    .Y(_1215_));
 sky130_fd_sc_hd__o221a_1 _1874_ (.A1(_0781_),
    .A2(_1214_),
    .B1(_1076_),
    .B2(_1168_),
    .C1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_1 _1875_ (.A0(_1175_),
    .A1(_1174_),
    .S(_1069_),
    .X(_1217_));
 sky130_fd_sc_hd__o211a_1 _1876_ (.A1(_1070_),
    .A2(_1172_),
    .B1(_1216_),
    .C1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__o221a_1 _1877_ (.A1(_1100_),
    .A2(_1210_),
    .B1(_1212_),
    .B2(_1213_),
    .C1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__or3b_1 _1878_ (.A(_1206_),
    .B(_1209_),
    .C_N(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__buf_2 _1879_ (.A(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _1880_ (.A0(_1025_),
    .A1(_1088_),
    .S(net48),
    .X(_1222_));
 sky130_fd_sc_hd__xor2_1 _1881_ (.A(_0718_),
    .B(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__and2_1 _1882_ (.A(_1092_),
    .B(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__a22o_1 _1883_ (.A1(_0655_),
    .A2(_1221_),
    .B1(_1224_),
    .B2(_0631_),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(\RegFile.A[6] ),
    .A1(_1225_),
    .S(_1203_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _1885_ (.A(_1226_),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _1886_ (.A(_1136_),
    .B(_1146_),
    .X(_1227_));
 sky130_fd_sc_hd__a21bo_1 _1887_ (.A1(_1134_),
    .A2(_1227_),
    .B1_N(_1207_),
    .X(_1228_));
 sky130_fd_sc_hd__xnor2_1 _1888_ (.A(_1132_),
    .B(_1154_),
    .Y(_1229_));
 sky130_fd_sc_hd__nand2_1 _1889_ (.A(_1069_),
    .B(_1165_),
    .Y(_1230_));
 sky130_fd_sc_hd__o221a_1 _1890_ (.A1(_1071_),
    .A2(_1172_),
    .B1(_1214_),
    .B2(_0922_),
    .C1(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__mux2_1 _1891_ (.A0(_1174_),
    .A1(_1175_),
    .S(_0781_),
    .X(_1232_));
 sky130_fd_sc_hd__o211a_1 _1892_ (.A1(_1073_),
    .A2(_1168_),
    .B1(_1231_),
    .C1(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__o221a_1 _1893_ (.A1(_0806_),
    .A2(_1210_),
    .B1(_1229_),
    .B2(_1213_),
    .C1(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__or2_1 _1894_ (.A(_1151_),
    .B(_1134_),
    .X(_1235_));
 sky130_fd_sc_hd__or2_1 _1895_ (.A(_1043_),
    .B(_1123_),
    .X(_1236_));
 sky130_fd_sc_hd__a31o_1 _1896_ (.A1(_1117_),
    .A2(_1105_),
    .A3(_1116_),
    .B1(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__o22a_1 _1897_ (.A1(_1049_),
    .A2(_1235_),
    .B1(_1237_),
    .B2(_1118_),
    .X(_1238_));
 sky130_fd_sc_hd__o211ai_4 _1898_ (.A1(_1147_),
    .A2(_1228_),
    .B1(_1234_),
    .C1(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__inv_2 _1899_ (.A(_1086_),
    .Y(_1240_));
 sky130_fd_sc_hd__a211o_1 _1900_ (.A1(_1022_),
    .A2(_1085_),
    .B1(_1240_),
    .C1(_1151_),
    .X(_1241_));
 sky130_fd_sc_hd__nand2_1 _1901_ (.A(_1151_),
    .B(_1021_),
    .Y(_1242_));
 sky130_fd_sc_hd__a21o_1 _1902_ (.A1(_1000_),
    .A2(_1020_),
    .B1(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__a21oi_1 _1903_ (.A1(_1241_),
    .A2(_1243_),
    .B1(_1011_),
    .Y(_1244_));
 sky130_fd_sc_hd__a31o_1 _1904_ (.A1(_1011_),
    .A2(_1241_),
    .A3(_1243_),
    .B1(_1049_),
    .X(_1245_));
 sky130_fd_sc_hd__nor2_2 _1905_ (.A(_1244_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a22o_1 _1906_ (.A1(_0655_),
    .A2(_1239_),
    .B1(_1246_),
    .B2(_0631_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _1907_ (.A0(\RegFile.A[5] ),
    .A1(_1247_),
    .S(_1203_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _1908_ (.A(_1248_),
    .X(_0155_));
 sky130_fd_sc_hd__a21boi_1 _1909_ (.A1(_1136_),
    .A2(_1146_),
    .B1_N(_1207_),
    .Y(_1249_));
 sky130_fd_sc_hd__o31a_1 _1910_ (.A1(_0832_),
    .A2(_0856_),
    .A3(_0912_),
    .B1(_0913_),
    .X(_1250_));
 sky130_fd_sc_hd__nor2_1 _1911_ (.A(_0937_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__or2_1 _1912_ (.A(_0938_),
    .B(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__inv_2 _1913_ (.A(_1165_),
    .Y(_1253_));
 sky130_fd_sc_hd__and2_1 _1914_ (.A(_1151_),
    .B(_1173_),
    .X(_1254_));
 sky130_fd_sc_hd__and3_1 _1915_ (.A(_1151_),
    .B(_1048_),
    .C(_1159_),
    .X(_1255_));
 sky130_fd_sc_hd__nor2_1 _1916_ (.A(_1254_),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__and2_1 _1917_ (.A(_0780_),
    .B(_0921_),
    .X(_1257_));
 sky130_fd_sc_hd__or2_1 _1918_ (.A(_1257_),
    .B(_1175_),
    .X(_1258_));
 sky130_fd_sc_hd__o221a_1 _1919_ (.A1(_0781_),
    .A2(_1253_),
    .B1(_1256_),
    .B2(_0922_),
    .C1(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a22o_1 _1920_ (.A1(_0934_),
    .A2(_1255_),
    .B1(_1164_),
    .B2(_0855_),
    .X(_1260_));
 sky130_fd_sc_hd__o21ba_1 _1921_ (.A1(_1072_),
    .A2(_1172_),
    .B1_N(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__o211a_1 _1922_ (.A1(_0937_),
    .A2(_1210_),
    .B1(_1259_),
    .C1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__o221ai_2 _1923_ (.A1(_1093_),
    .A2(_1136_),
    .B1(_1213_),
    .B2(_1252_),
    .C1(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__o211a_1 _1924_ (.A1(_0937_),
    .A2(_1114_),
    .B1(_1116_),
    .C1(_1124_),
    .X(_1264_));
 sky130_fd_sc_hd__a211o_4 _1925_ (.A1(_1227_),
    .A2(_1249_),
    .B1(_1263_),
    .C1(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _1926_ (.A0(_1000_),
    .A1(_1085_),
    .S(net48),
    .X(_1266_));
 sky130_fd_sc_hd__nand2_1 _1927_ (.A(_1022_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__o211a_1 _1928_ (.A1(_1022_),
    .A2(_1266_),
    .B1(_1267_),
    .C1(_1092_),
    .X(_1268_));
 sky130_fd_sc_hd__a22o_1 _1929_ (.A1(_0655_),
    .A2(_1265_),
    .B1(_1268_),
    .B2(_0631_),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _1930_ (.A0(\RegFile.A[4] ),
    .A1(_1269_),
    .S(_1203_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _1931_ (.A(_1270_),
    .X(_0154_));
 sky130_fd_sc_hd__nand2_1 _1932_ (.A(_1106_),
    .B(_1112_),
    .Y(_1271_));
 sky130_fd_sc_hd__or2_1 _1933_ (.A(_1113_),
    .B(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__a21oi_1 _1934_ (.A1(_1114_),
    .A2(_1272_),
    .B1(_1236_),
    .Y(_1273_));
 sky130_fd_sc_hd__o21a_1 _1935_ (.A1(_1143_),
    .A2(_1145_),
    .B1(_1207_),
    .X(_1274_));
 sky130_fd_sc_hd__nor2_1 _1936_ (.A(_0832_),
    .B(_0912_),
    .Y(_0174_));
 sky130_fd_sc_hd__xnor2_2 _1937_ (.A(_1113_),
    .B(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__o22a_1 _1938_ (.A1(_0855_),
    .A2(_1175_),
    .B1(_1214_),
    .B2(_0816_),
    .X(_0176_));
 sky130_fd_sc_hd__o211a_1 _1939_ (.A1(_0922_),
    .A2(_1253_),
    .B1(_0176_),
    .C1(_1093_),
    .X(_0177_));
 sky130_fd_sc_hd__o221a_1 _1940_ (.A1(_1061_),
    .A2(_1172_),
    .B1(_1256_),
    .B2(_1056_),
    .C1(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__o21ai_1 _1941_ (.A1(_1113_),
    .A2(_1210_),
    .B1(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__a221o_1 _1942_ (.A1(_1146_),
    .A2(_1274_),
    .B1(_0175_),
    .B2(_1161_),
    .C1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__nor2_1 _1943_ (.A(_1093_),
    .B(_1145_),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _1944_ (.A(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__o21a_2 _1945_ (.A1(_1273_),
    .A2(_0180_),
    .B1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__a21boi_1 _1946_ (.A1(_0736_),
    .A2(_1082_),
    .B1_N(_0734_),
    .Y(_0184_));
 sky130_fd_sc_hd__mux2_1 _1947_ (.A0(_0997_),
    .A1(_0184_),
    .S(net48),
    .X(_0185_));
 sky130_fd_sc_hd__nand2_1 _1948_ (.A(_0726_),
    .B(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__o211a_2 _1949_ (.A1(_0726_),
    .A2(_0185_),
    .B1(_0186_),
    .C1(_1092_),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_1 _1950_ (.A1(_0655_),
    .A2(_0183_),
    .B1(_0187_),
    .B2(_0631_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _1951_ (.A0(\RegFile.A[3] ),
    .A1(_0188_),
    .S(_1203_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _1952_ (.A(_0189_),
    .X(_0153_));
 sky130_fd_sc_hd__a21bo_1 _1953_ (.A1(_1137_),
    .A2(_1142_),
    .B1_N(_1207_),
    .X(_0190_));
 sky130_fd_sc_hd__nor2_1 _1954_ (.A(_1143_),
    .B(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__a21oi_1 _1955_ (.A1(_1107_),
    .A2(_1111_),
    .B1(_1057_),
    .Y(_0192_));
 sky130_fd_sc_hd__a31o_1 _1956_ (.A1(_1057_),
    .A2(_1107_),
    .A3(_1111_),
    .B1(_1236_),
    .X(_0193_));
 sky130_fd_sc_hd__and3_1 _1957_ (.A(_0911_),
    .B(_0882_),
    .C(_0910_),
    .X(_0194_));
 sky130_fd_sc_hd__or2_1 _1958_ (.A(_0912_),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__nor2_1 _1959_ (.A(_1062_),
    .B(_1172_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _1960_ (.A(_0675_),
    .B(_0867_),
    .Y(_0197_));
 sky130_fd_sc_hd__a221o_1 _1961_ (.A1(_0855_),
    .A2(_1165_),
    .B1(_1164_),
    .B2(_0197_),
    .C1(_1166_),
    .X(_0198_));
 sky130_fd_sc_hd__a21oi_1 _1962_ (.A1(_1210_),
    .A2(_1168_),
    .B1(_1057_),
    .Y(_0199_));
 sky130_fd_sc_hd__mux2_1 _1963_ (.A0(_1256_),
    .A1(_1175_),
    .S(_0816_),
    .X(_0200_));
 sky130_fd_sc_hd__or4b_1 _1964_ (.A(_0196_),
    .B(_0198_),
    .C(_0199_),
    .D_N(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__o21ba_1 _1965_ (.A1(_1213_),
    .A2(_0195_),
    .B1_N(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__o21ai_1 _1966_ (.A1(_0192_),
    .A2(_0193_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__o2bb2a_4 _1967_ (.A1_N(_1166_),
    .A2_N(_1137_),
    .B1(_0191_),
    .B2(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _1968_ (.A(_0746_),
    .B(_0994_),
    .Y(_0205_));
 sky130_fd_sc_hd__mux2_1 _1969_ (.A0(_0205_),
    .A1(_1082_),
    .S(net48),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _1970_ (.A(_0736_),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__a211o_2 _1971_ (.A1(_0736_),
    .A2(_0206_),
    .B1(_0207_),
    .C1(_1049_),
    .X(_0208_));
 sky130_fd_sc_hd__inv_2 _1972_ (.A(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__a22o_1 _1973_ (.A1(_0655_),
    .A2(_0204_),
    .B1(_0209_),
    .B2(_0631_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _1974_ (.A0(\RegFile.A[2] ),
    .A1(_0210_),
    .S(_1203_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _1975_ (.A(_0211_),
    .X(_0152_));
 sky130_fd_sc_hd__xnor2_1 _1976_ (.A(_1139_),
    .B(_1059_),
    .Y(_0212_));
 sky130_fd_sc_hd__or2_1 _1977_ (.A(_1141_),
    .B(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__nand2_1 _1978_ (.A(_1108_),
    .B(_1110_),
    .Y(_0214_));
 sky130_fd_sc_hd__xor2_1 _1979_ (.A(_1139_),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__o22a_1 _1980_ (.A1(_0883_),
    .A2(_1172_),
    .B1(_1168_),
    .B2(_1058_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_1 _1981_ (.A(_1139_),
    .B(_0909_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _1982_ (.A(_0910_),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__a2bb2o_1 _1983_ (.A1_N(_0197_),
    .A2_N(_1175_),
    .B1(_1162_),
    .B2(_1139_),
    .X(_0219_));
 sky130_fd_sc_hd__a221o_1 _1984_ (.A1(_0197_),
    .A2(_1254_),
    .B1(_1164_),
    .B2(_0908_),
    .C1(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__o21ba_1 _1985_ (.A1(_1213_),
    .A2(_0218_),
    .B1_N(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__o211ai_1 _1986_ (.A1(_0816_),
    .A2(_1253_),
    .B1(_0216_),
    .C1(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__a221o_1 _1987_ (.A1(_1166_),
    .A2(_0212_),
    .B1(_0215_),
    .B2(_1124_),
    .C1(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__a31o_4 _1988_ (.A1(_1142_),
    .A2(_1207_),
    .A3(_0213_),
    .B1(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__a21oi_1 _1989_ (.A1(_0756_),
    .A2(_0990_),
    .B1(_0993_),
    .Y(_0225_));
 sky130_fd_sc_hd__mux2_1 _1990_ (.A0(_0225_),
    .A1(_1080_),
    .S(net48),
    .X(_0226_));
 sky130_fd_sc_hd__a21oi_1 _1991_ (.A1(_1054_),
    .A2(_0226_),
    .B1(_1049_),
    .Y(_0227_));
 sky130_fd_sc_hd__o21ai_2 _1992_ (.A1(_1054_),
    .A2(_0226_),
    .B1(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _1993_ (.A(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__a22o_1 _1994_ (.A1(_0655_),
    .A2(_0224_),
    .B1(_0229_),
    .B2(_0631_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _1995_ (.A0(\RegFile.A[1] ),
    .A1(_0230_),
    .S(_1203_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _1996_ (.A(_0231_),
    .X(_0151_));
 sky130_fd_sc_hd__and2_1 _1997_ (.A(_1059_),
    .B(_1140_),
    .X(_0232_));
 sky130_fd_sc_hd__a21oi_1 _1998_ (.A1(_0885_),
    .A2(_0896_),
    .B1(_1172_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor2_1 _1999_ (.A(_1109_),
    .B(_1123_),
    .Y(_0234_));
 sky130_fd_sc_hd__a21oi_1 _2000_ (.A1(_1059_),
    .A2(_1123_),
    .B1(_1141_),
    .Y(_0235_));
 sky130_fd_sc_hd__o32a_1 _2001_ (.A1(_0232_),
    .A2(_0233_),
    .A3(_0234_),
    .B1(_1162_),
    .B2(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__a32o_1 _2002_ (.A1(\ALU.flags_to_alu[0] ),
    .A2(_1151_),
    .A3(_1164_),
    .B1(_1254_),
    .B2(_0908_),
    .X(_0237_));
 sky130_fd_sc_hd__a2bb2o_1 _2003_ (.A1_N(_0908_),
    .A2_N(_1175_),
    .B1(_1165_),
    .B2(_0197_),
    .X(_0238_));
 sky130_fd_sc_hd__a21o_1 _2004_ (.A1(_1059_),
    .A2(_1161_),
    .B1(_1255_),
    .X(_0239_));
 sky130_fd_sc_hd__nor2_1 _2005_ (.A(_0947_),
    .B(_1214_),
    .Y(_0240_));
 sky130_fd_sc_hd__a22o_1 _2006_ (.A1(_1140_),
    .A2(_0239_),
    .B1(_0240_),
    .B2(_1043_),
    .X(_0241_));
 sky130_fd_sc_hd__or3_1 _2007_ (.A(_0237_),
    .B(_0238_),
    .C(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__a211o_2 _2008_ (.A1(_1166_),
    .A2(_0232_),
    .B1(_0236_),
    .C1(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_1 _2009_ (.A(net48),
    .B(_1079_),
    .Y(_0244_));
 sky130_fd_sc_hd__or2_1 _2010_ (.A(net48),
    .B(_0990_),
    .X(_0245_));
 sky130_fd_sc_hd__a21oi_1 _2011_ (.A1(_0244_),
    .A2(_0245_),
    .B1(_0756_),
    .Y(_0246_));
 sky130_fd_sc_hd__a31o_1 _2012_ (.A1(_0756_),
    .A2(_0244_),
    .A3(_0245_),
    .B1(_1049_),
    .X(_0247_));
 sky130_fd_sc_hd__nor2_2 _2013_ (.A(_0246_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__a22o_1 _2014_ (.A1(_0655_),
    .A2(_0243_),
    .B1(_0248_),
    .B2(_0631_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(\RegFile.A[0] ),
    .A1(_0249_),
    .S(_1203_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _2016_ (.A(_0250_),
    .X(_0150_));
 sky130_fd_sc_hd__or4_1 _2017_ (.A(_1188_),
    .B(_1191_),
    .C(_1201_),
    .D(_1193_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_4 _2018_ (.A(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _2019_ (.A0(_1184_),
    .A1(\RegFile.B[7] ),
    .S(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_1 _2020_ (.A(_0253_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2021_ (.A0(_1225_),
    .A1(\RegFile.B[6] ),
    .S(_0252_),
    .X(_0254_));
 sky130_fd_sc_hd__clkbuf_1 _2022_ (.A(_0254_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(_1247_),
    .A1(\RegFile.B[5] ),
    .S(_0252_),
    .X(_0255_));
 sky130_fd_sc_hd__clkbuf_1 _2024_ (.A(_0255_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2025_ (.A0(_1269_),
    .A1(\RegFile.B[4] ),
    .S(_0252_),
    .X(_0256_));
 sky130_fd_sc_hd__clkbuf_1 _2026_ (.A(_0256_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2027_ (.A0(_0188_),
    .A1(\RegFile.B[3] ),
    .S(_0252_),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_1 _2028_ (.A(_0257_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2029_ (.A0(_0210_),
    .A1(\RegFile.B[2] ),
    .S(_0252_),
    .X(_0258_));
 sky130_fd_sc_hd__clkbuf_1 _2030_ (.A(_0258_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2031_ (.A0(_0230_),
    .A1(\RegFile.B[1] ),
    .S(_0252_),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _2032_ (.A(_0259_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2033_ (.A0(_0249_),
    .A1(\RegFile.B[0] ),
    .S(_0252_),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_1 _2034_ (.A(_0260_),
    .X(_0142_));
 sky130_fd_sc_hd__nor2_2 _2035_ (.A(_0621_),
    .B(_0628_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_4 _2036_ (.A(\ByteBuffer.instr[19] ),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__and4_2 _2037_ (.A(\ByteBuffer.instr[19] ),
    .B(net1),
    .C(net4),
    .D(_0261_),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_2 _2038_ (.A1(_1182_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net10),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_1 _2039_ (.A(_1188_),
    .B(_1191_),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_2 _2040_ (.A(_1188_),
    .Y(_0266_));
 sky130_fd_sc_hd__nor2_1 _2041_ (.A(_0266_),
    .B(_1191_),
    .Y(_0267_));
 sky130_fd_sc_hd__or2_2 _2042_ (.A(_0630_),
    .B(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__a21oi_2 _2043_ (.A1(_0655_),
    .A2(_1193_),
    .B1(_1201_),
    .Y(_0269_));
 sky130_fd_sc_hd__o211a_4 _2044_ (.A1(_0655_),
    .A2(_0265_),
    .B1(_0268_),
    .C1(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2045_ (.A0(\RegFile.C[7] ),
    .A1(_0264_),
    .S(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _2046_ (.A(_0271_),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_1 _2047_ (.A1(_1221_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net9),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _2048_ (.A0(\RegFile.C[6] ),
    .A1(_0272_),
    .S(_0270_),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _2049_ (.A(_0273_),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _2050_ (.A1(_1239_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net8),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2051_ (.A0(\RegFile.C[5] ),
    .A1(_0274_),
    .S(_0270_),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _2052_ (.A(_0275_),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_1 _2053_ (.A1(_1265_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net7),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2054_ (.A0(\RegFile.C[4] ),
    .A1(_0276_),
    .S(_0270_),
    .X(_0277_));
 sky130_fd_sc_hd__clkbuf_1 _2055_ (.A(_0277_),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_1 _2056_ (.A1(_0183_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net6),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2057_ (.A0(\RegFile.C[3] ),
    .A1(_0278_),
    .S(_0270_),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_1 _2058_ (.A(_0279_),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _2059_ (.A1(_0204_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net5),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2060_ (.A0(\RegFile.C[2] ),
    .A1(_0280_),
    .S(_0270_),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _2061_ (.A(_0281_),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _2062_ (.A1(_0224_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net3),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2063_ (.A0(\RegFile.C[1] ),
    .A1(_0282_),
    .S(_0270_),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_1 _2064_ (.A(_0283_),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _2065_ (.A1(_0243_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(net2),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(\RegFile.C[0] ),
    .A1(_0284_),
    .S(_0270_),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_1 _2067_ (.A(_0285_),
    .X(_0134_));
 sky130_fd_sc_hd__nand2_1 _2068_ (.A(_0266_),
    .B(_1191_),
    .Y(_0286_));
 sky130_fd_sc_hd__and2_2 _2069_ (.A(_0655_),
    .B(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__o21ai_4 _2070_ (.A1(_0655_),
    .A2(_0267_),
    .B1(_0269_),
    .Y(_0288_));
 sky130_fd_sc_hd__nor2_4 _2071_ (.A(_0287_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(\RegFile.D[7] ),
    .A1(_1184_),
    .S(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _2073_ (.A(_0290_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _2074_ (.A0(\RegFile.D[6] ),
    .A1(_1225_),
    .S(_0289_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _2075_ (.A(_0291_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2076_ (.A0(\RegFile.D[5] ),
    .A1(_1247_),
    .S(_0289_),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _2077_ (.A(_0292_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2078_ (.A0(\RegFile.D[4] ),
    .A1(_1269_),
    .S(_0289_),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _2079_ (.A(_0293_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2080_ (.A0(\RegFile.D[3] ),
    .A1(_0188_),
    .S(_0289_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _2081_ (.A(_0294_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2082_ (.A0(\RegFile.D[2] ),
    .A1(_0210_),
    .S(_0289_),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _2083_ (.A(_0295_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2084_ (.A0(\RegFile.D[1] ),
    .A1(_0230_),
    .S(_0289_),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _2085_ (.A(_0296_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _2086_ (.A0(\RegFile.D[0] ),
    .A1(_0249_),
    .S(_0289_),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _2087_ (.A(_0297_),
    .X(_0126_));
 sky130_fd_sc_hd__a21oi_4 _2088_ (.A1(_1192_),
    .A2(_0655_),
    .B1(_0288_),
    .Y(_0298_));
 sky130_fd_sc_hd__mux2_1 _2089_ (.A0(\RegFile.E[7] ),
    .A1(_0264_),
    .S(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _2090_ (.A(_0299_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2091_ (.A0(\RegFile.E[6] ),
    .A1(_0272_),
    .S(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _2092_ (.A(_0300_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2093_ (.A0(\RegFile.E[5] ),
    .A1(_0274_),
    .S(_0298_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _2094_ (.A(_0301_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2095_ (.A0(\RegFile.E[4] ),
    .A1(_0276_),
    .S(_0298_),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _2096_ (.A(_0302_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2097_ (.A0(\RegFile.E[3] ),
    .A1(_0278_),
    .S(_0298_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _2098_ (.A(_0303_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2099_ (.A0(\RegFile.E[2] ),
    .A1(_0280_),
    .S(_0298_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _2100_ (.A(_0304_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2101_ (.A0(\RegFile.E[1] ),
    .A1(_0282_),
    .S(_0298_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _2102_ (.A(_0305_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2103_ (.A0(\RegFile.E[0] ),
    .A1(_0284_),
    .S(_0298_),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _2104_ (.A(_0306_),
    .X(_0118_));
 sky130_fd_sc_hd__a21oi_2 _2105_ (.A1(_0630_),
    .A2(_0286_),
    .B1(_1202_),
    .Y(_0307_));
 sky130_fd_sc_hd__o21ai_4 _2106_ (.A1(_0630_),
    .A2(_0265_),
    .B1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(_1184_),
    .A1(\RegFile.H[7] ),
    .S(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _2108_ (.A(_0309_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(_1225_),
    .A1(\RegFile.H[6] ),
    .S(_0308_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _2110_ (.A(_0310_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2111_ (.A0(_1247_),
    .A1(\RegFile.H[5] ),
    .S(_0308_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_1 _2112_ (.A(_0311_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2113_ (.A0(_1269_),
    .A1(\RegFile.H[4] ),
    .S(_0308_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _2114_ (.A(_0312_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(_0188_),
    .A1(\RegFile.H[3] ),
    .S(_0308_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _2116_ (.A(_0313_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(_0210_),
    .A1(\RegFile.H[2] ),
    .S(_0308_),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _2118_ (.A(_0314_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2119_ (.A0(_0230_),
    .A1(\RegFile.H[1] ),
    .S(_0308_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _2120_ (.A(_0315_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _2121_ (.A0(_0249_),
    .A1(\RegFile.H[0] ),
    .S(_0308_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _2122_ (.A(_0316_),
    .X(_0110_));
 sky130_fd_sc_hd__nand2_4 _2123_ (.A(_0268_),
    .B(_0307_),
    .Y(_0317_));
 sky130_fd_sc_hd__mux2_1 _2124_ (.A0(_0264_),
    .A1(\RegFile.L[7] ),
    .S(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _2125_ (.A(_0318_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2126_ (.A0(_0272_),
    .A1(\RegFile.L[6] ),
    .S(_0317_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _2127_ (.A(_0319_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2128_ (.A0(_0274_),
    .A1(\RegFile.L[5] ),
    .S(_0317_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _2129_ (.A(_0320_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2130_ (.A0(_0276_),
    .A1(\RegFile.L[4] ),
    .S(_0317_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _2131_ (.A(_0321_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2132_ (.A0(_0278_),
    .A1(\RegFile.L[3] ),
    .S(_0317_),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _2133_ (.A(_0322_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2134_ (.A0(_0280_),
    .A1(\RegFile.L[2] ),
    .S(_0317_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _2135_ (.A(_0323_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2136_ (.A0(_0282_),
    .A1(\RegFile.L[1] ),
    .S(_0317_),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _2137_ (.A(_0324_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2138_ (.A0(_0284_),
    .A1(\RegFile.L[0] ),
    .S(_0317_),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _2139_ (.A(_0325_),
    .X(_0102_));
 sky130_fd_sc_hd__nand2_1 _2140_ (.A(_0630_),
    .B(_1094_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_1 _2141_ (.A(_1183_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__mux2_1 _2142_ (.A0(_0264_),
    .A1(_0327_),
    .S(_1201_),
    .X(_0328_));
 sky130_fd_sc_hd__a21oi_1 _2143_ (.A1(_0619_),
    .A2(_0668_),
    .B1(_0620_),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_1 _2144_ (.A(_0619_),
    .B(_0620_),
    .Y(_0330_));
 sky130_fd_sc_hd__a21o_1 _2145_ (.A1(_0330_),
    .A2(_0696_),
    .B1(_0618_),
    .X(_0331_));
 sky130_fd_sc_hd__o21a_1 _2146_ (.A1(_0647_),
    .A2(_0329_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__a2bb2o_1 _2147_ (.A1_N(_0332_),
    .A2_N(_0626_),
    .B1(_0645_),
    .B2(_1197_),
    .X(_0333_));
 sky130_fd_sc_hd__a211oi_4 _2148_ (.A1(_1192_),
    .A2(_0630_),
    .B1(_1202_),
    .C1(_0287_),
    .Y(_0334_));
 sky130_fd_sc_hd__a31o_2 _2149_ (.A1(_0659_),
    .A2(_1201_),
    .A3(_0333_),
    .B1(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _2150_ (.A0(\ALU.flags_to_alu[7] ),
    .A1(_0328_),
    .S(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_1 _2151_ (.A(_0336_),
    .X(_0101_));
 sky130_fd_sc_hd__inv_2 _2152_ (.A(_0335_),
    .Y(_0337_));
 sky130_fd_sc_hd__or4_1 _2153_ (.A(_1224_),
    .B(_1246_),
    .C(_1268_),
    .D(_0209_),
    .X(_0338_));
 sky130_fd_sc_hd__o31a_1 _2154_ (.A1(_1094_),
    .A2(_0187_),
    .A3(_0338_),
    .B1(_0630_),
    .X(_0339_));
 sky130_fd_sc_hd__o21a_1 _2155_ (.A1(_0229_),
    .A2(_0248_),
    .B1(_0630_),
    .X(_0340_));
 sky130_fd_sc_hd__or4_1 _2156_ (.A(_0183_),
    .B(_0204_),
    .C(_0224_),
    .D(_0243_),
    .X(_0341_));
 sky130_fd_sc_hd__or4_1 _2157_ (.A(_1221_),
    .B(_1239_),
    .C(_1265_),
    .D(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__or4_2 _2158_ (.A(_1182_),
    .B(_0339_),
    .C(_0340_),
    .D(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__nand2_1 _2159_ (.A(_1201_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__o21a_1 _2160_ (.A1(_1201_),
    .A2(_0272_),
    .B1(_0335_),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_1 _2161_ (.A1(net137),
    .A2(_0337_),
    .B1(_0344_),
    .B2(_0345_),
    .X(_0100_));
 sky130_fd_sc_hd__a22o_1 _2162_ (.A1(_0274_),
    .A2(_0334_),
    .B1(_0337_),
    .B2(net138),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _2163_ (.A1(_0276_),
    .A2(_0334_),
    .B1(_0337_),
    .B2(net136),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_1 _2164_ (.A1(_0278_),
    .A2(_0334_),
    .B1(_0337_),
    .B2(net135),
    .X(_0097_));
 sky130_fd_sc_hd__xor2_1 _2165_ (.A(_1094_),
    .B(_0187_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_2 _2166_ (.A(_1151_),
    .B(_1092_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _2167_ (.A(_1257_),
    .B(_1049_),
    .Y(_0348_));
 sky130_fd_sc_hd__o221a_1 _2168_ (.A1(_1093_),
    .A2(_1136_),
    .B1(_0347_),
    .B2(_1252_),
    .C1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__a22o_1 _2169_ (.A1(_0816_),
    .A2(_1049_),
    .B1(_1166_),
    .B2(_1137_),
    .X(_0350_));
 sky130_fd_sc_hd__a21oi_1 _2170_ (.A1(_1050_),
    .A2(_0195_),
    .B1(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _2171_ (.A(_1050_),
    .B(_0218_),
    .Y(_0352_));
 sky130_fd_sc_hd__o221a_1 _2172_ (.A1(_0197_),
    .A2(_1092_),
    .B1(_1093_),
    .B2(_0212_),
    .C1(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__xnor2_1 _2173_ (.A(_0351_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__xnor2_1 _2174_ (.A(_0349_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__o211a_1 _2175_ (.A1(_1043_),
    .A2(_1229_),
    .B1(_1235_),
    .C1(_1092_),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_1 _2176_ (.A1(_0781_),
    .A2(_1049_),
    .B1(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__mux2_1 _2177_ (.A0(_0908_),
    .A1(_0232_),
    .S(_1092_),
    .X(_0358_));
 sky130_fd_sc_hd__xnor2_1 _2178_ (.A(_0357_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__xnor2_1 _2179_ (.A(_0355_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__xnor2_1 _2180_ (.A(_0346_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__xnor2_1 _2181_ (.A(_1246_),
    .B(_1268_),
    .Y(_0362_));
 sky130_fd_sc_hd__a21oi_1 _2182_ (.A1(_1092_),
    .A2(_1223_),
    .B1(_0228_),
    .Y(_0363_));
 sky130_fd_sc_hd__and3_1 _2183_ (.A(_1092_),
    .B(_1223_),
    .C(_0228_),
    .X(_0364_));
 sky130_fd_sc_hd__or3_1 _2184_ (.A(_0362_),
    .B(_0363_),
    .C(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__o21ai_1 _2185_ (.A1(_0363_),
    .A2(_0364_),
    .B1(_0362_),
    .Y(_0366_));
 sky130_fd_sc_hd__o221a_1 _2186_ (.A1(_1066_),
    .A2(_1092_),
    .B1(_1158_),
    .B2(_0347_),
    .C1(_1181_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _2187_ (.A(_1050_),
    .B(_1212_),
    .Y(_0368_));
 sky130_fd_sc_hd__o221a_1 _2188_ (.A1(_1069_),
    .A2(_1092_),
    .B1(_1093_),
    .B2(_1131_),
    .C1(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__xnor2_1 _2189_ (.A(_0248_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__xnor2_1 _2190_ (.A(_0367_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__xnor2_1 _2191_ (.A(_0208_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21oi_1 _2192_ (.A1(_0365_),
    .A2(_0366_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__and3_1 _2193_ (.A(_0365_),
    .B(_0366_),
    .C(_0372_),
    .X(_0374_));
 sky130_fd_sc_hd__or3_1 _2194_ (.A(_0361_),
    .B(_0373_),
    .C(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__o21ai_1 _2195_ (.A1(_0373_),
    .A2(_0374_),
    .B1(_0361_),
    .Y(_0376_));
 sky130_fd_sc_hd__o221ai_4 _2196_ (.A1(_0855_),
    .A2(_1092_),
    .B1(_0347_),
    .B2(_0175_),
    .C1(_0182_),
    .Y(_0377_));
 sky130_fd_sc_hd__a21oi_1 _2197_ (.A1(_0375_),
    .A2(_0376_),
    .B1(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__and3_1 _2198_ (.A(_0377_),
    .B(_0375_),
    .C(_0376_),
    .X(_0379_));
 sky130_fd_sc_hd__xor2_1 _2199_ (.A(_1221_),
    .B(_1265_),
    .X(_0380_));
 sky130_fd_sc_hd__xnor2_1 _2200_ (.A(_0243_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__xor2_1 _2201_ (.A(_1182_),
    .B(_0204_),
    .X(_0382_));
 sky130_fd_sc_hd__xnor2_1 _2202_ (.A(_0381_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__xnor2_1 _2203_ (.A(_1239_),
    .B(_0224_),
    .Y(_0384_));
 sky130_fd_sc_hd__xnor2_1 _2204_ (.A(_0383_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__xnor2_1 _2205_ (.A(_0183_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__nand2_1 _2206_ (.A(_0655_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__o31ai_4 _2207_ (.A1(_0655_),
    .A2(_0378_),
    .A3(_0379_),
    .B1(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(_0280_),
    .A1(_0388_),
    .S(_1201_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2209_ (.A0(\ALU.flags_to_alu[2] ),
    .A1(_0389_),
    .S(_0335_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _2210_ (.A(_0390_),
    .X(_0096_));
 sky130_fd_sc_hd__inv_2 _2211_ (.A(_0334_),
    .Y(_0391_));
 sky130_fd_sc_hd__o22a_1 _2212_ (.A1(_0282_),
    .A2(_0391_),
    .B1(_0335_),
    .B2(net132),
    .X(_0095_));
 sky130_fd_sc_hd__a21o_1 _2213_ (.A1(_1096_),
    .A2(_1125_),
    .B1(_0986_),
    .X(_0392_));
 sky130_fd_sc_hd__nand2_1 _2214_ (.A(_1124_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__o21ai_1 _2215_ (.A1(_1149_),
    .A2(_1079_),
    .B1(_1207_),
    .Y(_0394_));
 sky130_fd_sc_hd__o21ai_1 _2216_ (.A1(\ALU.flags_to_alu[0] ),
    .A2(_1151_),
    .B1(_1173_),
    .Y(_0395_));
 sky130_fd_sc_hd__a31o_1 _2217_ (.A1(\ALU.flags_to_alu[0] ),
    .A2(_1151_),
    .A3(_1122_),
    .B1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__a21oi_1 _2218_ (.A1(_0908_),
    .A2(_1165_),
    .B1(_0240_),
    .Y(_0397_));
 sky130_fd_sc_hd__o2111a_1 _2219_ (.A1(_1213_),
    .A2(_0990_),
    .B1(_0394_),
    .C1(_0396_),
    .D1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__o211a_1 _2220_ (.A1(_1049_),
    .A2(_0244_),
    .B1(_0398_),
    .C1(_0655_),
    .X(_0399_));
 sky130_fd_sc_hd__inv_2 _2221_ (.A(_1029_),
    .Y(_0400_));
 sky130_fd_sc_hd__nor2_1 _2222_ (.A(_0400_),
    .B(_1033_),
    .Y(_0401_));
 sky130_fd_sc_hd__a211o_1 _2223_ (.A1(_1034_),
    .A2(_1089_),
    .B1(_1035_),
    .C1(_1093_),
    .X(_0402_));
 sky130_fd_sc_hd__o311a_1 _2224_ (.A1(_0347_),
    .A2(_1038_),
    .A3(_0401_),
    .B1(_0402_),
    .C1(_0630_),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_2 _2225_ (.A1(_0393_),
    .A2(_0399_),
    .B1(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__mux2_1 _2226_ (.A0(_0284_),
    .A1(_0404_),
    .S(_1201_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _2227_ (.A0(\ALU.flags_to_alu[0] ),
    .A1(_0405_),
    .S(_0335_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _2228_ (.A(_0406_),
    .X(_0094_));
 sky130_fd_sc_hd__nor2_1 _2229_ (.A(net128),
    .B(_0659_),
    .Y(\ByteBuffer.next_counter[0] ));
 sky130_fd_sc_hd__nand2_4 _2230_ (.A(\ByteBuffer.counter[1] ),
    .B(\ByteBuffer.next_counter[0] ),
    .Y(_0407_));
 sky130_fd_sc_hd__or3b_1 _2231_ (.A(\ByteBuffer.counter[1] ),
    .B(_0659_),
    .C_N(\ByteBuffer.counter[0] ),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_4 _2232_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _2233_ (.A(_0407_),
    .B(_0409_),
    .Y(\ByteBuffer.next_counter[1] ));
 sky130_fd_sc_hd__and2_1 _2234_ (.A(\MemControl.state[0] ),
    .B(_0261_),
    .X(_0410_));
 sky130_fd_sc_hd__and3_2 _2235_ (.A(_0670_),
    .B(_0659_),
    .C(_0662_),
    .X(_0411_));
 sky130_fd_sc_hd__o21ba_2 _2236_ (.A1(\MemControl.state[2] ),
    .A2(\MemControl.state[1] ),
    .B1_N(\MemControl.state[0] ),
    .X(_0412_));
 sky130_fd_sc_hd__or3_2 _2237_ (.A(_0410_),
    .B(_0411_),
    .C(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__nor3_1 _2238_ (.A(\ByteDecoder.state[1] ),
    .B(\ByteDecoder.num_bytes[2] ),
    .C(\ByteDecoder.num_bytes[3] ),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_2 _2239_ (.A(\ByteDecoder.state[0] ),
    .Y(_0415_));
 sky130_fd_sc_hd__a221o_1 _2240_ (.A1(\ByteDecoder.state[1] ),
    .A2(_0413_),
    .B1(_0414_),
    .B2(net129),
    .C1(_0415_),
    .X(\FSM.next_state[0] ));
 sky130_fd_sc_hd__or2_1 _2241_ (.A(\ByteDecoder.state[1] ),
    .B(\ByteDecoder.state[0] ),
    .X(_0416_));
 sky130_fd_sc_hd__and2b_2 _2242_ (.A_N(net4),
    .B(net1),
    .X(_0417_));
 sky130_fd_sc_hd__and2_2 _2243_ (.A(net10),
    .B(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _2244_ (.A(net9),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__or2b_1 _2245_ (.A(net5),
    .B_N(net3),
    .X(_0420_));
 sky130_fd_sc_hd__and2_1 _2246_ (.A(net8),
    .B(_0417_),
    .X(_0421_));
 sky130_fd_sc_hd__and2_1 _2247_ (.A(net7),
    .B(_0417_),
    .X(_0422_));
 sky130_fd_sc_hd__or2b_1 _2248_ (.A(net3),
    .B_N(net5),
    .X(_0423_));
 sky130_fd_sc_hd__a21o_1 _2249_ (.A1(_0420_),
    .A2(_0423_),
    .B1(net2),
    .X(_0424_));
 sky130_fd_sc_hd__o31a_1 _2250_ (.A1(_0420_),
    .A2(_0421_),
    .A3(_0422_),
    .B1(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__and2_1 _2251_ (.A(net2),
    .B(_0417_),
    .X(_0426_));
 sky130_fd_sc_hd__or4b_1 _2252_ (.A(net3),
    .B(net5),
    .C(net6),
    .D_N(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__or3b_1 _2253_ (.A(net2),
    .B(_0420_),
    .C_N(_0421_),
    .X(_0428_));
 sky130_fd_sc_hd__and2_1 _2254_ (.A(net9),
    .B(_0417_),
    .X(_0429_));
 sky130_fd_sc_hd__a211o_1 _2255_ (.A1(_0427_),
    .A2(_0428_),
    .B1(_0418_),
    .C1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_1 _2256_ (.A(\ByteDecoder.state[1] ),
    .B(\ByteDecoder.state[0] ),
    .Y(_0431_));
 sky130_fd_sc_hd__o211ai_1 _2257_ (.A1(_0419_),
    .A2(_0425_),
    .B1(_0430_),
    .C1(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__and4bb_1 _2258_ (.A_N(net8),
    .B_N(_0420_),
    .C(_0426_),
    .D(net7),
    .X(_0433_));
 sky130_fd_sc_hd__o21ai_1 _2259_ (.A1(_0418_),
    .A2(_0429_),
    .B1(_0419_),
    .Y(_0434_));
 sky130_fd_sc_hd__and2_1 _2260_ (.A(net5),
    .B(_0417_),
    .X(_0435_));
 sky130_fd_sc_hd__and2_1 _2261_ (.A(net3),
    .B(_0417_),
    .X(_0436_));
 sky130_fd_sc_hd__and4b_1 _2262_ (.A_N(net2),
    .B(_0434_),
    .C(_0435_),
    .D(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__a31o_1 _2263_ (.A1(net9),
    .A2(_0418_),
    .A3(_0433_),
    .B1(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_1 _2264_ (.A(_0432_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a221o_1 _2265_ (.A1(net139),
    .A2(_0413_),
    .B1(_0416_),
    .B2(_0627_),
    .C1(_0439_),
    .X(\FSM.next_state[1] ));
 sky130_fd_sc_hd__or2_1 _2266_ (.A(\ByteBuffer.instr[19] ),
    .B(_0621_),
    .X(_0440_));
 sky130_fd_sc_hd__or2_1 _2267_ (.A(_0440_),
    .B(_0655_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_8 _2268_ (.A(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__inv_4 _2269_ (.A(_0442_),
    .Y(net46));
 sky130_fd_sc_hd__a21o_1 _2270_ (.A1(net131),
    .A2(_0411_),
    .B1(_0410_),
    .X(_0001_));
 sky130_fd_sc_hd__inv_2 _2271_ (.A(_0261_),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_2 _2272_ (.A(_0411_),
    .Y(_0444_));
 sky130_fd_sc_hd__a22o_1 _2273_ (.A1(\MemControl.state[0] ),
    .A2(_0443_),
    .B1(_0444_),
    .B2(net133),
    .X(_0000_));
 sky130_fd_sc_hd__buf_6 _2274_ (.A(net1),
    .X(_0445_));
 sky130_fd_sc_hd__and2_1 _2275_ (.A(\RegFile.A[0] ),
    .B(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _2276_ (.A(_0446_),
    .X(net30));
 sky130_fd_sc_hd__and2_1 _2277_ (.A(\RegFile.A[1] ),
    .B(_0445_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _2278_ (.A(_0447_),
    .X(net31));
 sky130_fd_sc_hd__and2_1 _2279_ (.A(\RegFile.A[2] ),
    .B(net1),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _2280_ (.A(_0448_),
    .X(net32));
 sky130_fd_sc_hd__and2_1 _2281_ (.A(\RegFile.A[3] ),
    .B(net1),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _2282_ (.A(_0449_),
    .X(net33));
 sky130_fd_sc_hd__and2_1 _2283_ (.A(\RegFile.A[4] ),
    .B(net1),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _2284_ (.A(_0450_),
    .X(net35));
 sky130_fd_sc_hd__and2_1 _2285_ (.A(\RegFile.A[5] ),
    .B(net1),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _2286_ (.A(_0451_),
    .X(net36));
 sky130_fd_sc_hd__and2_1 _2287_ (.A(\RegFile.A[6] ),
    .B(net1),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _2288_ (.A(_0452_),
    .X(net37));
 sky130_fd_sc_hd__and2_1 _2289_ (.A(\RegFile.A[7] ),
    .B(net1),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _2290_ (.A(_0453_),
    .X(net38));
 sky130_fd_sc_hd__a21boi_2 _2291_ (.A1(_0262_),
    .A2(_0413_),
    .B1_N(_0445_),
    .Y(net28));
 sky130_fd_sc_hd__and2_1 _2292_ (.A(_0445_),
    .B(net46),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _2293_ (.A(_0454_),
    .X(net29));
 sky130_fd_sc_hd__inv_2 _2294_ (.A(\PC.i_mem_addr[0] ),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _2295_ (.A(_0455_),
    .B(_0442_),
    .Y(_0456_));
 sky130_fd_sc_hd__o211a_1 _2296_ (.A1(_0243_),
    .A2(_0442_),
    .B1(_0456_),
    .C1(_0445_),
    .X(net44));
 sky130_fd_sc_hd__or2_1 _2297_ (.A(\PC.i_mem_addr[1] ),
    .B(net46),
    .X(_0457_));
 sky130_fd_sc_hd__o211a_1 _2298_ (.A1(_0224_),
    .A2(_0442_),
    .B1(_0457_),
    .C1(_0445_),
    .X(net45));
 sky130_fd_sc_hd__or2_1 _2299_ (.A(\PC.i_mem_addr[2] ),
    .B(net46),
    .X(_0458_));
 sky130_fd_sc_hd__o211a_1 _2300_ (.A1(_0204_),
    .A2(_0442_),
    .B1(_0458_),
    .C1(_0445_),
    .X(net13));
 sky130_fd_sc_hd__or2_1 _2301_ (.A(\PC.i_mem_addr[3] ),
    .B(net46),
    .X(_0459_));
 sky130_fd_sc_hd__o211a_1 _2302_ (.A1(_0183_),
    .A2(_0442_),
    .B1(_0459_),
    .C1(_0445_),
    .X(net14));
 sky130_fd_sc_hd__or2_1 _2303_ (.A(\PC.i_mem_addr[4] ),
    .B(net46),
    .X(_0460_));
 sky130_fd_sc_hd__o211a_1 _2304_ (.A1(_1265_),
    .A2(_0442_),
    .B1(_0460_),
    .C1(_0445_),
    .X(net15));
 sky130_fd_sc_hd__or2_1 _2305_ (.A(\PC.i_mem_addr[5] ),
    .B(net46),
    .X(_0461_));
 sky130_fd_sc_hd__o211a_1 _2306_ (.A1(_1239_),
    .A2(_0442_),
    .B1(_0461_),
    .C1(_0445_),
    .X(net16));
 sky130_fd_sc_hd__or2_1 _2307_ (.A(\PC.i_mem_addr[6] ),
    .B(net46),
    .X(_0462_));
 sky130_fd_sc_hd__o211a_1 _2308_ (.A1(_1221_),
    .A2(_0442_),
    .B1(_0462_),
    .C1(_0445_),
    .X(net17));
 sky130_fd_sc_hd__or2_1 _2309_ (.A(\PC.i_mem_addr[7] ),
    .B(net46),
    .X(_0463_));
 sky130_fd_sc_hd__o211a_1 _2310_ (.A1(_1182_),
    .A2(_0442_),
    .B1(_0463_),
    .C1(_0445_),
    .X(net18));
 sky130_fd_sc_hd__mux2_1 _2311_ (.A0(\PC.i_mem_addr[8] ),
    .A1(_0248_),
    .S(net46),
    .X(_0464_));
 sky130_fd_sc_hd__and2_1 _2312_ (.A(_0445_),
    .B(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _2313_ (.A(_0465_),
    .X(net19));
 sky130_fd_sc_hd__mux2_1 _2314_ (.A0(\PC.i_mem_addr[9] ),
    .A1(_0229_),
    .S(net46),
    .X(_0466_));
 sky130_fd_sc_hd__and2_1 _2315_ (.A(_0445_),
    .B(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__buf_1 _2316_ (.A(_0467_),
    .X(net20));
 sky130_fd_sc_hd__nand2_1 _2317_ (.A(_0208_),
    .B(net46),
    .Y(_0468_));
 sky130_fd_sc_hd__o211a_1 _2318_ (.A1(\PC.i_mem_addr[10] ),
    .A2(net46),
    .B1(_0468_),
    .C1(_0445_),
    .X(net21));
 sky130_fd_sc_hd__or2_1 _2319_ (.A(\PC.i_mem_addr[11] ),
    .B(net46),
    .X(_0469_));
 sky130_fd_sc_hd__o211a_1 _2320_ (.A1(_0187_),
    .A2(_0442_),
    .B1(_0469_),
    .C1(_0445_),
    .X(net22));
 sky130_fd_sc_hd__or2_1 _2321_ (.A(\PC.i_mem_addr[12] ),
    .B(net46),
    .X(_0470_));
 sky130_fd_sc_hd__o211a_1 _2322_ (.A1(_1268_),
    .A2(_0442_),
    .B1(_0470_),
    .C1(_0445_),
    .X(net24));
 sky130_fd_sc_hd__or2_1 _2323_ (.A(\PC.i_mem_addr[13] ),
    .B(net46),
    .X(_0471_));
 sky130_fd_sc_hd__o211a_1 _2324_ (.A1(_1246_),
    .A2(_0442_),
    .B1(_0471_),
    .C1(_0445_),
    .X(net25));
 sky130_fd_sc_hd__or2_1 _2325_ (.A(\PC.i_mem_addr[14] ),
    .B(net46),
    .X(_0472_));
 sky130_fd_sc_hd__o211a_1 _2326_ (.A1(_1224_),
    .A2(_0442_),
    .B1(_0472_),
    .C1(_0445_),
    .X(net26));
 sky130_fd_sc_hd__a2bb2o_1 _2327_ (.A1_N(_0440_),
    .A2_N(_0326_),
    .B1(_0442_),
    .B2(\PC.i_mem_addr[15] ),
    .X(_0473_));
 sky130_fd_sc_hd__and2_1 _2328_ (.A(_0445_),
    .B(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__buf_1 _2329_ (.A(_0474_),
    .X(net27));
 sky130_fd_sc_hd__nand3_1 _2330_ (.A(net1),
    .B(net4),
    .C(net46),
    .Y(_0475_));
 sky130_fd_sc_hd__inv_2 _2331_ (.A(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__and2_1 _2332_ (.A(_0752_),
    .B(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_1 _2333_ (.A(_0477_),
    .X(net12));
 sky130_fd_sc_hd__and2_1 _2334_ (.A(_0744_),
    .B(_0476_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _2335_ (.A(_0478_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _2336_ (.A(_0732_),
    .B(_0476_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _2337_ (.A(_0479_),
    .X(net34));
 sky130_fd_sc_hd__and2_1 _2338_ (.A(_0724_),
    .B(_0476_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _2339_ (.A(_0480_),
    .X(net39));
 sky130_fd_sc_hd__and2_1 _2340_ (.A(_1017_),
    .B(_0476_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _2341_ (.A(_0481_),
    .X(net40));
 sky130_fd_sc_hd__and2_1 _2342_ (.A(_1006_),
    .B(_0476_),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _2343_ (.A(_0482_),
    .X(net41));
 sky130_fd_sc_hd__and2_1 _2344_ (.A(_0713_),
    .B(_0476_),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_1 _2345_ (.A(_0483_),
    .X(net42));
 sky130_fd_sc_hd__and2_1 _2346_ (.A(_1032_),
    .B(_0476_),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _2347_ (.A(_0484_),
    .X(net43));
 sky130_fd_sc_hd__mux2_1 _2348_ (.A0(\MemControl.state[2] ),
    .A1(\MemControl.state[1] ),
    .S(_0411_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_1 _2349_ (.A(_0485_),
    .X(_0066_));
 sky130_fd_sc_hd__o21a_1 _2350_ (.A1(net127),
    .A2(_0431_),
    .B1(_0432_),
    .X(_0067_));
 sky130_fd_sc_hd__a21o_1 _2351_ (.A1(net126),
    .A2(_0416_),
    .B1(_0439_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2352_ (.A0(net129),
    .A1(_0438_),
    .S(_0431_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _2353_ (.A(_0486_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(_0426_),
    .A1(\ALU.immediate[8] ),
    .S(_0407_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _2355_ (.A(_0487_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2356_ (.A0(_0436_),
    .A1(\ALU.immediate[9] ),
    .S(_0407_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _2357_ (.A(_0488_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2358_ (.A0(_0435_),
    .A1(\ALU.immediate[10] ),
    .S(_0407_),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _2359_ (.A(_0489_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _2360_ (.A(net6),
    .B(_0417_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _2361_ (.A0(_0490_),
    .A1(\ALU.immediate[11] ),
    .S(_0407_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_1 _2362_ (.A(_0491_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2363_ (.A0(_0422_),
    .A1(\ALU.immediate[12] ),
    .S(_0407_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _2364_ (.A(_0492_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2365_ (.A0(_0421_),
    .A1(\ALU.immediate[13] ),
    .S(_0407_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _2366_ (.A(_0493_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(_0429_),
    .A1(\ALU.immediate[14] ),
    .S(_0407_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _2368_ (.A(_0494_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2369_ (.A0(_0418_),
    .A1(\ALU.immediate[15] ),
    .S(_0407_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _2370_ (.A(_0495_),
    .X(_0077_));
 sky130_fd_sc_hd__or3_1 _2371_ (.A(\ByteBuffer.counter[0] ),
    .B(\ByteBuffer.counter[1] ),
    .C(_0659_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_4 _2372_ (.A(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _2373_ (.A0(_0426_),
    .A1(_0619_),
    .S(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _2374_ (.A(_0498_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(_0436_),
    .A1(_0622_),
    .S(_0497_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _2376_ (.A(_0499_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2377_ (.A0(_0435_),
    .A1(_0624_),
    .S(_0497_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _2378_ (.A(_0500_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2379_ (.A0(_0490_),
    .A1(\ByteBuffer.instr[19] ),
    .S(_0497_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _2380_ (.A(_0501_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2381_ (.A0(_0422_),
    .A1(\ByteBuffer.instr[20] ),
    .S(_0497_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _2382_ (.A(_0502_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(_0421_),
    .A1(\ByteBuffer.instr[21] ),
    .S(_0497_),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _2384_ (.A(_0503_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2385_ (.A0(_0429_),
    .A1(\ByteBuffer.instr[22] ),
    .S(_0497_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _2386_ (.A(_0504_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(_0418_),
    .A1(_0645_),
    .S(_0497_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _2388_ (.A(_0505_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(_0426_),
    .A1(\ALU.immediate[0] ),
    .S(_0409_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_0506_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(_0436_),
    .A1(\ALU.immediate[1] ),
    .S(_0409_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _2392_ (.A(_0507_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(_0435_),
    .A1(\ALU.immediate[2] ),
    .S(_0409_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _2394_ (.A(_0508_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2395_ (.A0(_0490_),
    .A1(\ALU.immediate[3] ),
    .S(_0409_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _2396_ (.A(_0509_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(_0422_),
    .A1(\ALU.immediate[4] ),
    .S(_0409_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_1 _2398_ (.A(_0510_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(_0421_),
    .A1(\ALU.immediate[5] ),
    .S(_0409_),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_1 _2400_ (.A(_0511_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2401_ (.A0(_0429_),
    .A1(\ALU.immediate[6] ),
    .S(_0409_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _2402_ (.A(_0512_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(_0418_),
    .A1(\ALU.immediate[7] ),
    .S(_0409_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_1 _2404_ (.A(_0513_),
    .X(_0093_));
 sky130_fd_sc_hd__buf_1 _2405_ (.A(clknet_2_1__leaf_clk),
    .X(_0514_));
 sky130_fd_sc_hd__buf_1 _2406_ (.A(clknet_1_0__leaf__0514_),
    .X(_0515_));
 sky130_fd_sc_hd__inv_2 _2407__8 (.A(clknet_1_1__leaf__0515_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _2408__9 (.A(clknet_1_0__leaf__0515_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _2409__10 (.A(clknet_1_1__leaf__0515_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _2410__11 (.A(clknet_1_0__leaf__0515_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _2411__12 (.A(clknet_1_0__leaf__0515_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _2412__13 (.A(clknet_1_0__leaf__0515_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _2413__14 (.A(clknet_1_1__leaf__0515_),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _2414__15 (.A(clknet_1_0__leaf__0515_),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _2415__16 (.A(clknet_1_1__leaf__0515_),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _2416__17 (.A(clknet_1_0__leaf__0515_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _2417__18 (.A(clknet_1_1__leaf__0515_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _2418__19 (.A(clknet_1_0__leaf__0515_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _2419__20 (.A(clknet_1_0__leaf__0515_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _2420__21 (.A(clknet_1_0__leaf__0515_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _2421__22 (.A(clknet_1_0__leaf__0515_),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _2422__23 (.A(clknet_1_0__leaf__0515_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _2423__24 (.A(clknet_1_1__leaf__0515_),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _2424__25 (.A(clknet_1_0__leaf__0515_),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _2425__26 (.A(clknet_1_1__leaf__0515_),
    .Y(net87));
 sky130_fd_sc_hd__buf_1 _2426_ (.A(clknet_1_1__leaf__0514_),
    .X(_0516_));
 sky130_fd_sc_hd__inv_2 _2427__27 (.A(clknet_1_1__leaf__0516_),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _2428__28 (.A(clknet_1_1__leaf__0516_),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _2429__29 (.A(clknet_1_1__leaf__0516_),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _2430__30 (.A(clknet_1_1__leaf__0516_),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _2431__31 (.A(clknet_1_1__leaf__0516_),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _2432__32 (.A(clknet_1_0__leaf__0516_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _2433__33 (.A(clknet_1_0__leaf__0516_),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _2434__34 (.A(clknet_1_0__leaf__0516_),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _2435__35 (.A(clknet_1_0__leaf__0516_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _2436__36 (.A(clknet_1_0__leaf__0516_),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _2437__37 (.A(clknet_1_0__leaf__0516_),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _2438__38 (.A(clknet_1_0__leaf__0516_),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _2439__39 (.A(clknet_1_0__leaf__0516_),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _2440__40 (.A(clknet_1_1__leaf__0516_),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _2441__41 (.A(clknet_1_1__leaf__0516_),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _2442__42 (.A(clknet_1_1__leaf__0516_),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _2443__43 (.A(clknet_1_1__leaf__0516_),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _2444__44 (.A(clknet_1_1__leaf__0516_),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _2445__45 (.A(clknet_1_1__leaf__0516_),
    .Y(net106));
 sky130_fd_sc_hd__buf_1 _2446_ (.A(clknet_1_0__leaf__0514_),
    .X(_0517_));
 sky130_fd_sc_hd__inv_2 _2447__46 (.A(clknet_1_1__leaf__0517_),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _2448__47 (.A(clknet_1_1__leaf__0517_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _2449__48 (.A(clknet_1_0__leaf__0517_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _2450__49 (.A(clknet_1_0__leaf__0517_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _2451__50 (.A(clknet_1_0__leaf__0517_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _2452__51 (.A(clknet_1_0__leaf__0517_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _2453__52 (.A(clknet_1_0__leaf__0517_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _2454__53 (.A(clknet_1_0__leaf__0517_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _2455__54 (.A(clknet_1_0__leaf__0517_),
    .Y(net115));
 sky130_fd_sc_hd__inv_2 _2456__55 (.A(clknet_1_0__leaf__0517_),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _2457__56 (.A(clknet_1_1__leaf__0517_),
    .Y(net117));
 sky130_fd_sc_hd__inv_2 _2458__57 (.A(clknet_1_1__leaf__0517_),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _2459__58 (.A(clknet_1_1__leaf__0517_),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _2460__59 (.A(clknet_1_1__leaf__0517_),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _2461__60 (.A(clknet_1_1__leaf__0517_),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _2462__61 (.A(clknet_1_1__leaf__0517_),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _2463__62 (.A(clknet_1_1__leaf__0517_),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _2464__63 (.A(clknet_1_1__leaf__0517_),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _2465__64 (.A(clknet_1_1__leaf__0517_),
    .Y(net125));
 sky130_fd_sc_hd__inv_2 _2466__1 (.A(clknet_1_0__leaf__0514_),
    .Y(net62));
 sky130_fd_sc_hd__inv_2 _2467__2 (.A(clknet_1_1__leaf__0514_),
    .Y(net63));
 sky130_fd_sc_hd__inv_2 _2468__3 (.A(clknet_1_1__leaf__0514_),
    .Y(net64));
 sky130_fd_sc_hd__inv_2 _2469__4 (.A(clknet_1_1__leaf__0514_),
    .Y(net65));
 sky130_fd_sc_hd__inv_2 _2470__5 (.A(clknet_1_0__leaf__0514_),
    .Y(net66));
 sky130_fd_sc_hd__inv_2 _2471__6 (.A(clknet_1_0__leaf__0514_),
    .Y(net67));
 sky130_fd_sc_hd__inv_2 _2472__7 (.A(clknet_1_1__leaf__0514_),
    .Y(net68));
 sky130_fd_sc_hd__and3_1 _2473_ (.A(_0659_),
    .B(_0669_),
    .C(_0648_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_4 _2474_ (.A(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__inv_2 _2475_ (.A(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__and3_1 _2476_ (.A(_0903_),
    .B(_0906_),
    .C(_0519_),
    .X(_0521_));
 sky130_fd_sc_hd__a21o_1 _2477_ (.A1(\ALU.immediate[0] ),
    .A2(_0520_),
    .B1(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__nor2_1 _2478_ (.A(_0678_),
    .B(_0636_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2_1 _2479_ (.A(\ByteBuffer.instr[19] ),
    .B(_0639_),
    .Y(_0524_));
 sky130_fd_sc_hd__nor2_1 _2480_ (.A(_0678_),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_1 _2481_ (.A(\ByteBuffer.instr[20] ),
    .B(_0639_),
    .Y(_0526_));
 sky130_fd_sc_hd__nor2_1 _2482_ (.A(_0678_),
    .B(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _2483_ (.A(_0404_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__mux2_1 _2484_ (.A0(_0524_),
    .A1(_0525_),
    .S(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__xnor2_1 _2485_ (.A(_0327_),
    .B(_0525_),
    .Y(_0530_));
 sky130_fd_sc_hd__or2_1 _2486_ (.A(_0678_),
    .B(_0524_),
    .X(_0531_));
 sky130_fd_sc_hd__or4b_1 _2487_ (.A(\ByteBuffer.instr[20] ),
    .B(_0343_),
    .C(_0531_),
    .D_N(_0636_),
    .X(_0532_));
 sky130_fd_sc_hd__o41a_1 _2488_ (.A1(_0678_),
    .A2(_0636_),
    .A3(_0526_),
    .A4(_0530_),
    .B1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__o21ai_2 _2489_ (.A1(_0523_),
    .A2(_0529_),
    .B1(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__o211a_1 _2490_ (.A1(_0678_),
    .A2(_0526_),
    .B1(_0531_),
    .C1(_0523_),
    .X(_0535_));
 sky130_fd_sc_hd__and3b_1 _2491_ (.A_N(_0636_),
    .B(_0525_),
    .C(_0697_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(_0535_),
    .A1(_0536_),
    .S(_0388_),
    .X(_0537_));
 sky130_fd_sc_hd__o211a_1 _2493_ (.A1(\ByteBuffer.instr[21] ),
    .A2(_0621_),
    .B1(_0648_),
    .C1(_0647_),
    .X(_0538_));
 sky130_fd_sc_hd__or3_2 _2494_ (.A(_0525_),
    .B(_0527_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__o21ai_4 _2495_ (.A1(_0534_),
    .A2(_0537_),
    .B1(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(_0522_),
    .A1(_0455_),
    .S(net47),
    .X(_0541_));
 sky130_fd_sc_hd__nor2_8 _2497_ (.A(_0659_),
    .B(_0412_),
    .Y(_0542_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(\PC.i_mem_addr[0] ),
    .A1(_0541_),
    .S(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _2499_ (.A(_0543_),
    .X(_0158_));
 sky130_fd_sc_hd__nor2_1 _2500_ (.A(\ALU.immediate[1] ),
    .B(_0519_),
    .Y(_0544_));
 sky130_fd_sc_hd__a21oi_1 _2501_ (.A1(_0867_),
    .A2(_0519_),
    .B1(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__xor2_1 _2502_ (.A(\PC.i_mem_addr[1] ),
    .B(\PC.i_mem_addr[0] ),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(_0545_),
    .A1(_0546_),
    .S(net47),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(\PC.i_mem_addr[1] ),
    .A1(_0547_),
    .S(_0542_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_1 _2505_ (.A(_0548_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(\ALU.immediate[2] ),
    .A1(_0815_),
    .S(_0519_),
    .X(_0549_));
 sky130_fd_sc_hd__a21oi_1 _2507_ (.A1(\PC.i_mem_addr[1] ),
    .A2(\PC.i_mem_addr[0] ),
    .B1(\PC.i_mem_addr[2] ),
    .Y(_0550_));
 sky130_fd_sc_hd__and3_1 _2508_ (.A(\PC.i_mem_addr[1] ),
    .B(\PC.i_mem_addr[0] ),
    .C(\PC.i_mem_addr[2] ),
    .X(_0551_));
 sky130_fd_sc_hd__nor2_1 _2509_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(_0549_),
    .A1(_0552_),
    .S(net47),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _2511_ (.A0(\PC.i_mem_addr[2] ),
    .A1(_0553_),
    .S(_0542_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _2512_ (.A(_0554_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2513_ (.A0(\ALU.immediate[3] ),
    .A1(_0853_),
    .S(_0519_),
    .X(_0555_));
 sky130_fd_sc_hd__and2_1 _2514_ (.A(\PC.i_mem_addr[3] ),
    .B(_0551_),
    .X(_0556_));
 sky130_fd_sc_hd__nor2_1 _2515_ (.A(\PC.i_mem_addr[3] ),
    .B(_0551_),
    .Y(_0557_));
 sky130_fd_sc_hd__nor2_1 _2516_ (.A(_0556_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(_0555_),
    .A1(_0558_),
    .S(net47),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(\PC.i_mem_addr[3] ),
    .A1(_0559_),
    .S(_0542_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(_0560_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(\ALU.immediate[4] ),
    .A1(_0921_),
    .S(_0519_),
    .X(_0561_));
 sky130_fd_sc_hd__xor2_1 _2521_ (.A(\PC.i_mem_addr[4] ),
    .B(_0556_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(_0561_),
    .A1(_0562_),
    .S(net47),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(\PC.i_mem_addr[4] ),
    .A1(_0563_),
    .S(_0542_),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(_0564_),
    .X(_0162_));
 sky130_fd_sc_hd__o21a_1 _2525_ (.A1(_0630_),
    .A2(_0775_),
    .B1(_0778_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\ALU.immediate[5] ),
    .A1(_0565_),
    .S(_0519_),
    .X(_0566_));
 sky130_fd_sc_hd__and3_1 _2527_ (.A(\PC.i_mem_addr[4] ),
    .B(\PC.i_mem_addr[5] ),
    .C(_0556_),
    .X(_0567_));
 sky130_fd_sc_hd__a21oi_1 _2528_ (.A1(\PC.i_mem_addr[4] ),
    .A2(_0556_),
    .B1(\PC.i_mem_addr[5] ),
    .Y(_0568_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(_0567_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(_0566_),
    .A1(_0569_),
    .S(net47),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(\PC.i_mem_addr[5] ),
    .A1(_0570_),
    .S(_0542_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _2532_ (.A(_0571_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(\ALU.immediate[6] ),
    .A1(_0969_),
    .S(_0519_),
    .X(_0572_));
 sky130_fd_sc_hd__and2_1 _2534_ (.A(\PC.i_mem_addr[6] ),
    .B(_0567_),
    .X(_0573_));
 sky130_fd_sc_hd__nor2_1 _2535_ (.A(\PC.i_mem_addr[6] ),
    .B(_0567_),
    .Y(_0574_));
 sky130_fd_sc_hd__nor2_1 _2536_ (.A(_0573_),
    .B(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(_0572_),
    .A1(_0575_),
    .S(net47),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\PC.i_mem_addr[6] ),
    .A1(_0576_),
    .S(_0542_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(_0577_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(\ALU.immediate[7] ),
    .A1(_0946_),
    .S(_0519_),
    .X(_0578_));
 sky130_fd_sc_hd__xor2_1 _2541_ (.A(\PC.i_mem_addr[7] ),
    .B(_0573_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(_0578_),
    .A1(_0579_),
    .S(net47),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(\PC.i_mem_addr[7] ),
    .A1(_0580_),
    .S(_0542_),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_1 _2544_ (.A(_0581_),
    .X(_0165_));
 sky130_fd_sc_hd__and3_1 _2545_ (.A(\PC.i_mem_addr[7] ),
    .B(\PC.i_mem_addr[8] ),
    .C(_0573_),
    .X(_0582_));
 sky130_fd_sc_hd__inv_2 _2546_ (.A(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__a31o_1 _2547_ (.A1(\PC.i_mem_addr[6] ),
    .A2(\PC.i_mem_addr[7] ),
    .A3(_0567_),
    .B1(\PC.i_mem_addr[8] ),
    .X(_0584_));
 sky130_fd_sc_hd__o211a_2 _2548_ (.A1(_0534_),
    .A2(_0537_),
    .B1(_0520_),
    .C1(_0539_),
    .X(_0585_));
 sky130_fd_sc_hd__a32o_1 _2549_ (.A1(net47),
    .A2(_0583_),
    .A3(_0584_),
    .B1(_0585_),
    .B2(\ALU.immediate[8] ),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(\PC.i_mem_addr[8] ),
    .A1(_0586_),
    .S(_0542_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_1 _2551_ (.A(_0587_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _2552_ (.A(\PC.i_mem_addr[9] ),
    .B(_0582_),
    .X(_0588_));
 sky130_fd_sc_hd__inv_2 _2553_ (.A(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__or2_1 _2554_ (.A(\PC.i_mem_addr[9] ),
    .B(_0582_),
    .X(_0590_));
 sky130_fd_sc_hd__a32o_1 _2555_ (.A1(_0540_),
    .A2(_0589_),
    .A3(_0590_),
    .B1(_0585_),
    .B2(\ALU.immediate[9] ),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _2556_ (.A0(\PC.i_mem_addr[9] ),
    .A1(_0591_),
    .S(_0542_),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_1 _2557_ (.A(_0592_),
    .X(_0167_));
 sky130_fd_sc_hd__nand2_1 _2558_ (.A(\PC.i_mem_addr[10] ),
    .B(_0588_),
    .Y(_0593_));
 sky130_fd_sc_hd__or2_1 _2559_ (.A(\PC.i_mem_addr[10] ),
    .B(_0588_),
    .X(_0594_));
 sky130_fd_sc_hd__a32o_1 _2560_ (.A1(_0540_),
    .A2(_0593_),
    .A3(_0594_),
    .B1(_0585_),
    .B2(\ALU.immediate[10] ),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(\PC.i_mem_addr[10] ),
    .A1(_0595_),
    .S(_0542_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_1 _2562_ (.A(_0596_),
    .X(_0168_));
 sky130_fd_sc_hd__and3_1 _2563_ (.A(\PC.i_mem_addr[10] ),
    .B(\PC.i_mem_addr[11] ),
    .C(_0588_),
    .X(_0597_));
 sky130_fd_sc_hd__inv_2 _2564_ (.A(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__a31o_1 _2565_ (.A1(\PC.i_mem_addr[9] ),
    .A2(\PC.i_mem_addr[10] ),
    .A3(_0582_),
    .B1(\PC.i_mem_addr[11] ),
    .X(_0599_));
 sky130_fd_sc_hd__a32o_1 _2566_ (.A1(_0540_),
    .A2(_0598_),
    .A3(_0599_),
    .B1(_0585_),
    .B2(\ALU.immediate[11] ),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(\PC.i_mem_addr[11] ),
    .A1(_0600_),
    .S(_0542_),
    .X(_0601_));
 sky130_fd_sc_hd__clkbuf_1 _2568_ (.A(_0601_),
    .X(_0169_));
 sky130_fd_sc_hd__nand2_1 _2569_ (.A(\PC.i_mem_addr[12] ),
    .B(_0597_),
    .Y(_0602_));
 sky130_fd_sc_hd__or2_1 _2570_ (.A(\PC.i_mem_addr[12] ),
    .B(_0597_),
    .X(_0603_));
 sky130_fd_sc_hd__a32o_1 _2571_ (.A1(_0540_),
    .A2(_0602_),
    .A3(_0603_),
    .B1(_0585_),
    .B2(\ALU.immediate[12] ),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(\PC.i_mem_addr[12] ),
    .A1(_0604_),
    .S(_0542_),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_1 _2573_ (.A(_0605_),
    .X(_0170_));
 sky130_fd_sc_hd__and3_1 _2574_ (.A(\PC.i_mem_addr[12] ),
    .B(\PC.i_mem_addr[13] ),
    .C(_0597_),
    .X(_0606_));
 sky130_fd_sc_hd__inv_2 _2575_ (.A(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__a21o_1 _2576_ (.A1(\PC.i_mem_addr[12] ),
    .A2(_0597_),
    .B1(\PC.i_mem_addr[13] ),
    .X(_0608_));
 sky130_fd_sc_hd__a32o_1 _2577_ (.A1(_0540_),
    .A2(_0607_),
    .A3(_0608_),
    .B1(_0585_),
    .B2(\ALU.immediate[13] ),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(\PC.i_mem_addr[13] ),
    .A1(_0609_),
    .S(_0542_),
    .X(_0610_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_0610_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_1 _2580_ (.A(\PC.i_mem_addr[14] ),
    .B(_0606_),
    .Y(_0611_));
 sky130_fd_sc_hd__or2_1 _2581_ (.A(\PC.i_mem_addr[14] ),
    .B(_0606_),
    .X(_0612_));
 sky130_fd_sc_hd__a32o_1 _2582_ (.A1(_0540_),
    .A2(_0611_),
    .A3(_0612_),
    .B1(_0585_),
    .B2(\ALU.immediate[14] ),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(\PC.i_mem_addr[14] ),
    .A1(_0613_),
    .S(_0542_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_1 _2584_ (.A(_0614_),
    .X(_0172_));
 sky130_fd_sc_hd__xnor2_1 _2585_ (.A(\PC.i_mem_addr[15] ),
    .B(_0611_),
    .Y(_0615_));
 sky130_fd_sc_hd__a22o_1 _2586_ (.A1(\ALU.immediate[15] ),
    .A2(_0585_),
    .B1(_0615_),
    .B2(_0540_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(\PC.i_mem_addr[15] ),
    .A1(_0616_),
    .S(_0542_),
    .X(_0617_));
 sky130_fd_sc_hd__clkbuf_1 _2588_ (.A(_0617_),
    .X(_0173_));
 sky130_fd_sc_hd__dfrtp_1 _2589_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0066_),
    .RESET_B(net55),
    .Q(\MemControl.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2590_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0067_),
    .RESET_B(net55),
    .Q(\ByteDecoder.num_bytes[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2591_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0068_),
    .RESET_B(net55),
    .Q(\ByteDecoder.num_bytes[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2592_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0069_),
    .RESET_B(net55),
    .Q(\ByteDecoder.num_bytes[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2593_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0070_),
    .RESET_B(net57),
    .Q(\ALU.immediate[8] ));
 sky130_fd_sc_hd__dfrtp_4 _2594_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0071_),
    .RESET_B(net55),
    .Q(\ALU.immediate[9] ));
 sky130_fd_sc_hd__dfrtp_4 _2595_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0072_),
    .RESET_B(net55),
    .Q(\ALU.immediate[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2596_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0073_),
    .RESET_B(net57),
    .Q(\ALU.immediate[11] ));
 sky130_fd_sc_hd__dfrtp_2 _2597_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0074_),
    .RESET_B(net57),
    .Q(\ALU.immediate[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2598_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0075_),
    .RESET_B(net57),
    .Q(\ALU.immediate[13] ));
 sky130_fd_sc_hd__dfrtp_4 _2599_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0076_),
    .RESET_B(net55),
    .Q(\ALU.immediate[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2600_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0077_),
    .RESET_B(net57),
    .Q(\ALU.immediate[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2601_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0078_),
    .RESET_B(net55),
    .Q(\ByteBuffer.instr[16] ));
 sky130_fd_sc_hd__dfrtp_4 _2602_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0079_),
    .RESET_B(net55),
    .Q(\ByteBuffer.instr[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2603_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0080_),
    .RESET_B(net55),
    .Q(\ByteBuffer.instr[18] ));
 sky130_fd_sc_hd__dfrtp_4 _2604_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0081_),
    .RESET_B(net55),
    .Q(\ByteBuffer.instr[19] ));
 sky130_fd_sc_hd__dfrtp_4 _2605_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0082_),
    .RESET_B(net57),
    .Q(\ByteBuffer.instr[20] ));
 sky130_fd_sc_hd__dfrtp_4 _2606_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0083_),
    .RESET_B(net55),
    .Q(\ByteBuffer.instr[21] ));
 sky130_fd_sc_hd__dfrtp_4 _2607_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0084_),
    .RESET_B(net55),
    .Q(\ByteBuffer.instr[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2608_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0085_),
    .RESET_B(net57),
    .Q(\ByteBuffer.instr[23] ));
 sky130_fd_sc_hd__dfrtp_2 _2609_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0086_),
    .RESET_B(net55),
    .Q(\ALU.immediate[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2610_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0087_),
    .RESET_B(net56),
    .Q(\ALU.immediate[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2611_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0088_),
    .RESET_B(net56),
    .Q(\ALU.immediate[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2612_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0089_),
    .RESET_B(net56),
    .Q(\ALU.immediate[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2613_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0090_),
    .RESET_B(net57),
    .Q(\ALU.immediate[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2614_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0091_),
    .RESET_B(net56),
    .Q(\ALU.immediate[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2615_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0092_),
    .RESET_B(net56),
    .Q(\ALU.immediate[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2616_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0093_),
    .RESET_B(net57),
    .Q(\ALU.immediate[7] ));
 sky130_fd_sc_hd__dfrtp_4 _2617_ (.CLK(net69),
    .D(_0094_),
    .RESET_B(net58),
    .Q(\ALU.flags_to_alu[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2618_ (.CLK(net70),
    .D(_0095_),
    .RESET_B(net58),
    .Q(\ALU.flags_to_alu[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2619_ (.CLK(net71),
    .D(_0096_),
    .RESET_B(net58),
    .Q(\ALU.flags_to_alu[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2620_ (.CLK(net72),
    .D(_0097_),
    .RESET_B(net58),
    .Q(\ALU.flags_to_alu[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2621_ (.CLK(net73),
    .D(_0098_),
    .RESET_B(net58),
    .Q(\ALU.flags_to_alu[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2622_ (.CLK(net74),
    .D(_0099_),
    .RESET_B(net59),
    .Q(\ALU.flags_to_alu[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2623_ (.CLK(net75),
    .D(_0100_),
    .RESET_B(net58),
    .Q(\ALU.flags_to_alu[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2624_ (.CLK(net76),
    .D(_0101_),
    .RESET_B(net59),
    .Q(\ALU.flags_to_alu[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2625_ (.CLK(net77),
    .D(_0102_),
    .RESET_B(net58),
    .Q(\RegFile.L[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2626_ (.CLK(net78),
    .D(_0103_),
    .RESET_B(net59),
    .Q(\RegFile.L[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2627_ (.CLK(net79),
    .D(_0104_),
    .RESET_B(net58),
    .Q(\RegFile.L[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2628_ (.CLK(net80),
    .D(_0105_),
    .RESET_B(net59),
    .Q(\RegFile.L[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2629_ (.CLK(net81),
    .D(_0106_),
    .RESET_B(net58),
    .Q(\RegFile.L[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2630_ (.CLK(net82),
    .D(_0107_),
    .RESET_B(net59),
    .Q(\RegFile.L[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2631_ (.CLK(net83),
    .D(_0108_),
    .RESET_B(net59),
    .Q(\RegFile.L[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2632_ (.CLK(net84),
    .D(_0109_),
    .RESET_B(net59),
    .Q(\RegFile.L[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2633_ (.CLK(net85),
    .D(_0110_),
    .RESET_B(net60),
    .Q(\RegFile.H[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2634_ (.CLK(net86),
    .D(_0111_),
    .RESET_B(net60),
    .Q(\RegFile.H[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2635_ (.CLK(net87),
    .D(_0112_),
    .RESET_B(net60),
    .Q(\RegFile.H[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2636_ (.CLK(net88),
    .D(_0113_),
    .RESET_B(net60),
    .Q(\RegFile.H[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2637_ (.CLK(net89),
    .D(_0114_),
    .RESET_B(net60),
    .Q(\RegFile.H[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2638_ (.CLK(net90),
    .D(_0115_),
    .RESET_B(net60),
    .Q(\RegFile.H[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2639_ (.CLK(net91),
    .D(_0116_),
    .RESET_B(net60),
    .Q(\RegFile.H[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2640_ (.CLK(net92),
    .D(_0117_),
    .RESET_B(net60),
    .Q(\RegFile.H[7] ));
 sky130_fd_sc_hd__dfrtp_4 _2641_ (.CLK(net93),
    .D(_0118_),
    .RESET_B(net58),
    .Q(\RegFile.E[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2642_ (.CLK(net94),
    .D(_0119_),
    .RESET_B(net59),
    .Q(\RegFile.E[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2643_ (.CLK(net95),
    .D(_0120_),
    .RESET_B(net58),
    .Q(\RegFile.E[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2644_ (.CLK(net96),
    .D(_0121_),
    .RESET_B(net59),
    .Q(\RegFile.E[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2645_ (.CLK(net97),
    .D(_0122_),
    .RESET_B(net58),
    .Q(\RegFile.E[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2646_ (.CLK(net98),
    .D(_0123_),
    .RESET_B(net59),
    .Q(\RegFile.E[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2647_ (.CLK(net99),
    .D(_0124_),
    .RESET_B(net59),
    .Q(\RegFile.E[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2648_ (.CLK(net100),
    .D(_0125_),
    .RESET_B(net60),
    .Q(\RegFile.E[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2649_ (.CLK(net101),
    .D(_0126_),
    .RESET_B(net60),
    .Q(\RegFile.D[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2650_ (.CLK(net102),
    .D(_0127_),
    .RESET_B(net60),
    .Q(\RegFile.D[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2651_ (.CLK(net103),
    .D(_0128_),
    .RESET_B(net60),
    .Q(\RegFile.D[2] ));
 sky130_fd_sc_hd__dfrtp_4 _2652_ (.CLK(net104),
    .D(_0129_),
    .RESET_B(net61),
    .Q(\RegFile.D[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2653_ (.CLK(net105),
    .D(_0130_),
    .RESET_B(net60),
    .Q(\RegFile.D[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2654_ (.CLK(net106),
    .D(_0131_),
    .RESET_B(net61),
    .Q(\RegFile.D[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2655_ (.CLK(net107),
    .D(_0132_),
    .RESET_B(net61),
    .Q(\RegFile.D[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2656_ (.CLK(net108),
    .D(_0133_),
    .RESET_B(net61),
    .Q(\RegFile.D[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2657_ (.CLK(net109),
    .D(_0134_),
    .RESET_B(net58),
    .Q(\RegFile.C[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2658_ (.CLK(net110),
    .D(_0135_),
    .RESET_B(net59),
    .Q(\RegFile.C[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2659_ (.CLK(net111),
    .D(_0136_),
    .RESET_B(net58),
    .Q(\RegFile.C[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2660_ (.CLK(net112),
    .D(_0137_),
    .RESET_B(net59),
    .Q(\RegFile.C[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2661_ (.CLK(net113),
    .D(_0138_),
    .RESET_B(net58),
    .Q(\RegFile.C[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2662_ (.CLK(net114),
    .D(_0139_),
    .RESET_B(net59),
    .Q(\RegFile.C[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2663_ (.CLK(net115),
    .D(_0140_),
    .RESET_B(net59),
    .Q(\RegFile.C[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2664_ (.CLK(net116),
    .D(_0141_),
    .RESET_B(net59),
    .Q(\RegFile.C[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2665_ (.CLK(net117),
    .D(_0142_),
    .RESET_B(net60),
    .Q(\RegFile.B[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2666_ (.CLK(net118),
    .D(_0143_),
    .RESET_B(net61),
    .Q(\RegFile.B[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2667_ (.CLK(net119),
    .D(_0144_),
    .RESET_B(net60),
    .Q(\RegFile.B[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2668_ (.CLK(net120),
    .D(_0145_),
    .RESET_B(net61),
    .Q(\RegFile.B[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2669_ (.CLK(net121),
    .D(_0146_),
    .RESET_B(net60),
    .Q(\RegFile.B[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2670_ (.CLK(net122),
    .D(_0147_),
    .RESET_B(net61),
    .Q(\RegFile.B[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2671_ (.CLK(net123),
    .D(_0148_),
    .RESET_B(net61),
    .Q(\RegFile.B[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2672_ (.CLK(net124),
    .D(_0149_),
    .RESET_B(net61),
    .Q(\RegFile.B[7] ));
 sky130_fd_sc_hd__dfrtp_4 _2673_ (.CLK(net125),
    .D(_0150_),
    .RESET_B(net60),
    .Q(\RegFile.A[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2674_ (.CLK(net62),
    .D(_0151_),
    .RESET_B(net61),
    .Q(\RegFile.A[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2675_ (.CLK(net63),
    .D(_0152_),
    .RESET_B(net60),
    .Q(\RegFile.A[2] ));
 sky130_fd_sc_hd__dfrtp_4 _2676_ (.CLK(net64),
    .D(_0153_),
    .RESET_B(net60),
    .Q(\RegFile.A[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2677_ (.CLK(net65),
    .D(_0154_),
    .RESET_B(net60),
    .Q(\RegFile.A[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2678_ (.CLK(net66),
    .D(_0155_),
    .RESET_B(net61),
    .Q(\RegFile.A[5] ));
 sky130_fd_sc_hd__dfrtp_4 _2679_ (.CLK(net67),
    .D(_0156_),
    .RESET_B(net61),
    .Q(\RegFile.A[6] ));
 sky130_fd_sc_hd__dfrtp_4 _2680_ (.CLK(net68),
    .D(_0157_),
    .RESET_B(net61),
    .Q(\RegFile.A[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2681_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0158_),
    .RESET_B(net55),
    .Q(\PC.i_mem_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2682_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0159_),
    .RESET_B(net55),
    .Q(\PC.i_mem_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2683_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0160_),
    .RESET_B(net55),
    .Q(\PC.i_mem_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2684_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0161_),
    .RESET_B(net55),
    .Q(\PC.i_mem_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2685_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0162_),
    .RESET_B(net55),
    .Q(\PC.i_mem_addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2686_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0163_),
    .RESET_B(net57),
    .Q(\PC.i_mem_addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2687_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0164_),
    .RESET_B(net57),
    .Q(\PC.i_mem_addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2688_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0165_),
    .RESET_B(net57),
    .Q(\PC.i_mem_addr[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2689_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0166_),
    .RESET_B(net57),
    .Q(\PC.i_mem_addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2690_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0167_),
    .RESET_B(net57),
    .Q(\PC.i_mem_addr[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2691_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0168_),
    .RESET_B(net58),
    .Q(\PC.i_mem_addr[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2692_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0169_),
    .RESET_B(net58),
    .Q(\PC.i_mem_addr[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2693_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0170_),
    .RESET_B(net58),
    .Q(\PC.i_mem_addr[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2694_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0171_),
    .RESET_B(net58),
    .Q(\PC.i_mem_addr[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2695_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0172_),
    .RESET_B(net58),
    .Q(\PC.i_mem_addr[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2696_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0173_),
    .RESET_B(net57),
    .Q(\PC.i_mem_addr[15] ));
 sky130_fd_sc_hd__dfstp_1 _2697_ (.CLK(clknet_2_3__leaf_clk),
    .D(net134),
    .SET_B(net56),
    .Q(\MemControl.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2698_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0001_),
    .RESET_B(net56),
    .Q(\MemControl.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2699_ (.CLK(clknet_2_3__leaf_clk),
    .D(net130),
    .RESET_B(net56),
    .Q(\ByteDecoder.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2700_ (.CLK(clknet_2_3__leaf_clk),
    .D(\FSM.next_state[1] ),
    .RESET_B(net56),
    .Q(\ByteDecoder.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2701_ (.CLK(clknet_2_3__leaf_clk),
    .D(\ByteBuffer.next_counter[0] ),
    .RESET_B(net56),
    .Q(\ByteBuffer.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2702_ (.CLK(clknet_2_3__leaf_clk),
    .D(\ByteBuffer.next_counter[1] ),
    .RESET_B(net55),
    .Q(\ByteBuffer.counter[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0514_ (.A(_0514_),
    .X(clknet_0__0514_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0515_ (.A(_0515_),
    .X(clknet_0__0515_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0516_ (.A(_0516_),
    .X(clknet_0__0516_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0517_ (.A(_0517_),
    .X(clknet_0__0517_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0514_ (.A(clknet_0__0514_),
    .X(clknet_1_0__leaf__0514_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0515_ (.A(clknet_0__0515_),
    .X(clknet_1_0__leaf__0515_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0516_ (.A(clknet_0__0516_),
    .X(clknet_1_0__leaf__0516_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0517_ (.A(clknet_0__0517_),
    .X(clknet_1_0__leaf__0517_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0514_ (.A(clknet_0__0514_),
    .X(clknet_1_1__leaf__0514_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0515_ (.A(clknet_0__0515_),
    .X(clknet_1_1__leaf__0515_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0516_ (.A(clknet_0__0516_),
    .X(clknet_1_1__leaf__0516_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0517_ (.A(clknet_0__0517_),
    .X(clknet_1_1__leaf__0517_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__buf_8 fanout55 (.A(net57),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__buf_6 fanout57 (.A(net11),
    .X(net57));
 sky130_fd_sc_hd__buf_6 fanout58 (.A(net11),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 fanout59 (.A(net11),
    .X(net59));
 sky130_fd_sc_hd__buf_8 fanout60 (.A(net11),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(net11),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\ByteDecoder.num_bytes[2] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\ALU.flags_to_alu[3] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\ALU.flags_to_alu[4] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\ALU.flags_to_alu[6] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\ALU.flags_to_alu[5] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\ByteDecoder.state[1] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\ByteDecoder.num_bytes[3] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\ByteBuffer.counter[0] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\ByteDecoder.num_bytes[1] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\FSM.next_state[0] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\MemControl.state[2] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\ALU.flags_to_alu[1] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\MemControl.state[1] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0000_),
    .X(net134));
 sky130_fd_sc_hd__buf_4 input1 (.A(cs),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(gpi[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(nrst),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(gpi[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(gpi[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(gpi[23]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(gpi[2]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(gpi[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(gpi[4]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(gpi[5]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(gpi[6]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 max_cap47 (.A(_0540_),
    .X(net47));
 sky130_fd_sc_hd__buf_6 max_cap48 (.A(_1043_),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 max_cap49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__buf_4 max_cap51 (.A(_0685_),
    .X(net51));
 sky130_fd_sc_hd__buf_4 max_cap52 (.A(_0680_),
    .X(net52));
 sky130_fd_sc_hd__buf_4 max_cap53 (.A(_0706_),
    .X(net53));
 sky130_fd_sc_hd__buf_2 max_cap54 (.A(_0646_),
    .X(net54));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(gpo[0]));
 sky130_fd_sc_hd__clkbuf_4 output13 (.A(net13),
    .X(gpo[10]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(gpo[11]));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(gpo[12]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(gpo[13]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(gpo[14]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(gpo[15]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(gpo[16]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(gpo[17]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(gpo[18]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(gpo[19]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(gpo[1]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(gpo[20]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(gpo[21]));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net26),
    .X(gpo[22]));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net27),
    .X(gpo[23]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(gpo[24]));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net29),
    .X(gpo[25]));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net30),
    .X(gpo[26]));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net31),
    .X(gpo[27]));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net32),
    .X(gpo[28]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(gpo[29]));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net34),
    .X(gpo[2]));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net35),
    .X(gpo[30]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(gpo[31]));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(gpo[32]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(gpo[33]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(gpo[3]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(gpo[4]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(gpo[5]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(gpo[6]));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(gpo[7]));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net44),
    .X(gpo[8]));
 sky130_fd_sc_hd__clkbuf_4 output45 (.A(net45),
    .X(gpo[9]));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(store_en));
 sky130_fd_sc_hd__clkbuf_2 wire50 (.A(_0772_),
    .X(net50));
endmodule

