magic
tech sky130A
magscale 1 2
timestamp 1693936176
<< obsli1 >>
rect 1104 2159 147016 147985
<< obsm1 >>
rect 14 2128 147076 148016
<< metal2 >>
rect 2594 149514 2650 150314
rect 20626 149514 20682 150314
rect 38658 149514 38714 150314
rect 57334 149514 57390 150314
rect 75366 149514 75422 150314
rect 93398 149514 93454 150314
rect 111430 149514 111486 150314
rect 129462 149514 129518 150314
rect 147494 149514 147550 150314
rect 18 0 74 800
rect 18050 0 18106 800
rect 36082 0 36138 800
rect 54114 0 54170 800
rect 72146 0 72202 800
rect 90178 0 90234 800
rect 108854 0 108910 800
rect 126886 0 126942 800
rect 144918 0 144974 800
<< obsm2 >>
rect 20 149458 2538 149514
rect 2706 149458 20570 149514
rect 20738 149458 38602 149514
rect 38770 149458 57278 149514
rect 57446 149458 75310 149514
rect 75478 149458 93342 149514
rect 93510 149458 111374 149514
rect 111542 149458 129406 149514
rect 129574 149458 147438 149514
rect 20 856 147550 149458
rect 130 800 17994 856
rect 18162 800 36026 856
rect 36194 800 54058 856
rect 54226 800 72090 856
rect 72258 800 90122 856
rect 90290 800 108798 856
rect 108966 800 126830 856
rect 126998 800 144862 856
rect 145030 800 147550 856
<< metal3 >>
rect 0 133968 800 134088
rect 147370 130568 148170 130688
rect 0 114928 800 115048
rect 147370 111528 148170 111648
rect 0 95208 800 95328
rect 147370 92488 148170 92608
rect 0 76168 800 76288
rect 147370 73448 148170 73568
rect 0 57128 800 57248
rect 147370 54408 148170 54528
rect 0 38088 800 38208
rect 147370 34688 148170 34808
rect 0 19048 800 19168
rect 147370 15648 148170 15768
<< obsm3 >>
rect 800 134168 147555 148001
rect 880 133888 147555 134168
rect 800 130768 147555 133888
rect 800 130488 147290 130768
rect 800 115128 147555 130488
rect 880 114848 147555 115128
rect 800 111728 147555 114848
rect 800 111448 147290 111728
rect 800 95408 147555 111448
rect 880 95128 147555 95408
rect 800 92688 147555 95128
rect 800 92408 147290 92688
rect 800 76368 147555 92408
rect 880 76088 147555 76368
rect 800 73648 147555 76088
rect 800 73368 147290 73648
rect 800 57328 147555 73368
rect 880 57048 147555 57328
rect 800 54608 147555 57048
rect 800 54328 147290 54608
rect 800 38288 147555 54328
rect 880 38008 147555 38288
rect 800 34888 147555 38008
rect 800 34608 147290 34888
rect 800 19248 147555 34608
rect 880 18968 147555 19248
rect 800 15848 147555 18968
rect 800 15568 147290 15848
rect 800 2143 147555 15568
<< metal4 >>
rect 4208 2128 4528 148016
rect 19568 2128 19888 148016
rect 34928 2128 35248 148016
rect 50288 2128 50608 148016
rect 65648 2128 65968 148016
rect 81008 2128 81328 148016
rect 96368 2128 96688 148016
rect 111728 2128 112048 148016
rect 127088 2128 127408 148016
rect 142448 2128 142768 148016
<< obsm4 >>
rect 3838 2619 4128 147797
rect 4608 2619 19488 147797
rect 19968 2619 34848 147797
rect 35328 2619 50208 147797
rect 50688 2619 65568 147797
rect 66048 2619 80928 147797
rect 81408 2619 96288 147797
rect 96768 2619 111648 147797
rect 112128 2619 127008 147797
rect 127488 2619 142368 147797
rect 142848 2619 146490 147797
<< obsm5 >>
rect 3796 21260 146532 138540
<< labels >>
rlabel metal2 s 147494 149514 147550 150314 6 clk
port 1 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 color[0]
port 2 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 color[10]
port 3 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 color[11]
port 4 nsew signal output
rlabel metal2 s 38658 149514 38714 150314 6 color[12]
port 5 nsew signal output
rlabel metal2 s 93398 149514 93454 150314 6 color[13]
port 6 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 color[14]
port 7 nsew signal output
rlabel metal3 s 147370 73448 148170 73568 6 color[15]
port 8 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 color[16]
port 9 nsew signal output
rlabel metal3 s 147370 92488 148170 92608 6 color[17]
port 10 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 color[18]
port 11 nsew signal output
rlabel metal2 s 18 0 74 800 6 color[19]
port 12 nsew signal output
rlabel metal2 s 111430 149514 111486 150314 6 color[1]
port 13 nsew signal output
rlabel metal2 s 129462 149514 129518 150314 6 color[20]
port 14 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 color[21]
port 15 nsew signal output
rlabel metal3 s 147370 15648 148170 15768 6 color[22]
port 16 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 color[23]
port 17 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 color[2]
port 18 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 color[3]
port 19 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 color[4]
port 20 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 color[5]
port 21 nsew signal output
rlabel metal2 s 20626 149514 20682 150314 6 color[6]
port 22 nsew signal output
rlabel metal3 s 147370 34688 148170 34808 6 color[7]
port 23 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 color[8]
port 24 nsew signal output
rlabel metal3 s 147370 111528 148170 111648 6 color[9]
port 25 nsew signal output
rlabel metal3 s 147370 130568 148170 130688 6 cs
port 26 nsew signal input
rlabel metal2 s 57334 149514 57390 150314 6 is_mandelbrot
port 27 nsew signal output
rlabel metal2 s 75366 149514 75422 150314 6 nrst
port 28 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 spi_clk
port 29 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 spi_data
port 30 nsew signal input
rlabel metal2 s 2594 149514 2650 150314 6 spi_en
port 31 nsew signal input
rlabel metal3 s 147370 54408 148170 54528 6 valid_out
port 32 nsew signal output
rlabel metal4 s 4208 2128 4528 148016 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 148016 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 148016 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 148016 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 148016 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 148016 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 148016 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 148016 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 148016 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 148016 6 vssd1
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 148170 150314
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 67229252
string GDS_FILE /home/designer-05/work/Caravel_STARS_2023/openlane/DigiDoggs/runs/23_09_05_10_15/results/signoff/pushing_pixels.magic.gds
string GDS_START 1578934
<< end >>

