magic
tech sky130A
magscale 1 2
timestamp 1694009411
<< viali >>
rect 1593 39049 1627 39083
rect 4997 39049 5031 39083
rect 9505 39049 9539 39083
rect 11713 39049 11747 39083
rect 13185 39049 13219 39083
rect 17877 39049 17911 39083
rect 22201 39049 22235 39083
rect 27169 39049 27203 39083
rect 33149 39049 33183 39083
rect 15669 38981 15703 39015
rect 31125 38981 31159 39015
rect 36001 38981 36035 39015
rect 1501 38913 1535 38947
rect 4813 38913 4847 38947
rect 9321 38913 9355 38947
rect 11621 38913 11655 38947
rect 12265 38913 12299 38947
rect 12725 38913 12759 38947
rect 13001 38913 13035 38947
rect 17693 38913 17727 38947
rect 20085 38913 20119 38947
rect 22109 38913 22143 38947
rect 24777 38913 24811 38947
rect 25881 38913 25915 38947
rect 27077 38913 27111 38947
rect 33057 38913 33091 38947
rect 35633 38913 35667 38947
rect 37473 38913 37507 38947
rect 20361 38845 20395 38879
rect 26157 38845 26191 38879
rect 37657 38777 37691 38811
rect 12357 38709 12391 38743
rect 12541 38709 12575 38743
rect 15761 38709 15795 38743
rect 24869 38709 24903 38743
rect 31217 38709 31251 38743
rect 4997 38505 5031 38539
rect 9321 38505 9355 38539
rect 12344 38505 12378 38539
rect 24409 38505 24443 38539
rect 32137 38505 32171 38539
rect 34713 38505 34747 38539
rect 37841 38505 37875 38539
rect 12081 38369 12115 38403
rect 22753 38369 22787 38403
rect 24685 38369 24719 38403
rect 28733 38369 28767 38403
rect 5181 38301 5215 38335
rect 8493 38301 8527 38335
rect 9505 38301 9539 38335
rect 9873 38301 9907 38335
rect 9965 38301 9999 38335
rect 10149 38301 10183 38335
rect 20177 38301 20211 38335
rect 20269 38301 20303 38335
rect 20361 38301 20395 38335
rect 20545 38301 20579 38335
rect 22569 38301 22603 38335
rect 24593 38301 24627 38335
rect 26709 38301 26743 38335
rect 26801 38301 26835 38335
rect 26985 38301 27019 38335
rect 29193 38301 29227 38335
rect 29285 38301 29319 38335
rect 29561 38301 29595 38335
rect 31861 38301 31895 38335
rect 32321 38301 32355 38335
rect 34897 38301 34931 38335
rect 10425 38233 10459 38267
rect 20821 38233 20855 38267
rect 24961 38233 24995 38267
rect 27261 38233 27295 38267
rect 29837 38233 29871 38267
rect 37565 38233 37599 38267
rect 8585 38165 8619 38199
rect 11897 38165 11931 38199
rect 13829 38165 13863 38199
rect 19993 38165 20027 38199
rect 22293 38165 22327 38199
rect 26433 38165 26467 38199
rect 31309 38165 31343 38199
rect 31953 38165 31987 38199
rect 10333 37961 10367 37995
rect 11069 37961 11103 37995
rect 11529 37961 11563 37995
rect 12265 37961 12299 37995
rect 14657 37961 14691 37995
rect 17877 37961 17911 37995
rect 20453 37961 20487 37995
rect 22109 37961 22143 37995
rect 25513 37961 25547 37995
rect 26617 37961 26651 37995
rect 28825 37961 28859 37995
rect 29285 37961 29319 37995
rect 29653 37961 29687 37995
rect 12633 37893 12667 37927
rect 17509 37893 17543 37927
rect 17601 37893 17635 37927
rect 18245 37893 18279 37927
rect 18613 37893 18647 37927
rect 18981 37893 19015 37927
rect 20821 37893 20855 37927
rect 21465 37893 21499 37927
rect 26157 37893 26191 37927
rect 26249 37893 26283 37927
rect 8401 37825 8435 37859
rect 10517 37825 10551 37859
rect 10977 37825 11011 37859
rect 11713 37825 11747 37859
rect 14105 37825 14139 37859
rect 14289 37825 14323 37859
rect 14565 37825 14599 37859
rect 14749 37825 14783 37859
rect 14933 37825 14967 37859
rect 15577 37825 15611 37859
rect 15669 37825 15703 37859
rect 15853 37825 15887 37859
rect 15945 37825 15979 37859
rect 16037 37825 16071 37859
rect 17325 37825 17359 37859
rect 17693 37825 17727 37859
rect 18429 37825 18463 37859
rect 18797 37825 18831 37859
rect 19073 37825 19107 37859
rect 19165 37825 19199 37859
rect 19441 37825 19475 37859
rect 19625 37825 19659 37859
rect 21281 37825 21315 37859
rect 22017 37825 22051 37859
rect 22201 37825 22235 37859
rect 22569 37825 22603 37859
rect 22753 37825 22787 37859
rect 22845 37825 22879 37859
rect 22937 37825 22971 37859
rect 24777 37825 24811 37859
rect 24961 37825 24995 37859
rect 25237 37825 25271 37859
rect 25421 37825 25455 37859
rect 25697 37825 25731 37859
rect 26801 37825 26835 37859
rect 27445 37825 27479 37859
rect 27997 37825 28031 37859
rect 28089 37825 28123 37859
rect 29193 37825 29227 37859
rect 29837 37825 29871 37859
rect 30021 37825 30055 37859
rect 32321 37825 32355 37859
rect 8677 37757 8711 37791
rect 11161 37757 11195 37791
rect 12725 37757 12759 37791
rect 12909 37757 12943 37791
rect 13921 37757 13955 37791
rect 20913 37757 20947 37791
rect 21005 37757 21039 37791
rect 24593 37757 24627 37791
rect 25053 37757 25087 37791
rect 26433 37757 26467 37791
rect 27537 37757 27571 37791
rect 27629 37757 27663 37791
rect 29377 37757 29411 37791
rect 30297 37757 30331 37791
rect 10609 37689 10643 37723
rect 14381 37689 14415 37723
rect 21833 37689 21867 37723
rect 25789 37689 25823 37723
rect 27077 37689 27111 37723
rect 28273 37689 28307 37723
rect 32137 37689 32171 37723
rect 10149 37621 10183 37655
rect 15577 37621 15611 37655
rect 19349 37621 19383 37655
rect 19809 37621 19843 37655
rect 21649 37621 21683 37655
rect 22385 37621 22419 37655
rect 23121 37621 23155 37655
rect 31769 37621 31803 37655
rect 8953 37417 8987 37451
rect 19441 37417 19475 37451
rect 23581 37417 23615 37451
rect 25145 37417 25179 37451
rect 1777 37281 1811 37315
rect 10057 37281 10091 37315
rect 19533 37281 19567 37315
rect 24777 37281 24811 37315
rect 26985 37281 27019 37315
rect 31217 37281 31251 37315
rect 31309 37281 31343 37315
rect 9137 37213 9171 37247
rect 9873 37213 9907 37247
rect 14289 37213 14323 37247
rect 19717 37213 19751 37247
rect 21925 37213 21959 37247
rect 22109 37213 22143 37247
rect 22201 37213 22235 37247
rect 22293 37213 22327 37247
rect 22569 37213 22603 37247
rect 22662 37213 22696 37247
rect 23075 37213 23109 37247
rect 23765 37213 23799 37247
rect 23857 37213 23891 37247
rect 24961 37213 24995 37247
rect 27169 37213 27203 37247
rect 27353 37213 27387 37247
rect 37657 37213 37691 37247
rect 1501 37145 1535 37179
rect 15117 37145 15151 37179
rect 19441 37145 19475 37179
rect 22845 37145 22879 37179
rect 22937 37145 22971 37179
rect 23581 37145 23615 37179
rect 37289 37145 37323 37179
rect 9505 37077 9539 37111
rect 9965 37077 9999 37111
rect 19901 37077 19935 37111
rect 22477 37077 22511 37111
rect 23213 37077 23247 37111
rect 24041 37077 24075 37111
rect 30757 37077 30791 37111
rect 31125 37077 31159 37111
rect 37841 37077 37875 37111
rect 23121 36873 23155 36907
rect 15945 36805 15979 36839
rect 25513 36805 25547 36839
rect 7021 36737 7055 36771
rect 16129 36737 16163 36771
rect 16221 36737 16255 36771
rect 16318 36737 16352 36771
rect 22937 36737 22971 36771
rect 25237 36737 25271 36771
rect 25421 36737 25455 36771
rect 25605 36737 25639 36771
rect 27629 36737 27663 36771
rect 32965 36737 32999 36771
rect 22753 36669 22787 36703
rect 7113 36533 7147 36567
rect 15945 36533 15979 36567
rect 25789 36533 25823 36567
rect 27721 36533 27755 36567
rect 32781 36533 32815 36567
rect 19073 36329 19107 36363
rect 20913 36329 20947 36363
rect 23489 36329 23523 36363
rect 12817 36261 12851 36295
rect 13553 36261 13587 36295
rect 26157 36261 26191 36295
rect 29285 36261 29319 36295
rect 30205 36261 30239 36295
rect 6929 36193 6963 36227
rect 10701 36193 10735 36227
rect 27537 36193 27571 36227
rect 32781 36193 32815 36227
rect 4721 36125 4755 36159
rect 4813 36125 4847 36159
rect 4997 36125 5031 36159
rect 8953 36125 8987 36159
rect 12265 36125 12299 36159
rect 12541 36125 12575 36159
rect 12633 36125 12667 36159
rect 13123 36125 13157 36159
rect 13645 36125 13679 36159
rect 15117 36125 15151 36159
rect 15209 36125 15243 36159
rect 15301 36125 15335 36159
rect 15577 36125 15611 36159
rect 17417 36125 17451 36159
rect 17693 36125 17727 36159
rect 17785 36125 17819 36159
rect 18061 36125 18095 36159
rect 18245 36125 18279 36159
rect 18429 36125 18463 36159
rect 18522 36125 18556 36159
rect 18797 36125 18831 36159
rect 18894 36125 18928 36159
rect 19717 36125 19751 36159
rect 19809 36125 19843 36159
rect 20085 36125 20119 36159
rect 20177 36125 20211 36159
rect 20361 36125 20395 36159
rect 20637 36125 20671 36159
rect 20729 36125 20763 36159
rect 22937 36125 22971 36159
rect 23121 36125 23155 36159
rect 23213 36125 23247 36159
rect 23305 36125 23339 36159
rect 25145 36125 25179 36159
rect 25237 36125 25271 36159
rect 25421 36125 25455 36159
rect 25513 36125 25547 36159
rect 25605 36125 25639 36159
rect 25973 36125 26007 36159
rect 26341 36125 26375 36159
rect 26434 36125 26468 36159
rect 26709 36125 26743 36159
rect 26806 36125 26840 36159
rect 27445 36125 27479 36159
rect 29561 36125 29595 36159
rect 29654 36125 29688 36159
rect 29929 36125 29963 36159
rect 30026 36125 30060 36159
rect 30297 36125 30331 36159
rect 30941 36125 30975 36159
rect 32229 36125 32263 36159
rect 32321 36125 32355 36159
rect 32505 36125 32539 36159
rect 5273 36057 5307 36091
rect 7205 36057 7239 36091
rect 9229 36057 9263 36091
rect 12449 36057 12483 36091
rect 15419 36057 15453 36091
rect 17601 36057 17635 36091
rect 18705 36057 18739 36091
rect 19993 36057 20027 36091
rect 20545 36057 20579 36091
rect 25789 36057 25823 36091
rect 25881 36057 25915 36091
rect 26617 36057 26651 36091
rect 27813 36057 27847 36091
rect 29837 36057 29871 36091
rect 6745 35989 6779 36023
rect 8677 35989 8711 36023
rect 13001 35989 13035 36023
rect 13185 35989 13219 36023
rect 14933 35989 14967 36023
rect 17969 35989 18003 36023
rect 18245 35989 18279 36023
rect 19717 35989 19751 36023
rect 24961 35989 24995 36023
rect 26985 35989 27019 36023
rect 27261 35989 27295 36023
rect 30389 35989 30423 36023
rect 30757 35989 30791 36023
rect 34253 35989 34287 36023
rect 5549 35785 5583 35819
rect 7481 35785 7515 35819
rect 7849 35785 7883 35819
rect 8217 35785 8251 35819
rect 9137 35785 9171 35819
rect 9321 35785 9355 35819
rect 10241 35785 10275 35819
rect 13553 35785 13587 35819
rect 14841 35785 14875 35819
rect 27261 35785 27295 35819
rect 32781 35785 32815 35819
rect 33149 35785 33183 35819
rect 33241 35785 33275 35819
rect 6377 35717 6411 35751
rect 11989 35717 12023 35751
rect 25237 35717 25271 35751
rect 29653 35717 29687 35751
rect 5733 35649 5767 35683
rect 7665 35649 7699 35683
rect 8309 35649 8343 35683
rect 9045 35649 9079 35683
rect 9505 35649 9539 35683
rect 10149 35649 10183 35683
rect 10793 35649 10827 35683
rect 11897 35649 11931 35683
rect 12909 35649 12943 35683
rect 13002 35649 13036 35683
rect 13139 35649 13173 35683
rect 13277 35649 13311 35683
rect 13374 35649 13408 35683
rect 14749 35649 14783 35683
rect 22109 35649 22143 35683
rect 22293 35649 22327 35683
rect 22385 35649 22419 35683
rect 22477 35649 22511 35683
rect 22753 35649 22787 35683
rect 22846 35649 22880 35683
rect 23029 35649 23063 35683
rect 23121 35649 23155 35683
rect 23218 35649 23252 35683
rect 25421 35649 25455 35683
rect 25513 35649 25547 35683
rect 25697 35649 25731 35683
rect 25789 35649 25823 35683
rect 27629 35649 27663 35683
rect 29469 35649 29503 35683
rect 29745 35649 29779 35683
rect 30113 35649 30147 35683
rect 7205 35581 7239 35615
rect 8401 35581 8435 35615
rect 10425 35581 10459 35615
rect 12173 35581 12207 35615
rect 27721 35581 27755 35615
rect 27905 35581 27939 35615
rect 30389 35581 30423 35615
rect 33333 35581 33367 35615
rect 9781 35513 9815 35547
rect 11529 35513 11563 35547
rect 10609 35445 10643 35479
rect 22661 35445 22695 35479
rect 23397 35445 23431 35479
rect 29285 35445 29319 35479
rect 31861 35445 31895 35479
rect 6009 35241 6043 35275
rect 11989 35241 12023 35275
rect 27813 35241 27847 35275
rect 30665 35241 30699 35275
rect 14105 35173 14139 35207
rect 25421 35173 25455 35207
rect 6561 35105 6595 35139
rect 10517 35105 10551 35139
rect 23489 35105 23523 35139
rect 23581 35105 23615 35139
rect 27169 35105 27203 35139
rect 31309 35105 31343 35139
rect 4445 35037 4479 35071
rect 7941 35037 7975 35071
rect 9965 35037 9999 35071
rect 10057 35037 10091 35071
rect 10241 35037 10275 35071
rect 14289 35037 14323 35071
rect 14473 35037 14507 35071
rect 19441 35037 19475 35071
rect 19625 35037 19659 35071
rect 19901 35037 19935 35071
rect 21005 35037 21039 35071
rect 21098 35037 21132 35071
rect 21373 35037 21407 35071
rect 21470 35037 21504 35071
rect 22201 35037 22235 35071
rect 22294 35037 22328 35071
rect 22477 35037 22511 35071
rect 22707 35037 22741 35071
rect 23305 35037 23339 35071
rect 23397 35037 23431 35071
rect 23765 35037 23799 35071
rect 24961 35037 24995 35071
rect 25053 35037 25087 35071
rect 25145 35037 25179 35071
rect 25329 35037 25363 35071
rect 25697 35037 25731 35071
rect 25789 35037 25823 35071
rect 25881 35037 25915 35071
rect 26065 35037 26099 35071
rect 27353 35037 27387 35071
rect 27537 35037 27571 35071
rect 27626 35015 27660 35049
rect 27721 35037 27755 35071
rect 31033 35037 31067 35071
rect 6377 34969 6411 35003
rect 19533 34969 19567 35003
rect 19763 34969 19797 35003
rect 21281 34969 21315 35003
rect 22569 34969 22603 35003
rect 4537 34901 4571 34935
rect 6469 34901 6503 34935
rect 8033 34901 8067 34935
rect 14381 34901 14415 34935
rect 14657 34901 14691 34935
rect 19257 34901 19291 34935
rect 21649 34901 21683 34935
rect 22845 34901 22879 34935
rect 23121 34901 23155 34935
rect 24685 34901 24719 34935
rect 31125 34901 31159 34935
rect 6745 34697 6779 34731
rect 9597 34697 9631 34731
rect 16865 34697 16899 34731
rect 20821 34697 20855 34731
rect 24041 34697 24075 34731
rect 30941 34697 30975 34731
rect 12541 34629 12575 34663
rect 17233 34629 17267 34663
rect 17417 34629 17451 34663
rect 20085 34629 20119 34663
rect 20453 34629 20487 34663
rect 20653 34629 20687 34663
rect 23673 34629 23707 34663
rect 29377 34629 29411 34663
rect 4353 34561 4387 34595
rect 6837 34561 6871 34595
rect 7849 34561 7883 34595
rect 12173 34561 12207 34595
rect 12266 34561 12300 34595
rect 12449 34561 12483 34595
rect 12679 34561 12713 34595
rect 17141 34561 17175 34595
rect 17601 34561 17635 34595
rect 17693 34561 17727 34595
rect 17785 34561 17819 34595
rect 19901 34561 19935 34595
rect 20177 34561 20211 34595
rect 20305 34561 20339 34595
rect 22017 34561 22051 34595
rect 22109 34561 22143 34595
rect 22293 34561 22327 34595
rect 22385 34561 22419 34595
rect 23029 34561 23063 34595
rect 23121 34561 23155 34595
rect 23489 34561 23523 34595
rect 23765 34561 23799 34595
rect 23857 34561 23891 34595
rect 25145 34561 25179 34595
rect 25329 34561 25363 34595
rect 25421 34561 25455 34595
rect 25513 34561 25547 34595
rect 26525 34561 26559 34595
rect 26985 34561 27019 34595
rect 29101 34561 29135 34595
rect 29194 34561 29228 34595
rect 29469 34561 29503 34595
rect 29607 34561 29641 34595
rect 30849 34561 30883 34595
rect 31309 34561 31343 34595
rect 37565 34561 37599 34595
rect 4629 34493 4663 34527
rect 6101 34493 6135 34527
rect 6929 34493 6963 34527
rect 8125 34493 8159 34527
rect 16957 34493 16991 34527
rect 17969 34493 18003 34527
rect 19993 34493 20027 34527
rect 22845 34493 22879 34527
rect 23305 34493 23339 34527
rect 23397 34493 23431 34527
rect 27261 34493 27295 34527
rect 31401 34493 31435 34527
rect 31493 34493 31527 34527
rect 37841 34493 37875 34527
rect 17049 34425 17083 34459
rect 26341 34425 26375 34459
rect 6377 34357 6411 34391
rect 12817 34357 12851 34391
rect 16865 34357 16899 34391
rect 20637 34357 20671 34391
rect 21833 34357 21867 34391
rect 25697 34357 25731 34391
rect 28733 34357 28767 34391
rect 29745 34357 29779 34391
rect 30665 34357 30699 34391
rect 5365 34153 5399 34187
rect 8401 34153 8435 34187
rect 14841 34153 14875 34187
rect 16129 34153 16163 34187
rect 17417 34153 17451 34187
rect 24961 34153 24995 34187
rect 25237 34153 25271 34187
rect 26985 34153 27019 34187
rect 32781 34153 32815 34187
rect 33885 34153 33919 34187
rect 12357 34085 12391 34119
rect 32965 34085 32999 34119
rect 9965 34017 9999 34051
rect 14473 34017 14507 34051
rect 18797 34017 18831 34051
rect 24593 34017 24627 34051
rect 27445 34017 27479 34051
rect 27537 34017 27571 34051
rect 31309 34017 31343 34051
rect 33609 34017 33643 34051
rect 4445 33949 4479 33983
rect 5549 33949 5583 33983
rect 7113 33949 7147 33983
rect 8585 33949 8619 33983
rect 9689 33949 9723 33983
rect 10149 33949 10183 33983
rect 12347 33949 12381 33983
rect 12633 33949 12667 33983
rect 14749 33949 14783 33983
rect 14933 33949 14967 33983
rect 15209 33949 15243 33983
rect 16405 33949 16439 33983
rect 16497 33949 16531 33983
rect 16589 33949 16623 33983
rect 16773 33949 16807 33983
rect 17233 33949 17267 33983
rect 17693 33949 17727 33983
rect 18061 33949 18095 33983
rect 18521 33949 18555 33983
rect 18613 33949 18647 33983
rect 20361 33949 20395 33983
rect 20637 33949 20671 33983
rect 20729 33949 20763 33983
rect 25421 33949 25455 33983
rect 25513 33949 25547 33983
rect 25697 33949 25731 33983
rect 25789 33949 25823 33983
rect 28273 33949 28307 33983
rect 30021 33949 30055 33983
rect 30297 33949 30331 33983
rect 30757 33949 30791 33983
rect 30849 33949 30883 33983
rect 31033 33949 31067 33983
rect 33793 33949 33827 33983
rect 34253 33949 34287 33983
rect 16865 33881 16899 33915
rect 17049 33881 17083 33915
rect 17877 33881 17911 33915
rect 17969 33881 18003 33915
rect 20545 33881 20579 33915
rect 29837 33881 29871 33915
rect 33425 33881 33459 33915
rect 4537 33813 4571 33847
rect 7205 33813 7239 33847
rect 9321 33813 9355 33847
rect 9781 33813 9815 33847
rect 10241 33813 10275 33847
rect 12541 33813 12575 33847
rect 15117 33813 15151 33847
rect 17141 33813 17175 33847
rect 18245 33813 18279 33847
rect 18521 33813 18555 33847
rect 20913 33813 20947 33847
rect 24961 33813 24995 33847
rect 25145 33813 25179 33847
rect 27353 33813 27387 33847
rect 28365 33813 28399 33847
rect 30205 33813 30239 33847
rect 33333 33813 33367 33847
rect 34069 33813 34103 33847
rect 14749 33609 14783 33643
rect 17049 33609 17083 33643
rect 23949 33609 23983 33643
rect 24501 33609 24535 33643
rect 34621 33609 34655 33643
rect 37381 33609 37415 33643
rect 14197 33541 14231 33575
rect 14473 33541 14507 33575
rect 16681 33541 16715 33575
rect 17417 33541 17451 33575
rect 17509 33541 17543 33575
rect 19993 33541 20027 33575
rect 22017 33541 22051 33575
rect 22109 33541 22143 33575
rect 22201 33541 22235 33575
rect 16911 33507 16945 33541
rect 4353 33473 4387 33507
rect 7021 33473 7055 33507
rect 9505 33473 9539 33507
rect 14381 33473 14415 33507
rect 14565 33473 14599 33507
rect 17141 33473 17175 33507
rect 17234 33473 17268 33507
rect 17647 33473 17681 33507
rect 18153 33473 18187 33507
rect 18337 33473 18371 33507
rect 18521 33473 18555 33507
rect 18797 33473 18831 33507
rect 19050 33473 19084 33507
rect 19717 33473 19751 33507
rect 23857 33473 23891 33507
rect 24041 33473 24075 33507
rect 24409 33473 24443 33507
rect 24593 33473 24627 33507
rect 28181 33473 28215 33507
rect 32873 33473 32907 33507
rect 37565 33473 37599 33507
rect 4629 33405 4663 33439
rect 7297 33405 7331 33439
rect 9781 33405 9815 33439
rect 11253 33405 11287 33439
rect 11621 33405 11655 33439
rect 19625 33405 19659 33439
rect 19993 33405 20027 33439
rect 28457 33405 28491 33439
rect 33149 33405 33183 33439
rect 21833 33337 21867 33371
rect 6101 33269 6135 33303
rect 8769 33269 8803 33303
rect 12173 33269 12207 33303
rect 16865 33269 16899 33303
rect 17785 33269 17819 33303
rect 19809 33269 19843 33303
rect 22385 33269 22419 33303
rect 29929 33269 29963 33303
rect 5181 33065 5215 33099
rect 7573 33065 7607 33099
rect 9781 33065 9815 33099
rect 16957 33065 16991 33099
rect 18337 33065 18371 33099
rect 27905 33065 27939 33099
rect 30297 33065 30331 33099
rect 5733 32997 5767 33031
rect 28181 32997 28215 33031
rect 32873 32997 32907 33031
rect 6377 32929 6411 32963
rect 8309 32929 8343 32963
rect 8493 32929 8527 32963
rect 10241 32929 10275 32963
rect 10517 32929 10551 32963
rect 21281 32929 21315 32963
rect 28733 32929 28767 32963
rect 33425 32929 33459 32963
rect 5365 32861 5399 32895
rect 6101 32861 6135 32895
rect 7757 32861 7791 32895
rect 8217 32861 8251 32895
rect 9965 32861 9999 32895
rect 10057 32861 10091 32895
rect 10333 32861 10367 32895
rect 10425 32861 10459 32895
rect 12377 32861 12411 32895
rect 12633 32861 12667 32895
rect 12725 32861 12759 32895
rect 18153 32861 18187 32895
rect 18429 32861 18463 32895
rect 21649 32861 21683 32895
rect 22201 32861 22235 32895
rect 22294 32861 22328 32895
rect 22666 32861 22700 32895
rect 22937 32861 22971 32895
rect 23030 32861 23064 32895
rect 23402 32861 23436 32895
rect 25789 32861 25823 32895
rect 25881 32861 25915 32895
rect 26065 32861 26099 32895
rect 26157 32861 26191 32895
rect 26617 32861 26651 32895
rect 27077 32861 27111 32895
rect 28089 32861 28123 32895
rect 28549 32861 28583 32895
rect 29929 32861 29963 32895
rect 30113 32861 30147 32895
rect 33241 32861 33275 32895
rect 33885 32861 33919 32895
rect 34713 32861 34747 32895
rect 34989 32861 35023 32895
rect 12541 32793 12575 32827
rect 16773 32793 16807 32827
rect 18061 32793 18095 32827
rect 18521 32793 18555 32827
rect 19441 32793 19475 32827
rect 21557 32793 21591 32827
rect 22477 32793 22511 32827
rect 22569 32793 22603 32827
rect 23213 32793 23247 32827
rect 23305 32793 23339 32827
rect 33333 32793 33367 32827
rect 6193 32725 6227 32759
rect 7849 32725 7883 32759
rect 12909 32725 12943 32759
rect 16957 32725 16991 32759
rect 17141 32725 17175 32759
rect 20729 32725 20763 32759
rect 21465 32725 21499 32759
rect 21833 32725 21867 32759
rect 22845 32725 22879 32759
rect 23581 32725 23615 32759
rect 25605 32725 25639 32759
rect 26433 32725 26467 32759
rect 27169 32725 27203 32759
rect 28641 32725 28675 32759
rect 33701 32725 33735 32759
rect 34805 32725 34839 32759
rect 35081 32725 35115 32759
rect 22937 32521 22971 32555
rect 26065 32521 26099 32555
rect 30297 32521 30331 32555
rect 30757 32521 30791 32555
rect 31585 32521 31619 32555
rect 20913 32453 20947 32487
rect 30021 32453 30055 32487
rect 31677 32453 31711 32487
rect 7757 32385 7791 32419
rect 10885 32385 10919 32419
rect 12265 32385 12299 32419
rect 12358 32385 12392 32419
rect 12541 32385 12575 32419
rect 12633 32385 12667 32419
rect 12771 32385 12805 32419
rect 13001 32385 13035 32419
rect 18429 32385 18463 32419
rect 18521 32385 18555 32419
rect 18705 32385 18739 32419
rect 18797 32385 18831 32419
rect 19257 32385 19291 32419
rect 20085 32385 20119 32419
rect 20637 32385 20671 32419
rect 20821 32385 20855 32419
rect 21005 32385 21039 32419
rect 21833 32385 21867 32419
rect 21981 32385 22015 32419
rect 22109 32385 22143 32419
rect 22201 32385 22235 32419
rect 22298 32385 22332 32419
rect 23213 32385 23247 32419
rect 23581 32385 23615 32419
rect 23673 32385 23707 32419
rect 23857 32385 23891 32419
rect 23949 32385 23983 32419
rect 24041 32385 24075 32419
rect 25605 32385 25639 32419
rect 25697 32385 25731 32419
rect 25789 32385 25823 32419
rect 25973 32385 26007 32419
rect 26433 32385 26467 32419
rect 26985 32385 27019 32419
rect 29653 32385 29687 32419
rect 29746 32385 29780 32419
rect 29929 32385 29963 32419
rect 30118 32385 30152 32419
rect 30573 32385 30607 32419
rect 30849 32385 30883 32419
rect 32321 32385 32355 32419
rect 32689 32385 32723 32419
rect 34621 32385 34655 32419
rect 23121 32317 23155 32351
rect 23305 32317 23339 32351
rect 23397 32317 23431 32351
rect 26525 32317 26559 32351
rect 26617 32317 26651 32351
rect 27261 32317 27295 32351
rect 29009 32317 29043 32351
rect 31861 32317 31895 32351
rect 32965 32317 32999 32351
rect 34897 32317 34931 32351
rect 36645 32317 36679 32351
rect 31217 32249 31251 32283
rect 34437 32249 34471 32283
rect 7849 32181 7883 32215
rect 10701 32181 10735 32215
rect 12909 32181 12943 32215
rect 14289 32181 14323 32215
rect 18245 32181 18279 32215
rect 20085 32181 20119 32215
rect 21189 32181 21223 32215
rect 22477 32181 22511 32215
rect 24225 32181 24259 32215
rect 25329 32181 25363 32215
rect 30389 32181 30423 32215
rect 32137 32181 32171 32215
rect 13461 31977 13495 32011
rect 18613 31977 18647 32011
rect 23305 31977 23339 32011
rect 25973 31977 26007 32011
rect 31480 31977 31514 32011
rect 34253 31977 34287 32011
rect 33425 31909 33459 31943
rect 6101 31841 6135 31875
rect 7573 31841 7607 31875
rect 20821 31841 20855 31875
rect 21741 31841 21775 31875
rect 21833 31841 21867 31875
rect 29837 31841 29871 31875
rect 31125 31841 31159 31875
rect 31217 31841 31251 31875
rect 33241 31841 33275 31875
rect 33977 31841 34011 31875
rect 3893 31773 3927 31807
rect 5825 31773 5859 31807
rect 7941 31773 7975 31807
rect 8125 31773 8159 31807
rect 9505 31773 9539 31807
rect 10057 31773 10091 31807
rect 10149 31773 10183 31807
rect 10333 31773 10367 31807
rect 13369 31773 13403 31807
rect 14381 31773 14415 31807
rect 18889 31773 18923 31807
rect 20269 31773 20303 31807
rect 21097 31773 21131 31807
rect 21649 31773 21683 31807
rect 21925 31773 21959 31807
rect 22753 31773 22787 31807
rect 23029 31773 23063 31807
rect 23121 31773 23155 31807
rect 25421 31773 25455 31807
rect 25605 31773 25639 31807
rect 25697 31773 25731 31807
rect 25789 31773 25823 31807
rect 30205 31773 30239 31807
rect 30389 31773 30423 31807
rect 30757 31773 30791 31807
rect 33885 31773 33919 31807
rect 34437 31773 34471 31807
rect 4169 31705 4203 31739
rect 10609 31705 10643 31739
rect 13185 31705 13219 31739
rect 14749 31705 14783 31739
rect 18429 31705 18463 31739
rect 18613 31705 18647 31739
rect 22937 31705 22971 31739
rect 5641 31637 5675 31671
rect 7757 31637 7791 31671
rect 8677 31637 8711 31671
rect 9597 31637 9631 31671
rect 12081 31637 12115 31671
rect 14565 31637 14599 31671
rect 14657 31637 14691 31671
rect 14933 31637 14967 31671
rect 21465 31637 21499 31671
rect 33793 31637 33827 31671
rect 4077 31433 4111 31467
rect 4905 31433 4939 31467
rect 6009 31433 6043 31467
rect 6745 31433 6779 31467
rect 6837 31433 6871 31467
rect 11529 31433 11563 31467
rect 14289 31433 14323 31467
rect 18705 31433 18739 31467
rect 20729 31433 20763 31467
rect 22569 31433 22603 31467
rect 29561 31433 29595 31467
rect 31769 31433 31803 31467
rect 7757 31365 7791 31399
rect 16681 31365 16715 31399
rect 17325 31365 17359 31399
rect 19441 31365 19475 31399
rect 22385 31365 22419 31399
rect 3985 31297 4019 31331
rect 5089 31297 5123 31331
rect 5917 31297 5951 31331
rect 7481 31297 7515 31331
rect 11897 31297 11931 31331
rect 13001 31297 13035 31331
rect 16865 31297 16899 31331
rect 17141 31297 17175 31331
rect 17417 31297 17451 31331
rect 17509 31297 17543 31331
rect 18613 31297 18647 31331
rect 19165 31297 19199 31331
rect 22201 31297 22235 31331
rect 22661 31297 22695 31331
rect 22845 31297 22879 31331
rect 22937 31297 22971 31331
rect 23029 31297 23063 31331
rect 23397 31297 23431 31331
rect 25237 31297 25271 31331
rect 25329 31297 25363 31331
rect 27905 31297 27939 31331
rect 27997 31297 28031 31331
rect 28089 31297 28123 31331
rect 28273 31297 28307 31331
rect 28917 31297 28951 31331
rect 29009 31297 29043 31331
rect 29101 31297 29135 31331
rect 29285 31297 29319 31331
rect 29377 31297 29411 31331
rect 30481 31297 30515 31331
rect 31217 31297 31251 31331
rect 31309 31297 31343 31331
rect 31401 31297 31435 31331
rect 31585 31297 31619 31331
rect 31677 31297 31711 31331
rect 32321 31297 32355 31331
rect 34805 31297 34839 31331
rect 6929 31229 6963 31263
rect 9413 31229 9447 31263
rect 9689 31229 9723 31263
rect 11989 31229 12023 31263
rect 12173 31229 12207 31263
rect 6377 31161 6411 31195
rect 30665 31161 30699 31195
rect 9229 31093 9263 31127
rect 11161 31093 11195 31127
rect 17049 31093 17083 31127
rect 17693 31093 17727 31127
rect 23213 31093 23247 31127
rect 24685 31093 24719 31127
rect 25237 31093 25271 31127
rect 25605 31093 25639 31127
rect 27629 31093 27663 31127
rect 28641 31093 28675 31127
rect 30941 31093 30975 31127
rect 32137 31093 32171 31127
rect 34897 31093 34931 31127
rect 8033 30889 8067 30923
rect 8953 30889 8987 30923
rect 10057 30889 10091 30923
rect 16497 30889 16531 30923
rect 18153 30889 18187 30923
rect 19257 30889 19291 30923
rect 10609 30821 10643 30855
rect 18797 30821 18831 30855
rect 23857 30821 23891 30855
rect 28641 30821 28675 30855
rect 9505 30753 9539 30787
rect 11161 30753 11195 30787
rect 14933 30753 14967 30787
rect 16589 30753 16623 30787
rect 25237 30753 25271 30787
rect 25881 30753 25915 30787
rect 34713 30753 34747 30787
rect 6469 30685 6503 30719
rect 7481 30685 7515 30719
rect 7849 30685 7883 30719
rect 8217 30685 8251 30719
rect 9321 30685 9355 30719
rect 10241 30685 10275 30719
rect 12449 30685 12483 30719
rect 12633 30685 12667 30719
rect 12725 30685 12759 30719
rect 12817 30685 12851 30719
rect 14841 30685 14875 30719
rect 15025 30685 15059 30719
rect 15301 30685 15335 30719
rect 16313 30685 16347 30719
rect 16681 30685 16715 30719
rect 16774 30685 16808 30719
rect 17049 30685 17083 30719
rect 17187 30685 17221 30719
rect 17601 30685 17635 30719
rect 17969 30685 18003 30719
rect 18245 30685 18279 30719
rect 18613 30685 18647 30719
rect 19257 30685 19291 30719
rect 19349 30685 19383 30719
rect 20913 30685 20947 30719
rect 21005 30685 21039 30719
rect 21189 30685 21223 30719
rect 21281 30685 21315 30719
rect 21373 30685 21407 30719
rect 21557 30685 21591 30719
rect 23121 30685 23155 30719
rect 23397 30685 23431 30719
rect 23765 30685 23799 30719
rect 23949 30685 23983 30719
rect 24041 30685 24075 30719
rect 24777 30685 24811 30719
rect 25053 30685 25087 30719
rect 25605 30685 25639 30719
rect 27077 30685 27111 30719
rect 28825 30685 28859 30719
rect 29193 30685 29227 30719
rect 32781 30685 32815 30719
rect 34345 30685 34379 30719
rect 7665 30617 7699 30651
rect 7757 30617 7791 30651
rect 10977 30617 11011 30651
rect 16129 30617 16163 30651
rect 16957 30617 16991 30651
rect 17785 30617 17819 30651
rect 17877 30617 17911 30651
rect 18429 30617 18463 30651
rect 18521 30617 18555 30651
rect 21741 30617 21775 30651
rect 23581 30617 23615 30651
rect 30941 30617 30975 30651
rect 34989 30617 35023 30651
rect 36737 30617 36771 30651
rect 6561 30549 6595 30583
rect 8769 30549 8803 30583
rect 9413 30549 9447 30583
rect 11069 30549 11103 30583
rect 13001 30549 13035 30583
rect 14565 30549 14599 30583
rect 15209 30549 15243 30583
rect 17325 30549 17359 30583
rect 19625 30549 19659 30583
rect 20729 30549 20763 30583
rect 22937 30549 22971 30583
rect 23305 30549 23339 30583
rect 27169 30549 27203 30583
rect 29285 30549 29319 30583
rect 32229 30549 32263 30583
rect 32873 30549 32907 30583
rect 34161 30549 34195 30583
rect 19257 30345 19291 30379
rect 26433 30345 26467 30379
rect 34069 30345 34103 30379
rect 8493 30277 8527 30311
rect 12541 30277 12575 30311
rect 13001 30277 13035 30311
rect 14841 30277 14875 30311
rect 15393 30277 15427 30311
rect 17969 30277 18003 30311
rect 20453 30277 20487 30311
rect 20637 30277 20671 30311
rect 21097 30277 21131 30311
rect 21281 30277 21315 30311
rect 25605 30277 25639 30311
rect 26525 30277 26559 30311
rect 29377 30277 29411 30311
rect 34437 30277 34471 30311
rect 8309 30209 8343 30243
rect 8581 30209 8615 30243
rect 8677 30209 8711 30243
rect 10057 30209 10091 30243
rect 12265 30209 12299 30243
rect 12358 30209 12392 30243
rect 12633 30209 12667 30243
rect 12771 30209 12805 30243
rect 15025 30209 15059 30243
rect 15117 30209 15151 30243
rect 15209 30209 15243 30243
rect 16957 30209 16991 30243
rect 17050 30209 17084 30243
rect 17233 30209 17267 30243
rect 17325 30209 17359 30243
rect 17463 30209 17497 30243
rect 19993 30209 20027 30243
rect 20177 30209 20211 30243
rect 20269 30209 20303 30243
rect 23397 30209 23431 30243
rect 25329 30209 25363 30243
rect 25513 30209 25547 30243
rect 25697 30209 25731 30243
rect 31217 30209 31251 30243
rect 31401 30209 31435 30243
rect 31493 30209 31527 30243
rect 32137 30209 32171 30243
rect 6377 30141 6411 30175
rect 6653 30141 6687 30175
rect 26709 30141 26743 30175
rect 26985 30141 27019 30175
rect 27261 30141 27295 30175
rect 29009 30141 29043 30175
rect 29101 30141 29135 30175
rect 32413 30141 32447 30175
rect 34529 30141 34563 30175
rect 34621 30141 34655 30175
rect 8861 30073 8895 30107
rect 14289 30073 14323 30107
rect 17601 30073 17635 30107
rect 20821 30073 20855 30107
rect 24685 30073 24719 30107
rect 8125 30005 8159 30039
rect 10149 30005 10183 30039
rect 12909 30005 12943 30039
rect 19809 30005 19843 30039
rect 20637 30005 20671 30039
rect 21281 30005 21315 30039
rect 21465 30005 21499 30039
rect 25881 30005 25915 30039
rect 26065 30005 26099 30039
rect 30849 30005 30883 30039
rect 31033 30005 31067 30039
rect 33885 30005 33919 30039
rect 12541 29801 12575 29835
rect 16865 29801 16899 29835
rect 20085 29801 20119 29835
rect 20269 29801 20303 29835
rect 20637 29801 20671 29835
rect 23949 29801 23983 29835
rect 26433 29801 26467 29835
rect 28365 29801 28399 29835
rect 30389 29801 30423 29835
rect 14933 29733 14967 29767
rect 16221 29733 16255 29767
rect 24133 29733 24167 29767
rect 33793 29733 33827 29767
rect 13829 29665 13863 29699
rect 14657 29665 14691 29699
rect 15025 29665 15059 29699
rect 28825 29665 28859 29699
rect 28917 29665 28951 29699
rect 34345 29665 34379 29699
rect 4445 29597 4479 29631
rect 5733 29597 5767 29631
rect 7573 29597 7607 29631
rect 9597 29597 9631 29631
rect 12265 29597 12299 29631
rect 12357 29597 12391 29631
rect 13553 29597 13587 29631
rect 13645 29597 13679 29631
rect 13921 29597 13955 29631
rect 14841 29597 14875 29631
rect 15117 29597 15151 29631
rect 15301 29597 15335 29631
rect 15669 29597 15703 29631
rect 15853 29597 15887 29631
rect 15945 29597 15979 29631
rect 16037 29597 16071 29631
rect 16313 29597 16347 29631
rect 16681 29597 16715 29631
rect 18199 29597 18233 29631
rect 18337 29597 18371 29631
rect 18429 29597 18463 29631
rect 18613 29597 18647 29631
rect 19901 29597 19935 29631
rect 20085 29597 20119 29631
rect 22293 29597 22327 29631
rect 22661 29597 22695 29631
rect 23765 29597 23799 29631
rect 23949 29597 23983 29631
rect 25513 29597 25547 29631
rect 25605 29597 25639 29631
rect 25789 29597 25823 29631
rect 25881 29597 25915 29631
rect 26617 29597 26651 29631
rect 29745 29597 29779 29631
rect 29838 29597 29872 29631
rect 30210 29597 30244 29631
rect 30481 29597 30515 29631
rect 30665 29597 30699 29631
rect 30757 29597 30791 29631
rect 30883 29591 30917 29625
rect 31217 29597 31251 29631
rect 34713 29597 34747 29631
rect 35173 29597 35207 29631
rect 6285 29529 6319 29563
rect 20453 29529 20487 29563
rect 20637 29529 20671 29563
rect 22477 29529 22511 29563
rect 22569 29529 22603 29563
rect 30021 29529 30055 29563
rect 30113 29529 30147 29563
rect 31125 29529 31159 29563
rect 32965 29529 32999 29563
rect 34161 29529 34195 29563
rect 4537 29461 4571 29495
rect 7665 29461 7699 29495
rect 9689 29461 9723 29495
rect 13369 29461 13403 29495
rect 16497 29461 16531 29495
rect 16589 29461 16623 29495
rect 17969 29461 18003 29495
rect 20821 29461 20855 29495
rect 22845 29461 22879 29495
rect 25329 29461 25363 29495
rect 28733 29461 28767 29495
rect 34253 29461 34287 29495
rect 34805 29461 34839 29495
rect 34989 29461 35023 29495
rect 6837 29257 6871 29291
rect 22201 29257 22235 29291
rect 29929 29257 29963 29291
rect 32597 29257 32631 29291
rect 6193 29189 6227 29223
rect 18429 29189 18463 29223
rect 28641 29189 28675 29223
rect 32505 29189 32539 29223
rect 36369 29189 36403 29223
rect 4169 29121 4203 29155
rect 6745 29121 6779 29155
rect 7481 29121 7515 29155
rect 9505 29121 9539 29155
rect 12449 29121 12483 29155
rect 13185 29121 13219 29155
rect 18246 29121 18280 29155
rect 18339 29121 18373 29155
rect 18613 29121 18647 29155
rect 18705 29121 18739 29155
rect 18820 29127 18854 29161
rect 21833 29121 21867 29155
rect 22017 29121 22051 29155
rect 22293 29121 22327 29155
rect 22477 29121 22511 29155
rect 22569 29121 22603 29155
rect 22661 29121 22695 29155
rect 23213 29121 23247 29155
rect 23489 29121 23523 29155
rect 23673 29121 23707 29155
rect 25329 29121 25363 29155
rect 25421 29121 25455 29155
rect 25513 29121 25547 29155
rect 25697 29121 25731 29155
rect 26985 29121 27019 29155
rect 31585 29121 31619 29155
rect 34345 29121 34379 29155
rect 36645 29121 36679 29155
rect 36829 29121 36863 29155
rect 7021 29053 7055 29087
rect 7757 29053 7791 29087
rect 11253 29053 11287 29087
rect 11529 29053 11563 29087
rect 12265 29053 12299 29087
rect 13001 29053 13035 29087
rect 18889 29053 18923 29087
rect 32781 29053 32815 29087
rect 34621 29053 34655 29087
rect 12633 28985 12667 29019
rect 13369 28985 13403 29019
rect 18061 28985 18095 29019
rect 19165 28985 19199 29019
rect 22845 28985 22879 29019
rect 23305 28985 23339 29019
rect 23397 28985 23431 29019
rect 25053 28985 25087 29019
rect 32137 28985 32171 29019
rect 37013 28985 37047 29019
rect 4432 28917 4466 28951
rect 6377 28917 6411 28951
rect 9229 28917 9263 28951
rect 9768 28917 9802 28951
rect 12173 28917 12207 28951
rect 18797 28917 18831 28951
rect 22937 28917 22971 28951
rect 27077 28917 27111 28951
rect 31677 28917 31711 28951
rect 4997 28713 5031 28747
rect 8769 28713 8803 28747
rect 10701 28713 10735 28747
rect 24225 28645 24259 28679
rect 13737 28577 13771 28611
rect 20361 28577 20395 28611
rect 26801 28577 26835 28611
rect 28825 28577 28859 28611
rect 1961 28509 1995 28543
rect 4261 28509 4295 28543
rect 5181 28509 5215 28543
rect 6837 28509 6871 28543
rect 8217 28509 8251 28543
rect 8401 28509 8435 28543
rect 8585 28509 8619 28543
rect 9137 28509 9171 28543
rect 10149 28509 10183 28543
rect 10425 28509 10459 28543
rect 10517 28509 10551 28543
rect 10977 28509 11011 28543
rect 11161 28509 11195 28543
rect 11253 28509 11287 28543
rect 11621 28509 11655 28543
rect 12909 28509 12943 28543
rect 17233 28509 17267 28543
rect 17693 28509 17727 28543
rect 20269 28509 20303 28543
rect 20453 28509 20487 28543
rect 20545 28509 20579 28543
rect 22845 28509 22879 28543
rect 23121 28509 23155 28543
rect 23213 28509 23247 28543
rect 23673 28509 23707 28543
rect 23857 28509 23891 28543
rect 24041 28509 24075 28543
rect 25421 28509 25455 28543
rect 25789 28509 25823 28543
rect 26249 28509 26283 28543
rect 26341 28509 26375 28543
rect 26525 28509 26559 28543
rect 26617 28509 26651 28543
rect 28733 28509 28767 28543
rect 29193 28525 29227 28559
rect 29561 28509 29595 28543
rect 31493 28509 31527 28543
rect 34161 28509 34195 28543
rect 34897 28509 34931 28543
rect 8493 28441 8527 28475
rect 10333 28441 10367 28475
rect 10793 28441 10827 28475
rect 23029 28441 23063 28475
rect 23949 28441 23983 28475
rect 25605 28441 25639 28475
rect 25697 28441 25731 28475
rect 27077 28441 27111 28475
rect 29837 28441 29871 28475
rect 31769 28441 31803 28475
rect 1777 28373 1811 28407
rect 4353 28373 4387 28407
rect 6929 28373 6963 28407
rect 9689 28373 9723 28407
rect 11713 28373 11747 28407
rect 17877 28373 17911 28407
rect 20085 28373 20119 28407
rect 23397 28373 23431 28407
rect 25973 28373 26007 28407
rect 26065 28373 26099 28407
rect 28549 28373 28583 28407
rect 29009 28373 29043 28407
rect 31309 28373 31343 28407
rect 33241 28373 33275 28407
rect 34253 28373 34287 28407
rect 34713 28373 34747 28407
rect 17693 28169 17727 28203
rect 19273 28169 19307 28203
rect 19441 28169 19475 28203
rect 20821 28169 20855 28203
rect 22017 28169 22051 28203
rect 22109 28169 22143 28203
rect 22201 28169 22235 28203
rect 27077 28169 27111 28203
rect 28733 28169 28767 28203
rect 30297 28169 30331 28203
rect 31769 28169 31803 28203
rect 32137 28169 32171 28203
rect 4445 28101 4479 28135
rect 14565 28101 14599 28135
rect 17325 28101 17359 28135
rect 19073 28101 19107 28135
rect 20453 28101 20487 28135
rect 21833 28101 21867 28135
rect 23673 28101 23707 28135
rect 29929 28101 29963 28135
rect 30021 28101 30055 28135
rect 30757 28101 30791 28135
rect 33701 28101 33735 28135
rect 34345 28101 34379 28135
rect 4169 28033 4203 28067
rect 6745 28033 6779 28067
rect 11345 28033 11379 28067
rect 11529 28033 11563 28067
rect 14381 28033 14415 28067
rect 14473 28033 14507 28067
rect 14841 28033 14875 28067
rect 15393 28033 15427 28067
rect 15577 28033 15611 28067
rect 17141 28033 17175 28067
rect 17417 28033 17451 28067
rect 17509 28033 17543 28067
rect 19717 28033 19751 28067
rect 19993 28033 20027 28067
rect 20177 28033 20211 28067
rect 20270 28033 20304 28067
rect 20545 28033 20579 28067
rect 20642 28033 20676 28067
rect 21189 28033 21223 28067
rect 21281 28033 21315 28067
rect 22385 28033 22419 28067
rect 22661 28033 22695 28067
rect 22809 28033 22843 28067
rect 22937 28033 22971 28067
rect 23029 28033 23063 28067
rect 23126 28033 23160 28067
rect 23397 28033 23431 28067
rect 23490 28033 23524 28067
rect 23765 28033 23799 28067
rect 23862 28033 23896 28067
rect 26065 28033 26099 28067
rect 26157 28033 26191 28067
rect 26249 28033 26283 28067
rect 26433 28033 26467 28067
rect 27261 28033 27295 28067
rect 29101 28033 29135 28067
rect 29193 28033 29227 28067
rect 29653 28033 29687 28067
rect 29746 28033 29780 28067
rect 30118 28033 30152 28067
rect 30573 28033 30607 28067
rect 30849 28033 30883 28067
rect 31953 28033 31987 28067
rect 32505 28033 32539 28067
rect 33609 28033 33643 28067
rect 34069 28033 34103 28067
rect 7021 27965 7055 27999
rect 11805 27965 11839 27999
rect 13277 27965 13311 27999
rect 15301 27965 15335 27999
rect 21557 27965 21591 27999
rect 25789 27965 25823 27999
rect 29285 27965 29319 27999
rect 32597 27965 32631 27999
rect 32781 27965 32815 27999
rect 33793 27965 33827 27999
rect 35817 27965 35851 27999
rect 11161 27897 11195 27931
rect 14197 27897 14231 27931
rect 14749 27897 14783 27931
rect 15209 27897 15243 27931
rect 19809 27897 19843 27931
rect 19901 27897 19935 27931
rect 33241 27897 33275 27931
rect 5917 27829 5951 27863
rect 8493 27829 8527 27863
rect 15117 27829 15151 27863
rect 19257 27829 19291 27863
rect 19533 27829 19567 27863
rect 21005 27829 21039 27863
rect 21465 27829 21499 27863
rect 23305 27829 23339 27863
rect 24041 27829 24075 27863
rect 30389 27829 30423 27863
rect 4721 27625 4755 27659
rect 7205 27625 7239 27659
rect 11621 27625 11655 27659
rect 19993 27625 20027 27659
rect 21097 27625 21131 27659
rect 27169 27625 27203 27659
rect 33701 27625 33735 27659
rect 7665 27557 7699 27591
rect 14565 27557 14599 27591
rect 15117 27557 15151 27591
rect 30573 27557 30607 27591
rect 6101 27489 6135 27523
rect 8125 27489 8159 27523
rect 8217 27489 8251 27523
rect 12265 27489 12299 27523
rect 23029 27489 23063 27523
rect 23305 27489 23339 27523
rect 23397 27489 23431 27523
rect 27721 27489 27755 27523
rect 4905 27421 4939 27455
rect 5825 27421 5859 27455
rect 7389 27421 7423 27455
rect 8033 27421 8067 27455
rect 8493 27421 8527 27455
rect 11989 27421 12023 27455
rect 13093 27421 13127 27455
rect 13369 27421 13403 27455
rect 13461 27421 13495 27455
rect 14933 27421 14967 27455
rect 15761 27421 15795 27455
rect 16037 27421 16071 27455
rect 16129 27421 16163 27455
rect 16681 27421 16715 27455
rect 16829 27421 16863 27455
rect 16957 27421 16991 27455
rect 17187 27421 17221 27455
rect 19441 27421 19475 27455
rect 19625 27421 19659 27455
rect 19717 27421 19751 27455
rect 19809 27421 19843 27455
rect 20565 27421 20599 27455
rect 20821 27421 20855 27455
rect 20913 27421 20947 27455
rect 22385 27421 22419 27455
rect 22569 27421 22603 27455
rect 23213 27421 23247 27455
rect 23489 27421 23523 27455
rect 23673 27421 23707 27455
rect 27629 27421 27663 27455
rect 30757 27421 30791 27455
rect 31033 27421 31067 27455
rect 33517 27421 33551 27455
rect 13277 27353 13311 27387
rect 15945 27353 15979 27387
rect 17049 27353 17083 27387
rect 20729 27353 20763 27387
rect 30665 27353 30699 27387
rect 31401 27353 31435 27387
rect 5457 27285 5491 27319
rect 5917 27285 5951 27319
rect 8585 27285 8619 27319
rect 12081 27285 12115 27319
rect 13645 27285 13679 27319
rect 14749 27285 14783 27319
rect 14841 27285 14875 27319
rect 16313 27285 16347 27319
rect 17325 27285 17359 27319
rect 27537 27285 27571 27319
rect 11529 27081 11563 27115
rect 16681 27081 16715 27115
rect 26433 27081 26467 27115
rect 11897 27013 11931 27047
rect 13185 27013 13219 27047
rect 17601 27013 17635 27047
rect 19073 27013 19107 27047
rect 5917 26945 5951 26979
rect 8125 26945 8159 26979
rect 10333 26945 10367 26979
rect 10977 26945 11011 26979
rect 12909 26945 12943 26979
rect 13002 26945 13036 26979
rect 13277 26945 13311 26979
rect 13374 26945 13408 26979
rect 14657 26945 14691 26979
rect 15025 26945 15059 26979
rect 15117 26945 15151 26979
rect 15485 26945 15519 26979
rect 15669 26945 15703 26979
rect 15761 26945 15795 26979
rect 15945 26945 15979 26979
rect 16865 26945 16899 26979
rect 17049 26945 17083 26979
rect 17233 26945 17267 26979
rect 17417 26945 17451 26979
rect 18153 26945 18187 26979
rect 18337 26945 18371 26979
rect 18429 26945 18463 26979
rect 18521 26945 18555 26979
rect 18797 26945 18831 26979
rect 18981 26945 19015 26979
rect 19165 26945 19199 26979
rect 25605 26945 25639 26979
rect 25789 26945 25823 26979
rect 25881 26945 25915 26979
rect 25973 26945 26007 26979
rect 26249 26945 26283 26979
rect 27629 26945 27663 26979
rect 28641 26945 28675 26979
rect 28734 26945 28768 26979
rect 28917 26945 28951 26979
rect 29009 26945 29043 26979
rect 29147 26945 29181 26979
rect 34345 26945 34379 26979
rect 34805 26945 34839 26979
rect 8401 26877 8435 26911
rect 10425 26877 10459 26911
rect 10609 26877 10643 26911
rect 11989 26877 12023 26911
rect 12173 26877 12207 26911
rect 14473 26877 14507 26911
rect 15301 26877 15335 26911
rect 17141 26877 17175 26911
rect 9965 26809 9999 26843
rect 13553 26809 13587 26843
rect 15577 26809 15611 26843
rect 18705 26809 18739 26843
rect 5733 26741 5767 26775
rect 9873 26741 9907 26775
rect 10793 26741 10827 26775
rect 14289 26741 14323 26775
rect 19349 26741 19383 26775
rect 26157 26741 26191 26775
rect 27445 26741 27479 26775
rect 29285 26741 29319 26775
rect 34161 26741 34195 26775
rect 34897 26741 34931 26775
rect 10504 26537 10538 26571
rect 11989 26537 12023 26571
rect 17877 26537 17911 26571
rect 21833 26537 21867 26571
rect 29929 26537 29963 26571
rect 33333 26537 33367 26571
rect 8953 26469 8987 26503
rect 14197 26469 14231 26503
rect 17693 26469 17727 26503
rect 30573 26469 30607 26503
rect 33149 26469 33183 26503
rect 17877 26401 17911 26435
rect 27353 26401 27387 26435
rect 33885 26401 33919 26435
rect 34713 26401 34747 26435
rect 4813 26333 4847 26367
rect 4905 26333 4939 26367
rect 5089 26333 5123 26367
rect 9137 26333 9171 26367
rect 9965 26333 9999 26367
rect 10057 26333 10091 26367
rect 10241 26333 10275 26367
rect 14105 26333 14139 26367
rect 14657 26333 14691 26367
rect 14933 26333 14967 26367
rect 16405 26333 16439 26367
rect 16589 26333 16623 26367
rect 16773 26333 16807 26367
rect 17049 26333 17083 26367
rect 17142 26333 17176 26367
rect 17325 26333 17359 26367
rect 17555 26333 17589 26367
rect 17785 26333 17819 26367
rect 20821 26333 20855 26367
rect 21005 26333 21039 26367
rect 21189 26333 21223 26367
rect 24041 26333 24075 26367
rect 24133 26333 24167 26367
rect 24409 26333 24443 26367
rect 26617 26333 26651 26367
rect 26709 26333 26743 26367
rect 26801 26333 26835 26367
rect 26985 26333 27019 26367
rect 27077 26333 27111 26367
rect 29193 26333 29227 26367
rect 30113 26333 30147 26367
rect 30297 26333 30331 26367
rect 30389 26333 30423 26367
rect 30849 26333 30883 26367
rect 30941 26333 30975 26367
rect 31033 26333 31067 26367
rect 31217 26333 31251 26367
rect 31401 26333 31435 26367
rect 34345 26333 34379 26367
rect 5365 26265 5399 26299
rect 7113 26265 7147 26299
rect 16221 26265 16255 26299
rect 17417 26265 17451 26299
rect 21089 26265 21123 26299
rect 21465 26265 21499 26299
rect 21649 26265 21683 26299
rect 24685 26265 24719 26299
rect 26341 26265 26375 26299
rect 31677 26265 31711 26299
rect 33701 26265 33735 26299
rect 34989 26265 35023 26299
rect 36737 26265 36771 26299
rect 16497 26197 16531 26231
rect 18153 26197 18187 26231
rect 21373 26197 21407 26231
rect 26157 26197 26191 26231
rect 28825 26197 28859 26231
rect 29285 26197 29319 26231
rect 33793 26197 33827 26231
rect 34437 26197 34471 26231
rect 6469 25993 6503 26027
rect 23857 25993 23891 26027
rect 24409 25993 24443 26027
rect 24501 25993 24535 26027
rect 25789 25993 25823 26027
rect 27261 25993 27295 26027
rect 27537 25993 27571 26027
rect 28825 25993 28859 26027
rect 31585 25993 31619 26027
rect 31769 25993 31803 26027
rect 32137 25993 32171 26027
rect 32597 25993 32631 26027
rect 33977 25993 34011 26027
rect 6837 25925 6871 25959
rect 13001 25925 13035 25959
rect 15761 25925 15795 25959
rect 23029 25925 23063 25959
rect 29377 25925 29411 25959
rect 32505 25925 32539 25959
rect 36369 25925 36403 25959
rect 6009 25857 6043 25891
rect 10425 25857 10459 25891
rect 11805 25857 11839 25891
rect 11897 25857 11931 25891
rect 15025 25857 15059 25891
rect 15485 25857 15519 25891
rect 18245 25857 18279 25891
rect 20637 25857 20671 25891
rect 20913 25857 20947 25891
rect 22385 25857 22419 25891
rect 22569 25857 22603 25891
rect 22661 25857 22695 25891
rect 22845 25857 22879 25891
rect 23121 25857 23155 25891
rect 23213 25857 23247 25891
rect 23673 25857 23707 25891
rect 23949 25857 23983 25891
rect 24041 25857 24075 25891
rect 24685 25857 24719 25891
rect 25973 25857 26007 25891
rect 26065 25857 26099 25891
rect 26249 25857 26283 25891
rect 26341 25857 26375 25891
rect 27169 25857 27203 25891
rect 27905 25857 27939 25891
rect 29009 25857 29043 25891
rect 31493 25857 31527 25891
rect 31953 25857 31987 25891
rect 33885 25857 33919 25891
rect 6929 25789 6963 25823
rect 7021 25789 7055 25823
rect 18337 25789 18371 25823
rect 24133 25789 24167 25823
rect 27997 25789 28031 25823
rect 28181 25789 28215 25823
rect 29101 25789 29135 25823
rect 31125 25789 31159 25823
rect 32781 25789 32815 25823
rect 34069 25789 34103 25823
rect 34345 25789 34379 25823
rect 34621 25789 34655 25823
rect 22477 25721 22511 25755
rect 5825 25653 5859 25687
rect 10241 25653 10275 25687
rect 12081 25653 12115 25687
rect 14473 25653 14507 25687
rect 18429 25653 18463 25687
rect 18613 25653 18647 25687
rect 20453 25653 20487 25687
rect 20821 25653 20855 25687
rect 22201 25653 22235 25687
rect 23397 25653 23431 25687
rect 23489 25653 23523 25687
rect 24041 25653 24075 25687
rect 33517 25653 33551 25687
rect 5536 25449 5570 25483
rect 7205 25449 7239 25483
rect 11621 25449 11655 25483
rect 20361 25449 20395 25483
rect 22661 25449 22695 25483
rect 23029 25449 23063 25483
rect 24409 25449 24443 25483
rect 25329 25449 25363 25483
rect 28365 25449 28399 25483
rect 34069 25449 34103 25483
rect 7021 25381 7055 25415
rect 11437 25381 11471 25415
rect 7757 25313 7791 25347
rect 9965 25313 9999 25347
rect 12173 25313 12207 25347
rect 12633 25313 12667 25347
rect 13737 25313 13771 25347
rect 17325 25313 17359 25347
rect 22753 25313 22787 25347
rect 24869 25313 24903 25347
rect 24961 25313 24995 25347
rect 29009 25313 29043 25347
rect 1685 25245 1719 25279
rect 4997 25245 5031 25279
rect 5089 25245 5123 25279
rect 5273 25245 5307 25279
rect 7573 25245 7607 25279
rect 8033 25245 8067 25279
rect 8585 25245 8619 25279
rect 9413 25245 9447 25279
rect 9505 25245 9539 25279
rect 9689 25245 9723 25279
rect 11989 25245 12023 25279
rect 12817 25245 12851 25279
rect 13461 25245 13495 25279
rect 13645 25245 13679 25279
rect 14197 25245 14231 25279
rect 14657 25245 14691 25279
rect 15117 25245 15151 25279
rect 16589 25245 16623 25279
rect 17233 25245 17267 25279
rect 18429 25245 18463 25279
rect 18797 25245 18831 25279
rect 18889 25245 18923 25279
rect 19809 25245 19843 25279
rect 19993 25245 20027 25279
rect 20177 25245 20211 25279
rect 20637 25245 20671 25279
rect 21005 25245 21039 25279
rect 21281 25245 21315 25279
rect 22661 25245 22695 25279
rect 25605 25245 25639 25279
rect 25697 25245 25731 25279
rect 25789 25245 25823 25279
rect 25973 25245 26007 25279
rect 26249 25245 26283 25279
rect 26341 25245 26375 25279
rect 26525 25245 26559 25279
rect 26617 25245 26651 25279
rect 28733 25245 28767 25279
rect 34253 25245 34287 25279
rect 1961 25177 1995 25211
rect 13001 25177 13035 25211
rect 18521 25177 18555 25211
rect 18613 25177 18647 25211
rect 20085 25177 20119 25211
rect 21557 25177 21591 25211
rect 26065 25177 26099 25211
rect 28825 25177 28859 25211
rect 3433 25109 3467 25143
rect 7665 25109 7699 25143
rect 8125 25109 8159 25143
rect 8401 25109 8435 25143
rect 12081 25109 12115 25143
rect 14866 25109 14900 25143
rect 18245 25109 18279 25143
rect 24777 25109 24811 25143
rect 1593 24905 1627 24939
rect 2145 24905 2179 24939
rect 9781 24905 9815 24939
rect 10149 24905 10183 24939
rect 21005 24905 21039 24939
rect 22753 24905 22787 24939
rect 28273 24905 28307 24939
rect 28457 24905 28491 24939
rect 2789 24837 2823 24871
rect 8125 24837 8159 24871
rect 20637 24837 20671 24871
rect 20729 24837 20763 24871
rect 25697 24837 25731 24871
rect 1501 24769 1535 24803
rect 2329 24769 2363 24803
rect 12173 24769 12207 24803
rect 12633 24769 12667 24803
rect 13369 24769 13403 24803
rect 13737 24769 13771 24803
rect 14381 24769 14415 24803
rect 14841 24769 14875 24803
rect 16129 24769 16163 24803
rect 16313 24769 16347 24803
rect 17049 24769 17083 24803
rect 17877 24769 17911 24803
rect 17969 24769 18003 24803
rect 18061 24769 18095 24803
rect 18245 24769 18279 24803
rect 18613 24769 18647 24803
rect 19165 24769 19199 24803
rect 20361 24769 20395 24803
rect 20509 24769 20543 24803
rect 20867 24769 20901 24803
rect 22109 24769 22143 24803
rect 22202 24769 22236 24803
rect 22385 24769 22419 24803
rect 22477 24769 22511 24803
rect 22574 24769 22608 24803
rect 25513 24769 25547 24803
rect 25789 24769 25823 24803
rect 25881 24769 25915 24803
rect 28181 24769 28215 24803
rect 28641 24769 28675 24803
rect 29377 24769 29411 24803
rect 29561 24769 29595 24803
rect 29653 24769 29687 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 32413 24769 32447 24803
rect 32597 24769 32631 24803
rect 32689 24769 32723 24803
rect 32873 24769 32907 24803
rect 34805 24769 34839 24803
rect 2881 24701 2915 24735
rect 3065 24701 3099 24735
rect 3433 24701 3467 24735
rect 3709 24701 3743 24735
rect 7849 24701 7883 24735
rect 10241 24701 10275 24735
rect 10425 24701 10459 24735
rect 12725 24701 12759 24735
rect 13277 24701 13311 24735
rect 13921 24701 13955 24735
rect 14197 24701 14231 24735
rect 15117 24701 15151 24735
rect 17325 24701 17359 24735
rect 17601 24701 17635 24735
rect 18889 24701 18923 24735
rect 19441 24701 19475 24735
rect 2421 24633 2455 24667
rect 11989 24633 12023 24667
rect 26065 24633 26099 24667
rect 32413 24633 32447 24667
rect 5181 24565 5215 24599
rect 9597 24565 9631 24599
rect 16497 24565 16531 24599
rect 29193 24565 29227 24599
rect 32229 24565 32263 24599
rect 32689 24565 32723 24599
rect 34897 24565 34931 24599
rect 3985 24361 4019 24395
rect 11253 24361 11287 24395
rect 14841 24361 14875 24395
rect 16405 24361 16439 24395
rect 17693 24361 17727 24395
rect 17877 24361 17911 24395
rect 21557 24361 21591 24395
rect 22753 24361 22787 24395
rect 26433 24361 26467 24395
rect 28273 24361 28307 24395
rect 31401 24361 31435 24395
rect 33241 24361 33275 24395
rect 4445 24293 4479 24327
rect 12633 24293 12667 24327
rect 13645 24293 13679 24327
rect 14565 24293 14599 24327
rect 19625 24293 19659 24327
rect 23489 24293 23523 24327
rect 24501 24293 24535 24327
rect 32505 24293 32539 24327
rect 4997 24225 5031 24259
rect 6469 24225 6503 24259
rect 11805 24225 11839 24259
rect 14105 24225 14139 24259
rect 14657 24225 14691 24259
rect 16865 24225 16899 24259
rect 18797 24225 18831 24259
rect 21005 24225 21039 24259
rect 25053 24225 25087 24259
rect 28733 24225 28767 24259
rect 28825 24225 28859 24259
rect 32321 24225 32355 24259
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 12541 24157 12575 24191
rect 12725 24157 12759 24191
rect 12909 24157 12943 24191
rect 13369 24157 13403 24191
rect 13645 24157 13679 24191
rect 14289 24157 14323 24191
rect 14749 24157 14783 24191
rect 15301 24157 15335 24191
rect 15761 24157 15795 24191
rect 15854 24157 15888 24191
rect 16037 24157 16071 24191
rect 16129 24157 16163 24191
rect 16226 24157 16260 24191
rect 16773 24157 16807 24191
rect 17233 24157 17267 24191
rect 18153 24157 18187 24191
rect 18245 24157 18279 24191
rect 18337 24157 18371 24191
rect 19993 24157 20027 24191
rect 20177 24157 20211 24191
rect 20269 24157 20303 24191
rect 20417 24157 20451 24191
rect 20637 24157 20671 24191
rect 20775 24157 20809 24191
rect 21189 24157 21223 24191
rect 22753 24157 22787 24191
rect 22845 24157 22879 24191
rect 24041 24157 24075 24191
rect 25789 24157 25823 24191
rect 25882 24157 25916 24191
rect 26295 24157 26329 24191
rect 26709 24157 26743 24191
rect 27077 24157 27111 24191
rect 27721 24157 27755 24191
rect 27905 24157 27939 24191
rect 28181 24157 28215 24191
rect 30297 24157 30331 24191
rect 30389 24157 30423 24191
rect 30481 24157 30515 24191
rect 30665 24157 30699 24191
rect 30757 24157 30791 24191
rect 30941 24157 30975 24191
rect 31033 24157 31067 24191
rect 31217 24157 31251 24191
rect 31309 24157 31343 24191
rect 32045 24157 32079 24191
rect 32137 24157 32171 24191
rect 32413 24157 32447 24191
rect 32505 24157 32539 24191
rect 32781 24157 32815 24191
rect 32873 24157 32907 24191
rect 33149 24157 33183 24191
rect 33977 24157 34011 24191
rect 34345 24157 34379 24191
rect 34805 24157 34839 24191
rect 34989 24157 35023 24191
rect 6745 24089 6779 24123
rect 17509 24089 17543 24123
rect 20545 24089 20579 24123
rect 23305 24089 23339 24123
rect 26065 24089 26099 24123
rect 26157 24089 26191 24123
rect 26893 24089 26927 24123
rect 26985 24089 27019 24123
rect 34161 24089 34195 24123
rect 34253 24089 34287 24123
rect 4905 24021 4939 24055
rect 8217 24021 8251 24055
rect 11621 24021 11655 24055
rect 11713 24021 11747 24055
rect 17693 24021 17727 24055
rect 19809 24021 19843 24055
rect 19901 24021 19935 24055
rect 20913 24021 20947 24055
rect 21281 24021 21315 24055
rect 21373 24021 21407 24055
rect 23121 24021 23155 24055
rect 24133 24021 24167 24055
rect 24869 24021 24903 24055
rect 24961 24021 24995 24055
rect 27261 24021 27295 24055
rect 28641 24021 28675 24055
rect 30021 24021 30055 24055
rect 30849 24021 30883 24055
rect 31217 24021 31251 24055
rect 31769 24021 31803 24055
rect 31861 24021 31895 24055
rect 32689 24021 32723 24055
rect 32965 24021 32999 24055
rect 34529 24021 34563 24055
rect 35817 24021 35851 24055
rect 6929 23817 6963 23851
rect 7205 23817 7239 23851
rect 10793 23817 10827 23851
rect 13829 23817 13863 23851
rect 14105 23817 14139 23851
rect 18429 23817 18463 23851
rect 26065 23817 26099 23851
rect 29837 23817 29871 23851
rect 31769 23817 31803 23851
rect 32413 23817 32447 23851
rect 12909 23749 12943 23783
rect 13277 23749 13311 23783
rect 24041 23749 24075 23783
rect 27169 23749 27203 23783
rect 28365 23749 28399 23783
rect 1409 23681 1443 23715
rect 7113 23681 7147 23715
rect 7573 23681 7607 23715
rect 10517 23681 10551 23715
rect 10701 23681 10735 23715
rect 10885 23681 10919 23715
rect 13093 23681 13127 23715
rect 13461 23681 13495 23715
rect 13737 23681 13771 23715
rect 13915 23681 13949 23715
rect 14013 23681 14047 23715
rect 14197 23681 14231 23715
rect 15853 23681 15887 23715
rect 16037 23681 16071 23715
rect 16129 23681 16163 23715
rect 16221 23681 16255 23715
rect 17141 23681 17175 23715
rect 17325 23681 17359 23715
rect 17509 23681 17543 23715
rect 18153 23681 18187 23715
rect 18429 23681 18463 23715
rect 18613 23681 18647 23715
rect 22293 23681 22327 23715
rect 22477 23681 22511 23715
rect 22569 23681 22603 23715
rect 22662 23681 22696 23715
rect 23029 23681 23063 23715
rect 23213 23681 23247 23715
rect 23305 23681 23339 23715
rect 23398 23681 23432 23715
rect 23673 23681 23707 23715
rect 23765 23681 23799 23715
rect 24317 23681 24351 23715
rect 26985 23681 27019 23715
rect 27261 23681 27295 23715
rect 27353 23681 27387 23715
rect 28089 23681 28123 23715
rect 31677 23681 31711 23715
rect 32321 23681 32355 23715
rect 34805 23681 34839 23715
rect 35173 23681 35207 23715
rect 35357 23681 35391 23715
rect 1685 23613 1719 23647
rect 7665 23613 7699 23647
rect 7757 23613 7791 23647
rect 13553 23613 13587 23647
rect 19441 23613 19475 23647
rect 24593 23613 24627 23647
rect 34989 23613 35023 23647
rect 35081 23613 35115 23647
rect 16957 23545 16991 23579
rect 22937 23545 22971 23579
rect 27537 23545 27571 23579
rect 35173 23545 35207 23579
rect 3157 23477 3191 23511
rect 10333 23477 10367 23511
rect 16405 23477 16439 23511
rect 34621 23477 34655 23511
rect 1777 23273 1811 23307
rect 3801 23273 3835 23307
rect 8033 23273 8067 23307
rect 15393 23273 15427 23307
rect 17693 23273 17727 23307
rect 17877 23273 17911 23307
rect 24685 23273 24719 23307
rect 27353 23273 27387 23307
rect 13829 23205 13863 23239
rect 16313 23205 16347 23239
rect 25789 23205 25823 23239
rect 2973 23137 3007 23171
rect 4813 23137 4847 23171
rect 7205 23137 7239 23171
rect 10149 23137 10183 23171
rect 14841 23137 14875 23171
rect 17049 23137 17083 23171
rect 19257 23137 19291 23171
rect 22201 23137 22235 23171
rect 22477 23137 22511 23171
rect 22845 23137 22879 23171
rect 23489 23137 23523 23171
rect 36093 23137 36127 23171
rect 1961 23069 1995 23103
rect 2697 23069 2731 23103
rect 3985 23069 4019 23103
rect 4169 23069 4203 23103
rect 4445 23069 4479 23103
rect 8217 23069 8251 23103
rect 8401 23069 8435 23103
rect 8519 23069 8553 23103
rect 8677 23069 8711 23103
rect 9597 23069 9631 23103
rect 9689 23069 9723 23103
rect 9873 23069 9907 23103
rect 13369 23069 13403 23103
rect 13553 23069 13587 23103
rect 13921 23069 13955 23103
rect 14105 23069 14139 23103
rect 14933 23069 14967 23103
rect 16221 23069 16255 23103
rect 16773 23069 16807 23103
rect 17969 23069 18003 23103
rect 18613 23069 18647 23103
rect 18797 23069 18831 23103
rect 19533 23069 19567 23103
rect 21741 23069 21775 23103
rect 22109 23069 22143 23103
rect 22937 23069 22971 23103
rect 23305 23069 23339 23103
rect 24869 23069 24903 23103
rect 25237 23069 25271 23103
rect 25421 23069 25455 23103
rect 25610 23069 25644 23103
rect 31759 23069 31793 23103
rect 31953 23069 31987 23103
rect 35265 23069 35299 23103
rect 35449 23069 35483 23103
rect 35725 23069 35759 23103
rect 36001 23069 36035 23103
rect 36277 23069 36311 23103
rect 36461 23069 36495 23103
rect 37565 23069 37599 23103
rect 4077 23001 4111 23035
rect 4307 23001 4341 23035
rect 5089 23001 5123 23035
rect 7021 23001 7055 23035
rect 8309 23001 8343 23035
rect 8953 23001 8987 23035
rect 9137 23001 9171 23035
rect 11897 23001 11931 23035
rect 17509 23001 17543 23035
rect 17725 23001 17759 23035
rect 19625 23001 19659 23035
rect 19993 23001 20027 23035
rect 21833 23001 21867 23035
rect 25513 23001 25547 23035
rect 27077 23001 27111 23035
rect 35541 23001 35575 23035
rect 36369 23001 36403 23035
rect 2329 22933 2363 22967
rect 2789 22933 2823 22967
rect 6561 22933 6595 22967
rect 6653 22933 6687 22967
rect 7113 22933 7147 22967
rect 9321 22933 9355 22967
rect 18061 22933 18095 22967
rect 19441 22933 19475 22967
rect 21465 22933 21499 22967
rect 21925 22933 21959 22967
rect 31953 22933 31987 22967
rect 35357 22933 35391 22967
rect 35909 22933 35943 22967
rect 37381 22933 37415 22967
rect 2145 22729 2179 22763
rect 3341 22729 3375 22763
rect 4445 22729 4479 22763
rect 5365 22729 5399 22763
rect 8309 22729 8343 22763
rect 10057 22729 10091 22763
rect 11529 22729 11563 22763
rect 11897 22729 11931 22763
rect 21281 22729 21315 22763
rect 22201 22729 22235 22763
rect 34621 22729 34655 22763
rect 3157 22661 3191 22695
rect 3709 22661 3743 22695
rect 4261 22661 4295 22695
rect 4537 22661 4571 22695
rect 7021 22661 7055 22695
rect 10517 22661 10551 22695
rect 14013 22661 14047 22695
rect 16221 22661 16255 22695
rect 22293 22661 22327 22695
rect 27169 22661 27203 22695
rect 28825 22661 28859 22695
rect 34437 22661 34471 22695
rect 4767 22627 4801 22661
rect 2421 22593 2455 22627
rect 2513 22593 2547 22627
rect 2605 22593 2639 22627
rect 2789 22593 2823 22627
rect 3065 22593 3099 22627
rect 3249 22593 3283 22627
rect 3525 22593 3559 22627
rect 3617 22593 3651 22627
rect 3847 22593 3881 22627
rect 3985 22593 4019 22627
rect 4077 22593 4111 22627
rect 4997 22593 5031 22627
rect 5549 22593 5583 22627
rect 6653 22593 6687 22627
rect 6837 22593 6871 22627
rect 6929 22593 6963 22627
rect 7139 22593 7173 22627
rect 7592 22593 7626 22627
rect 7757 22593 7791 22627
rect 7849 22593 7883 22627
rect 8217 22593 8251 22627
rect 8401 22593 8435 22627
rect 10425 22593 10459 22627
rect 14289 22593 14323 22627
rect 15025 22593 15059 22627
rect 15209 22593 15243 22627
rect 15485 22593 15519 22627
rect 17325 22593 17359 22627
rect 17693 22593 17727 22627
rect 18429 22593 18463 22627
rect 18981 22593 19015 22627
rect 19073 22593 19107 22627
rect 20453 22593 20487 22627
rect 20545 22593 20579 22627
rect 20729 22593 20763 22627
rect 21097 22593 21131 22627
rect 21189 22593 21223 22627
rect 22109 22593 22143 22627
rect 26985 22593 27019 22627
rect 27261 22593 27295 22627
rect 27353 22593 27387 22627
rect 28733 22593 28767 22627
rect 28917 22593 28951 22627
rect 29009 22593 29043 22627
rect 29285 22593 29319 22627
rect 29469 22593 29503 22627
rect 31217 22593 31251 22627
rect 31401 22593 31435 22627
rect 31677 22593 31711 22627
rect 31861 22593 31895 22627
rect 31953 22593 31987 22627
rect 32321 22593 32355 22627
rect 32413 22593 32447 22627
rect 32597 22593 32631 22627
rect 32689 22593 32723 22627
rect 34161 22593 34195 22627
rect 34345 22593 34379 22627
rect 34713 22593 34747 22627
rect 35633 22593 35667 22627
rect 35725 22593 35759 22627
rect 37657 22593 37691 22627
rect 7297 22525 7331 22559
rect 10701 22525 10735 22559
rect 11989 22525 12023 22559
rect 12173 22525 12207 22559
rect 14105 22525 14139 22559
rect 16865 22525 16899 22559
rect 17141 22525 17175 22559
rect 17601 22525 17635 22559
rect 21557 22525 21591 22559
rect 22569 22525 22603 22559
rect 5089 22457 5123 22491
rect 7389 22457 7423 22491
rect 14473 22457 14507 22491
rect 15209 22457 15243 22491
rect 18337 22457 18371 22491
rect 20269 22457 20303 22491
rect 31309 22457 31343 22491
rect 37841 22457 37875 22491
rect 4721 22389 4755 22423
rect 4905 22389 4939 22423
rect 14289 22389 14323 22423
rect 19993 22389 20027 22423
rect 20361 22389 20395 22423
rect 20821 22389 20855 22423
rect 21465 22389 21499 22423
rect 21833 22389 21867 22423
rect 22477 22389 22511 22423
rect 27537 22389 27571 22423
rect 29101 22389 29135 22423
rect 29285 22389 29319 22423
rect 31493 22389 31527 22423
rect 32137 22389 32171 22423
rect 34253 22389 34287 22423
rect 34437 22389 34471 22423
rect 35909 22389 35943 22423
rect 3801 22185 3835 22219
rect 7205 22185 7239 22219
rect 10885 22185 10919 22219
rect 20637 22185 20671 22219
rect 20913 22185 20947 22219
rect 21005 22185 21039 22219
rect 21097 22185 21131 22219
rect 29193 22185 29227 22219
rect 31401 22185 31435 22219
rect 7573 22117 7607 22151
rect 16589 22117 16623 22151
rect 18153 22117 18187 22151
rect 24409 22117 24443 22151
rect 25697 22117 25731 22151
rect 28089 22117 28123 22151
rect 31677 22117 31711 22151
rect 32045 22117 32079 22151
rect 4077 22049 4111 22083
rect 5273 22049 5307 22083
rect 5917 22049 5951 22083
rect 8125 22049 8159 22083
rect 9321 22049 9355 22083
rect 11529 22049 11563 22083
rect 15853 22049 15887 22083
rect 16129 22049 16163 22083
rect 18797 22049 18831 22083
rect 22661 22049 22695 22083
rect 26893 22049 26927 22083
rect 28825 22049 28859 22083
rect 30573 22049 30607 22083
rect 33701 22049 33735 22083
rect 34437 22049 34471 22083
rect 35265 22049 35299 22083
rect 35541 22049 35575 22083
rect 3985 21981 4019 22015
rect 4169 21981 4203 22015
rect 4261 21981 4295 22015
rect 4813 21981 4847 22015
rect 5457 21981 5491 22015
rect 5641 21981 5675 22015
rect 5759 21981 5793 22015
rect 7481 21981 7515 22015
rect 7941 21981 7975 22015
rect 9137 21981 9171 22015
rect 12541 21981 12575 22015
rect 12633 21981 12667 22015
rect 12725 21981 12759 22015
rect 12909 21981 12943 22015
rect 15117 21981 15151 22015
rect 15301 21981 15335 22015
rect 16497 21981 16531 22015
rect 16865 21981 16899 22015
rect 17141 21981 17175 22015
rect 18061 21981 18095 22015
rect 18337 21981 18371 22015
rect 21189 21981 21223 22015
rect 21373 21981 21407 22015
rect 21557 21981 21591 22015
rect 22017 21981 22051 22015
rect 22201 21981 22235 22015
rect 22293 21981 22327 22015
rect 7251 21947 7285 21981
rect 22386 21959 22420 21993
rect 24685 21981 24719 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 25053 21981 25087 22015
rect 25145 21981 25179 22015
rect 25421 21981 25455 22015
rect 25513 21981 25547 22015
rect 27077 21981 27111 22015
rect 27537 21981 27571 22015
rect 27905 21981 27939 22015
rect 28181 21981 28215 22015
rect 28549 21981 28583 22015
rect 29009 21981 29043 22015
rect 29561 21981 29595 22015
rect 29745 21981 29779 22015
rect 29837 21981 29871 22015
rect 30389 21981 30423 22015
rect 31033 21981 31067 22015
rect 31217 21981 31251 22015
rect 31585 21981 31619 22015
rect 31769 21981 31803 22015
rect 31861 21981 31895 22015
rect 32045 21981 32079 22015
rect 32229 21981 32263 22015
rect 32321 21981 32355 22015
rect 32689 21981 32723 22015
rect 32781 21981 32815 22015
rect 32873 21981 32907 22015
rect 33057 21981 33091 22015
rect 34161 21981 34195 22015
rect 34253 21981 34287 22015
rect 34345 21981 34379 22015
rect 36001 21981 36035 22015
rect 4629 21913 4663 21947
rect 5549 21913 5583 21947
rect 6009 21913 6043 21947
rect 6193 21913 6227 21947
rect 7021 21913 7055 21947
rect 7757 21913 7791 21947
rect 8953 21913 8987 21947
rect 11253 21913 11287 21947
rect 25329 21913 25363 21947
rect 27721 21913 27755 21947
rect 27813 21913 27847 21947
rect 28365 21913 28399 21947
rect 28457 21913 28491 21947
rect 33517 21913 33551 21947
rect 35909 21913 35943 21947
rect 4997 21845 5031 21879
rect 6377 21845 6411 21879
rect 7389 21845 7423 21879
rect 11345 21845 11379 21879
rect 12265 21845 12299 21879
rect 21741 21845 21775 21879
rect 27261 21845 27295 21879
rect 28733 21845 28767 21879
rect 29659 21845 29693 21879
rect 30021 21845 30055 21879
rect 30481 21845 30515 21879
rect 31217 21845 31251 21879
rect 32413 21845 32447 21879
rect 33149 21845 33183 21879
rect 33609 21845 33643 21879
rect 33977 21845 34011 21879
rect 34713 21845 34747 21879
rect 35081 21845 35115 21879
rect 35173 21845 35207 21879
rect 35817 21845 35851 21879
rect 2421 21641 2455 21675
rect 9597 21641 9631 21675
rect 10241 21641 10275 21675
rect 13369 21641 13403 21675
rect 15025 21641 15059 21675
rect 16865 21641 16899 21675
rect 18981 21641 19015 21675
rect 20821 21641 20855 21675
rect 26157 21641 26191 21675
rect 27905 21641 27939 21675
rect 30205 21641 30239 21675
rect 31401 21641 31435 21675
rect 32873 21641 32907 21675
rect 34805 21641 34839 21675
rect 5365 21573 5399 21607
rect 12817 21573 12851 21607
rect 14841 21573 14875 21607
rect 16405 21573 16439 21607
rect 18521 21573 18555 21607
rect 21925 21573 21959 21607
rect 22293 21573 22327 21607
rect 27537 21573 27571 21607
rect 2237 21505 2271 21539
rect 2421 21505 2455 21539
rect 2881 21505 2915 21539
rect 5181 21505 5215 21539
rect 5641 21505 5675 21539
rect 5825 21505 5859 21539
rect 9045 21505 9079 21539
rect 9229 21505 9263 21539
rect 9321 21505 9355 21539
rect 9413 21505 9447 21539
rect 9689 21505 9723 21539
rect 9873 21505 9907 21539
rect 9965 21505 9999 21539
rect 10057 21505 10091 21539
rect 13369 21505 13403 21539
rect 14657 21505 14691 21539
rect 16037 21505 16071 21539
rect 16221 21505 16255 21539
rect 16681 21505 16715 21539
rect 16865 21505 16899 21539
rect 17417 21505 17451 21539
rect 17877 21505 17911 21539
rect 17969 21505 18003 21539
rect 19349 21505 19383 21539
rect 19717 21505 19751 21539
rect 21097 21505 21131 21539
rect 22201 21505 22235 21539
rect 22937 21505 22971 21539
rect 23029 21505 23063 21539
rect 23121 21505 23155 21539
rect 23305 21505 23339 21539
rect 25053 21505 25087 21539
rect 25697 21505 25731 21539
rect 25881 21505 25915 21539
rect 25973 21505 26007 21539
rect 26065 21505 26099 21539
rect 27353 21505 27387 21539
rect 27629 21505 27663 21539
rect 27721 21505 27755 21539
rect 29009 21505 29043 21539
rect 29193 21505 29227 21539
rect 29653 21505 29687 21539
rect 30113 21505 30147 21539
rect 30297 21505 30331 21539
rect 31585 21505 31619 21539
rect 31677 21505 31711 21539
rect 31861 21505 31895 21539
rect 32321 21505 32355 21539
rect 32413 21505 32447 21539
rect 32597 21505 32631 21539
rect 32781 21505 32815 21539
rect 32965 21505 32999 21539
rect 33885 21505 33919 21539
rect 34069 21505 34103 21539
rect 34161 21505 34195 21539
rect 34287 21505 34321 21539
rect 34713 21505 34747 21539
rect 2973 21437 3007 21471
rect 3065 21437 3099 21471
rect 13461 21437 13495 21471
rect 17325 21437 17359 21471
rect 19165 21437 19199 21471
rect 19625 21437 19659 21471
rect 21005 21437 21039 21471
rect 21189 21437 21223 21471
rect 21281 21437 21315 21471
rect 22109 21437 22143 21471
rect 24869 21437 24903 21471
rect 29745 21437 29779 21471
rect 31769 21437 31803 21471
rect 32505 21437 32539 21471
rect 21925 21369 21959 21403
rect 25789 21369 25823 21403
rect 32137 21369 32171 21403
rect 34529 21369 34563 21403
rect 2513 21301 2547 21335
rect 5549 21301 5583 21335
rect 5733 21301 5767 21335
rect 22661 21301 22695 21335
rect 25237 21301 25271 21335
rect 29009 21301 29043 21335
rect 30021 21301 30055 21335
rect 4169 21097 4203 21131
rect 10149 21097 10183 21131
rect 10793 21097 10827 21131
rect 12817 21097 12851 21131
rect 14749 21097 14783 21131
rect 16497 21097 16531 21131
rect 17325 21097 17359 21131
rect 17601 21097 17635 21131
rect 18153 21097 18187 21131
rect 23765 21097 23799 21131
rect 27261 21097 27295 21131
rect 34713 21097 34747 21131
rect 22017 21029 22051 21063
rect 1409 20961 1443 20995
rect 3157 20961 3191 20995
rect 3801 20961 3835 20995
rect 19257 20961 19291 20995
rect 19533 20961 19567 20995
rect 19993 20961 20027 20995
rect 23949 20961 23983 20995
rect 25053 20961 25087 20995
rect 25421 20961 25455 20995
rect 30205 20961 30239 20995
rect 32413 20961 32447 20995
rect 34989 20961 35023 20995
rect 35081 20961 35115 20995
rect 35633 20961 35667 20995
rect 3985 20893 4019 20927
rect 4261 20893 4295 20927
rect 5549 20893 5583 20927
rect 5641 20893 5675 20927
rect 5733 20893 5767 20927
rect 5917 20893 5951 20927
rect 9597 20893 9631 20927
rect 9781 20893 9815 20927
rect 9965 20893 9999 20927
rect 10241 20893 10275 20927
rect 10425 20893 10459 20927
rect 10609 20893 10643 20927
rect 12265 20893 12299 20927
rect 12541 20893 12575 20927
rect 12685 20893 12719 20927
rect 14105 20893 14139 20927
rect 14253 20893 14287 20927
rect 14381 20893 14415 20927
rect 14611 20893 14645 20927
rect 14933 20893 14967 20927
rect 15117 20893 15151 20927
rect 15393 20893 15427 20927
rect 16313 20893 16347 20927
rect 16773 20893 16807 20927
rect 17233 20893 17267 20927
rect 17417 20893 17451 20927
rect 17783 20893 17817 20927
rect 18245 20893 18279 20927
rect 18337 20893 18371 20927
rect 18430 20893 18464 20927
rect 18705 20893 18739 20927
rect 18843 20893 18877 20927
rect 19717 20893 19751 20927
rect 20085 20893 20119 20927
rect 20821 20893 20855 20927
rect 21005 20893 21039 20927
rect 21373 20893 21407 20927
rect 21741 20893 21775 20927
rect 24041 20893 24075 20927
rect 24409 20893 24443 20927
rect 24777 20893 24811 20927
rect 25237 20893 25271 20927
rect 26709 20893 26743 20927
rect 26893 20893 26927 20927
rect 27077 20893 27111 20927
rect 29837 20893 29871 20927
rect 30021 20893 30055 20927
rect 32321 20893 32355 20927
rect 34897 20893 34931 20927
rect 35173 20893 35207 20927
rect 35541 20893 35575 20927
rect 37381 20893 37415 20927
rect 1685 20825 1719 20859
rect 9873 20825 9907 20859
rect 10517 20825 10551 20859
rect 12449 20825 12483 20859
rect 14473 20825 14507 20859
rect 18613 20825 18647 20859
rect 19441 20825 19475 20859
rect 23765 20825 23799 20859
rect 24593 20825 24627 20859
rect 24685 20825 24719 20859
rect 26985 20825 27019 20859
rect 37565 20825 37599 20859
rect 4353 20757 4387 20791
rect 5273 20757 5307 20791
rect 15301 20757 15335 20791
rect 16681 20757 16715 20791
rect 17785 20757 17819 20791
rect 18981 20757 19015 20791
rect 24225 20757 24259 20791
rect 24961 20757 24995 20791
rect 32689 20757 32723 20791
rect 37197 20757 37231 20791
rect 37841 20757 37875 20791
rect 1593 20553 1627 20587
rect 2329 20553 2363 20587
rect 3433 20553 3467 20587
rect 8585 20553 8619 20587
rect 9597 20553 9631 20587
rect 10885 20553 10919 20587
rect 11897 20553 11931 20587
rect 11989 20553 12023 20587
rect 14473 20553 14507 20587
rect 15301 20553 15335 20587
rect 24225 20553 24259 20587
rect 35725 20553 35759 20587
rect 1501 20485 1535 20519
rect 3801 20485 3835 20519
rect 3939 20485 3973 20519
rect 9873 20485 9907 20519
rect 14933 20485 14967 20519
rect 15025 20485 15059 20519
rect 16865 20485 16899 20519
rect 22937 20485 22971 20519
rect 25329 20485 25363 20519
rect 2237 20417 2271 20451
rect 2513 20417 2547 20451
rect 2697 20417 2731 20451
rect 3617 20417 3651 20451
rect 3709 20417 3743 20451
rect 4077 20417 4111 20451
rect 4169 20417 4203 20451
rect 4353 20417 4387 20451
rect 9045 20417 9079 20451
rect 9229 20417 9263 20451
rect 9321 20417 9355 20451
rect 9413 20417 9447 20451
rect 9689 20417 9723 20451
rect 9965 20417 9999 20451
rect 10057 20417 10091 20451
rect 10333 20417 10367 20451
rect 10517 20417 10551 20451
rect 10609 20417 10643 20451
rect 10701 20417 10735 20451
rect 11805 20417 11839 20451
rect 12173 20417 12207 20451
rect 12633 20417 12667 20451
rect 12725 20417 12759 20451
rect 12909 20417 12943 20451
rect 13829 20417 13863 20451
rect 13977 20417 14011 20451
rect 14105 20417 14139 20451
rect 14197 20417 14231 20451
rect 14335 20417 14369 20451
rect 14657 20417 14691 20451
rect 14805 20417 14839 20451
rect 15122 20417 15156 20451
rect 16681 20417 16715 20451
rect 20085 20417 20119 20451
rect 20269 20417 20303 20451
rect 20361 20417 20395 20451
rect 20729 20417 20763 20451
rect 20821 20417 20855 20451
rect 21281 20417 21315 20451
rect 23213 20417 23247 20451
rect 24133 20417 24167 20451
rect 25145 20417 25179 20451
rect 25421 20417 25455 20451
rect 25513 20417 25547 20451
rect 28825 20417 28859 20451
rect 28917 20417 28951 20451
rect 29101 20417 29135 20451
rect 29193 20417 29227 20451
rect 29653 20417 29687 20451
rect 29837 20417 29871 20451
rect 35173 20417 35207 20451
rect 35909 20417 35943 20451
rect 36001 20417 36035 20451
rect 36185 20417 36219 20451
rect 36277 20417 36311 20451
rect 3249 20349 3283 20383
rect 6837 20349 6871 20383
rect 7113 20349 7147 20383
rect 17049 20349 17083 20383
rect 19901 20349 19935 20383
rect 23121 20349 23155 20383
rect 29929 20349 29963 20383
rect 35265 20349 35299 20383
rect 35449 20349 35483 20383
rect 4537 20281 4571 20315
rect 10241 20281 10275 20315
rect 11621 20281 11655 20315
rect 23397 20281 23431 20315
rect 34805 20281 34839 20315
rect 2053 20213 2087 20247
rect 20545 20213 20579 20247
rect 23213 20213 23247 20247
rect 25697 20213 25731 20247
rect 28641 20213 28675 20247
rect 29469 20213 29503 20247
rect 7389 20009 7423 20043
rect 14657 20009 14691 20043
rect 16129 20009 16163 20043
rect 17877 20009 17911 20043
rect 18429 20009 18463 20043
rect 18981 20009 19015 20043
rect 20821 20009 20855 20043
rect 21465 20009 21499 20043
rect 24409 20009 24443 20043
rect 26709 20009 26743 20043
rect 28457 20009 28491 20043
rect 35173 20009 35207 20043
rect 11989 19941 12023 19975
rect 14381 19941 14415 19975
rect 15393 19941 15427 19975
rect 24777 19941 24811 19975
rect 27813 19941 27847 19975
rect 34069 19941 34103 19975
rect 34437 19941 34471 19975
rect 34989 19941 35023 19975
rect 3341 19873 3375 19907
rect 5733 19873 5767 19907
rect 8309 19873 8343 19907
rect 11713 19873 11747 19907
rect 12357 19873 12391 19907
rect 14841 19873 14875 19907
rect 15301 19873 15335 19907
rect 20545 19873 20579 19907
rect 27261 19873 27295 19907
rect 28825 19873 28859 19907
rect 3065 19805 3099 19839
rect 4077 19805 4111 19839
rect 5641 19805 5675 19839
rect 7573 19805 7607 19839
rect 8217 19805 8251 19839
rect 12541 19805 12575 19839
rect 14289 19805 14323 19839
rect 14473 19805 14507 19839
rect 14933 19805 14967 19839
rect 15669 19805 15703 19839
rect 15761 19805 15795 19839
rect 15853 19805 15887 19839
rect 16037 19805 16071 19839
rect 16129 19805 16163 19839
rect 16313 19805 16347 19839
rect 17325 19805 17359 19839
rect 17601 19805 17635 19839
rect 17721 19805 17755 19839
rect 18554 19805 18588 19839
rect 19073 19805 19107 19839
rect 20637 19805 20671 19839
rect 22753 19805 22787 19839
rect 23857 19805 23891 19839
rect 24041 19805 24075 19839
rect 24593 19805 24627 19839
rect 24685 19805 24719 19839
rect 24869 19805 24903 19839
rect 25513 19805 25547 19839
rect 25881 19805 25915 19839
rect 26802 19805 26836 19839
rect 27169 19805 27203 19839
rect 27813 19805 27847 19839
rect 27997 19805 28031 19839
rect 28089 19805 28123 19839
rect 28365 19805 28399 19839
rect 28549 19805 28583 19839
rect 28917 19805 28951 19839
rect 29561 19805 29595 19839
rect 29929 19805 29963 19839
rect 30113 19805 30147 19839
rect 33149 19805 33183 19839
rect 33333 19805 33367 19839
rect 33793 19805 33827 19839
rect 34345 19805 34379 19839
rect 34529 19805 34563 19839
rect 34897 19805 34931 19839
rect 35081 19805 35115 19839
rect 35173 19805 35207 19839
rect 35357 19805 35391 19839
rect 15209 19737 15243 19771
rect 17509 19737 17543 19771
rect 21189 19737 21223 19771
rect 23581 19737 23615 19771
rect 25697 19737 25731 19771
rect 25789 19737 25823 19771
rect 30297 19737 30331 19771
rect 30389 19737 30423 19771
rect 2697 19669 2731 19703
rect 3157 19669 3191 19703
rect 3893 19669 3927 19703
rect 6009 19669 6043 19703
rect 7757 19669 7791 19703
rect 8125 19669 8159 19703
rect 12173 19669 12207 19703
rect 12725 19669 12759 19703
rect 18613 19669 18647 19703
rect 20177 19669 20211 19703
rect 23949 19669 23983 19703
rect 26065 19669 26099 19703
rect 28181 19669 28215 19703
rect 29285 19669 29319 19703
rect 33241 19669 33275 19703
rect 34253 19669 34287 19703
rect 9321 19465 9355 19499
rect 10793 19465 10827 19499
rect 24317 19465 24351 19499
rect 25881 19465 25915 19499
rect 26617 19465 26651 19499
rect 27445 19465 27479 19499
rect 34437 19465 34471 19499
rect 6561 19397 6595 19431
rect 6653 19397 6687 19431
rect 17601 19397 17635 19431
rect 24501 19397 24535 19431
rect 26249 19397 26283 19431
rect 31677 19397 31711 19431
rect 33977 19397 34011 19431
rect 1961 19329 1995 19363
rect 2237 19329 2271 19363
rect 4261 19329 4295 19363
rect 6377 19329 6411 19363
rect 6745 19329 6779 19363
rect 7665 19329 7699 19363
rect 9137 19329 9171 19363
rect 10425 19329 10459 19363
rect 13369 19329 13403 19363
rect 13553 19329 13587 19363
rect 16865 19329 16899 19363
rect 18705 19329 18739 19363
rect 18889 19329 18923 19363
rect 19349 19329 19383 19363
rect 19717 19329 19751 19363
rect 20545 19329 20579 19363
rect 20729 19329 20763 19363
rect 21005 19329 21039 19363
rect 22201 19329 22235 19363
rect 22477 19329 22511 19363
rect 23029 19329 23063 19363
rect 23765 19329 23799 19363
rect 23949 19329 23983 19363
rect 24041 19329 24075 19363
rect 24133 19329 24167 19363
rect 24409 19329 24443 19363
rect 24593 19329 24627 19363
rect 25697 19329 25731 19363
rect 25881 19329 25915 19363
rect 26065 19329 26099 19363
rect 26341 19329 26375 19363
rect 26433 19329 26467 19363
rect 27169 19329 27203 19363
rect 27353 19329 27387 19363
rect 28089 19329 28123 19363
rect 28273 19329 28307 19363
rect 28549 19329 28583 19363
rect 28824 19329 28858 19363
rect 29009 19329 29043 19363
rect 29101 19329 29135 19363
rect 29469 19329 29503 19363
rect 30021 19329 30055 19363
rect 30389 19329 30423 19363
rect 30481 19329 30515 19363
rect 31125 19329 31159 19363
rect 31585 19329 31619 19363
rect 32137 19329 32171 19363
rect 32321 19329 32355 19363
rect 32597 19329 32631 19363
rect 32689 19329 32723 19363
rect 32873 19329 32907 19363
rect 32965 19329 32999 19363
rect 33885 19329 33919 19363
rect 34621 19329 34655 19363
rect 34805 19329 34839 19363
rect 34897 19329 34931 19363
rect 34989 19329 35023 19363
rect 35173 19329 35207 19363
rect 2053 19261 2087 19295
rect 4537 19261 4571 19295
rect 8953 19261 8987 19295
rect 10517 19261 10551 19295
rect 13645 19261 13679 19295
rect 18613 19261 18647 19295
rect 19901 19261 19935 19295
rect 22661 19261 22695 19295
rect 28181 19261 28215 19295
rect 28733 19261 28767 19295
rect 31033 19261 31067 19295
rect 31493 19261 31527 19295
rect 32229 19261 32263 19295
rect 17233 19193 17267 19227
rect 17785 19193 17819 19227
rect 20913 19193 20947 19227
rect 23305 19193 23339 19227
rect 28641 19193 28675 19227
rect 30849 19193 30883 19227
rect 32413 19193 32447 19227
rect 1777 19125 1811 19159
rect 2421 19125 2455 19159
rect 6009 19125 6043 19159
rect 6929 19125 6963 19159
rect 7481 19125 7515 19159
rect 13185 19125 13219 19159
rect 16957 19125 16991 19159
rect 17601 19125 17635 19159
rect 28365 19125 28399 19159
rect 29193 19125 29227 19159
rect 35081 19125 35115 19159
rect 2329 18921 2363 18955
rect 3801 18921 3835 18955
rect 4813 18921 4847 18955
rect 8677 18921 8711 18955
rect 11069 18921 11103 18955
rect 11897 18921 11931 18955
rect 12541 18921 12575 18955
rect 15301 18921 15335 18955
rect 20085 18921 20119 18955
rect 20453 18921 20487 18955
rect 20637 18921 20671 18955
rect 21925 18921 21959 18955
rect 23397 18921 23431 18955
rect 23673 18921 23707 18955
rect 23765 18921 23799 18955
rect 28733 18921 28767 18955
rect 32965 18921 32999 18955
rect 10977 18853 11011 18887
rect 26709 18853 26743 18887
rect 31861 18853 31895 18887
rect 32321 18853 32355 18887
rect 34713 18853 34747 18887
rect 35541 18853 35575 18887
rect 5917 18785 5951 18819
rect 6101 18785 6135 18819
rect 6929 18785 6963 18819
rect 11161 18785 11195 18819
rect 12173 18785 12207 18819
rect 13645 18785 13679 18819
rect 17049 18785 17083 18819
rect 19073 18785 19107 18819
rect 19809 18785 19843 18819
rect 19901 18785 19935 18819
rect 22017 18785 22051 18819
rect 22477 18785 22511 18819
rect 23305 18785 23339 18819
rect 24231 18785 24265 18819
rect 31125 18785 31159 18819
rect 35173 18785 35207 18819
rect 35357 18785 35391 18819
rect 1501 18717 1535 18751
rect 2053 18717 2087 18751
rect 2145 18717 2179 18751
rect 2513 18717 2547 18751
rect 2605 18717 2639 18751
rect 4077 18717 4111 18751
rect 4169 18717 4203 18751
rect 4261 18717 4295 18751
rect 4445 18717 4479 18751
rect 4997 18717 5031 18751
rect 10333 18717 10367 18751
rect 10517 18717 10551 18751
rect 10885 18717 10919 18751
rect 11345 18717 11379 18751
rect 11437 18717 11471 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 13450 18717 13484 18751
rect 13737 18727 13771 18761
rect 14105 18717 14139 18751
rect 15209 18717 15243 18751
rect 15393 18717 15427 18751
rect 15669 18717 15703 18751
rect 16221 18717 16255 18751
rect 16497 18717 16531 18751
rect 16865 18717 16899 18751
rect 17141 18717 17175 18751
rect 17509 18717 17543 18751
rect 18521 18717 18555 18751
rect 22201 18717 22235 18751
rect 22753 18717 22787 18751
rect 22845 18717 22879 18751
rect 22937 18717 22971 18751
rect 23121 18717 23155 18751
rect 23489 18717 23523 18751
rect 23949 18717 23983 18751
rect 24133 18717 24167 18751
rect 25329 18717 25363 18751
rect 25697 18717 25731 18751
rect 25881 18717 25915 18751
rect 26157 18717 26191 18751
rect 26525 18717 26559 18751
rect 28641 18717 28675 18751
rect 28825 18717 28859 18751
rect 31033 18717 31067 18751
rect 31217 18717 31251 18751
rect 31493 18717 31527 18751
rect 31677 18717 31711 18751
rect 31769 18717 31803 18751
rect 32045 18717 32079 18751
rect 32321 18717 32355 18751
rect 32597 18717 32631 18751
rect 32873 18717 32907 18751
rect 35817 18717 35851 18751
rect 7205 18649 7239 18683
rect 12817 18649 12851 18683
rect 13001 18649 13035 18683
rect 13277 18649 13311 18683
rect 14933 18649 14967 18683
rect 18061 18649 18095 18683
rect 18153 18649 18187 18683
rect 18613 18649 18647 18683
rect 20269 18649 20303 18683
rect 21925 18649 21959 18683
rect 23213 18649 23247 18683
rect 26341 18649 26375 18683
rect 26433 18649 26467 18683
rect 31309 18649 31343 18683
rect 35081 18649 35115 18683
rect 35541 18649 35575 18683
rect 35725 18649 35759 18683
rect 1593 18581 1627 18615
rect 2789 18581 2823 18615
rect 5457 18581 5491 18615
rect 5825 18581 5859 18615
rect 10425 18581 10459 18615
rect 10609 18581 10643 18615
rect 12081 18581 12115 18615
rect 12541 18581 12575 18615
rect 12725 18581 12759 18615
rect 13185 18581 13219 18615
rect 13829 18581 13863 18615
rect 19441 18581 19475 18615
rect 20479 18581 20513 18615
rect 22385 18581 22419 18615
rect 32505 18581 32539 18615
rect 3617 18377 3651 18411
rect 6377 18377 6411 18411
rect 9137 18377 9171 18411
rect 10701 18377 10735 18411
rect 12081 18377 12115 18411
rect 15669 18377 15703 18411
rect 16865 18377 16899 18411
rect 18705 18377 18739 18411
rect 19441 18377 19475 18411
rect 32137 18377 32171 18411
rect 32781 18377 32815 18411
rect 6929 18309 6963 18343
rect 7021 18309 7055 18343
rect 10517 18309 10551 18343
rect 11989 18309 12023 18343
rect 20545 18309 20579 18343
rect 35081 18309 35115 18343
rect 1777 18241 1811 18275
rect 2145 18241 2179 18275
rect 3249 18241 3283 18275
rect 3433 18241 3467 18275
rect 6653 18241 6687 18275
rect 7113 18241 7147 18275
rect 7849 18241 7883 18275
rect 10149 18241 10183 18275
rect 10977 18241 11011 18275
rect 11069 18241 11103 18275
rect 11182 18244 11216 18278
rect 11345 18241 11379 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 15853 18241 15887 18275
rect 16037 18241 16071 18275
rect 17049 18241 17083 18275
rect 18153 18241 18187 18275
rect 18521 18241 18555 18275
rect 19073 18241 19107 18275
rect 19257 18241 19291 18275
rect 20177 18241 20211 18275
rect 20361 18241 20395 18275
rect 28549 18241 28583 18275
rect 28917 18241 28951 18275
rect 32597 18241 32631 18275
rect 32873 18241 32907 18275
rect 34713 18241 34747 18275
rect 37565 18241 37599 18275
rect 6546 18173 6580 18207
rect 7297 18173 7331 18207
rect 10333 18173 10367 18207
rect 12173 18173 12207 18207
rect 16681 18173 16715 18207
rect 18061 18173 18095 18207
rect 28365 18173 28399 18207
rect 32505 18173 32539 18207
rect 32965 18173 32999 18207
rect 34805 18173 34839 18207
rect 10149 18105 10183 18139
rect 11621 18105 11655 18139
rect 28825 18105 28859 18139
rect 34713 18105 34747 18139
rect 1961 18037 1995 18071
rect 2329 18037 2363 18071
rect 15945 18037 15979 18071
rect 17233 18037 17267 18071
rect 18521 18037 18555 18071
rect 19073 18037 19107 18071
rect 37841 18037 37875 18071
rect 7665 17833 7699 17867
rect 10333 17833 10367 17867
rect 11437 17833 11471 17867
rect 12173 17833 12207 17867
rect 16221 17833 16255 17867
rect 20361 17833 20395 17867
rect 33333 17833 33367 17867
rect 33701 17833 33735 17867
rect 9873 17765 9907 17799
rect 11621 17765 11655 17799
rect 24961 17765 24995 17799
rect 25789 17765 25823 17799
rect 26433 17765 26467 17799
rect 29929 17765 29963 17799
rect 32781 17765 32815 17799
rect 3065 17697 3099 17731
rect 7481 17697 7515 17731
rect 8217 17697 8251 17731
rect 9229 17697 9263 17731
rect 10793 17697 10827 17731
rect 10977 17697 11011 17731
rect 14105 17697 14139 17731
rect 16681 17697 16715 17731
rect 16773 17697 16807 17731
rect 23857 17697 23891 17731
rect 24133 17697 24167 17731
rect 24501 17697 24535 17731
rect 25329 17697 25363 17731
rect 25973 17697 26007 17731
rect 26617 17697 26651 17731
rect 28365 17697 28399 17731
rect 31401 17697 31435 17731
rect 31770 17697 31804 17731
rect 33793 17697 33827 17731
rect 34253 17697 34287 17731
rect 34437 17697 34471 17731
rect 3985 17629 4019 17663
rect 4169 17629 4203 17663
rect 4445 17629 4479 17663
rect 4537 17629 4571 17663
rect 5273 17629 5307 17663
rect 8125 17629 8159 17663
rect 9597 17629 9631 17663
rect 9965 17629 9999 17663
rect 11253 17629 11287 17663
rect 11437 17629 11471 17663
rect 14381 17629 14415 17663
rect 14473 17629 14507 17663
rect 14565 17629 14599 17663
rect 14749 17629 14783 17663
rect 14933 17629 14967 17663
rect 15025 17629 15059 17663
rect 15577 17629 15611 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 16405 17629 16439 17663
rect 16497 17629 16531 17663
rect 18153 17629 18187 17663
rect 19349 17629 19383 17663
rect 20637 17629 20671 17663
rect 20729 17629 20763 17663
rect 20821 17629 20855 17663
rect 21005 17629 21039 17663
rect 22661 17629 22695 17663
rect 23765 17629 23799 17663
rect 24593 17629 24627 17663
rect 25421 17629 25455 17663
rect 26065 17629 26099 17663
rect 26709 17629 26743 17663
rect 27261 17629 27295 17663
rect 27445 17629 27479 17663
rect 27537 17629 27571 17663
rect 27997 17629 28031 17663
rect 28641 17629 28675 17663
rect 28825 17629 28859 17663
rect 29837 17629 29871 17663
rect 30021 17629 30055 17663
rect 30297 17629 30331 17663
rect 30481 17629 30515 17663
rect 31585 17629 31619 17663
rect 31677 17629 31711 17663
rect 31861 17629 31895 17663
rect 33057 17629 33091 17663
rect 33701 17629 33735 17663
rect 34161 17629 34195 17663
rect 33379 17595 33413 17629
rect 4077 17561 4111 17595
rect 4307 17561 4341 17595
rect 4629 17561 4663 17595
rect 5549 17561 5583 17595
rect 7113 17561 7147 17595
rect 7297 17561 7331 17595
rect 10701 17561 10735 17595
rect 11805 17561 11839 17595
rect 11989 17561 12023 17595
rect 19533 17561 19567 17595
rect 23213 17561 23247 17595
rect 27353 17561 27387 17595
rect 32781 17561 32815 17595
rect 33149 17561 33183 17595
rect 2513 17493 2547 17527
rect 2881 17493 2915 17527
rect 2973 17493 3007 17527
rect 3801 17493 3835 17527
rect 7021 17493 7055 17527
rect 8033 17493 8067 17527
rect 14933 17493 14967 17527
rect 15393 17493 15427 17527
rect 18245 17493 18279 17527
rect 19717 17493 19751 17527
rect 27077 17493 27111 17527
rect 30389 17493 30423 17527
rect 32965 17493 32999 17527
rect 33517 17493 33551 17527
rect 34069 17493 34103 17527
rect 34437 17493 34471 17527
rect 5365 17289 5399 17323
rect 5733 17289 5767 17323
rect 10977 17289 11011 17323
rect 11253 17289 11287 17323
rect 11621 17289 11655 17323
rect 12173 17289 12207 17323
rect 13185 17289 13219 17323
rect 16221 17289 16255 17323
rect 17417 17289 17451 17323
rect 18889 17289 18923 17323
rect 20269 17289 20303 17323
rect 21005 17289 21039 17323
rect 24225 17289 24259 17323
rect 28365 17289 28399 17323
rect 29469 17289 29503 17323
rect 31585 17289 31619 17323
rect 31861 17289 31895 17323
rect 34161 17289 34195 17323
rect 34713 17289 34747 17323
rect 4537 17221 4571 17255
rect 4737 17221 4771 17255
rect 12909 17221 12943 17255
rect 13461 17221 13495 17255
rect 15945 17221 15979 17255
rect 19993 17221 20027 17255
rect 20729 17221 20763 17255
rect 29101 17221 29135 17255
rect 29301 17221 29335 17255
rect 34345 17221 34379 17255
rect 34545 17221 34579 17255
rect 35541 17221 35575 17255
rect 1409 17153 1443 17187
rect 4169 17153 4203 17187
rect 5273 17153 5307 17187
rect 9229 17153 9263 17187
rect 9413 17153 9447 17187
rect 9505 17153 9539 17187
rect 9598 17153 9632 17187
rect 10885 17153 10919 17187
rect 11069 17153 11103 17187
rect 11161 17153 11195 17187
rect 11345 17153 11379 17187
rect 11529 17153 11563 17187
rect 11713 17153 11747 17187
rect 11805 17153 11839 17187
rect 11989 17153 12023 17187
rect 12081 17153 12115 17187
rect 12265 17153 12299 17187
rect 13093 17153 13127 17187
rect 13317 17153 13351 17187
rect 14933 17153 14967 17187
rect 15577 17153 15611 17187
rect 15731 17153 15765 17187
rect 16037 17153 16071 17187
rect 16313 17153 16347 17187
rect 16865 17153 16899 17187
rect 17233 17153 17267 17187
rect 17509 17153 17543 17187
rect 17693 17153 17727 17187
rect 18613 17153 18647 17187
rect 19625 17153 19659 17187
rect 19718 17153 19752 17187
rect 19901 17153 19935 17187
rect 20090 17153 20124 17187
rect 20361 17153 20395 17187
rect 20509 17153 20543 17187
rect 20637 17153 20671 17187
rect 20867 17153 20901 17187
rect 21281 17153 21315 17187
rect 22201 17153 22235 17187
rect 22661 17153 22695 17187
rect 23213 17153 23247 17187
rect 23857 17153 23891 17187
rect 27997 17153 28031 17187
rect 28181 17153 28215 17187
rect 28273 17153 28307 17187
rect 28641 17153 28675 17187
rect 28733 17153 28767 17187
rect 28825 17153 28859 17187
rect 29009 17153 29043 17187
rect 31217 17153 31251 17187
rect 31401 17153 31435 17187
rect 31677 17153 31711 17187
rect 31953 17153 31987 17187
rect 32137 17153 32171 17187
rect 32321 17153 32355 17187
rect 33977 17153 34011 17187
rect 34253 17153 34287 17187
rect 34805 17153 34839 17187
rect 35265 17153 35299 17187
rect 1685 17085 1719 17119
rect 3893 17085 3927 17119
rect 4077 17085 4111 17119
rect 4261 17085 4295 17119
rect 4353 17085 4387 17119
rect 5825 17085 5859 17119
rect 6009 17085 6043 17119
rect 15209 17085 15243 17119
rect 16773 17085 16807 17119
rect 18245 17085 18279 17119
rect 18705 17085 18739 17119
rect 21097 17085 21131 17119
rect 21557 17085 21591 17119
rect 21925 17085 21959 17119
rect 23121 17085 23155 17119
rect 23581 17085 23615 17119
rect 23765 17085 23799 17119
rect 34897 17085 34931 17119
rect 35357 17085 35391 17119
rect 35541 17085 35575 17119
rect 4905 17017 4939 17051
rect 9873 17017 9907 17051
rect 15117 17017 15151 17051
rect 16037 17017 16071 17051
rect 22661 17017 22695 17051
rect 27997 17017 28031 17051
rect 31677 17017 31711 17051
rect 32413 17017 32447 17051
rect 35173 17017 35207 17051
rect 3157 16949 3191 16983
rect 4721 16949 4755 16983
rect 5089 16949 5123 16983
rect 11897 16949 11931 16983
rect 14749 16949 14783 16983
rect 17141 16949 17175 16983
rect 17509 16949 17543 16983
rect 21465 16949 21499 16983
rect 29285 16949 29319 16983
rect 33977 16949 34011 16983
rect 34529 16949 34563 16983
rect 34805 16949 34839 16983
rect 1961 16745 1995 16779
rect 21005 16745 21039 16779
rect 21189 16745 21223 16779
rect 35173 16745 35207 16779
rect 5825 16677 5859 16711
rect 8677 16677 8711 16711
rect 18705 16677 18739 16711
rect 22569 16677 22603 16711
rect 4629 16609 4663 16643
rect 5089 16609 5123 16643
rect 6285 16609 6319 16643
rect 6469 16609 6503 16643
rect 6929 16609 6963 16643
rect 9137 16609 9171 16643
rect 13093 16609 13127 16643
rect 14381 16609 14415 16643
rect 18061 16609 18095 16643
rect 18153 16609 18187 16643
rect 19257 16609 19291 16643
rect 20545 16609 20579 16643
rect 22825 16609 22859 16643
rect 23121 16609 23155 16643
rect 34805 16609 34839 16643
rect 2145 16541 2179 16575
rect 4721 16541 4755 16575
rect 9321 16541 9355 16575
rect 13001 16541 13035 16575
rect 14473 16541 14507 16575
rect 14749 16541 14783 16575
rect 18429 16541 18463 16575
rect 19717 16541 19751 16575
rect 19901 16541 19935 16575
rect 20085 16541 20119 16575
rect 20637 16541 20671 16575
rect 21465 16541 21499 16575
rect 31217 16541 31251 16575
rect 34897 16541 34931 16575
rect 7205 16473 7239 16507
rect 14841 16473 14875 16507
rect 17969 16473 18003 16507
rect 20821 16473 20855 16507
rect 21037 16473 21071 16507
rect 22017 16473 22051 16507
rect 22569 16473 22603 16507
rect 23029 16473 23063 16507
rect 6193 16405 6227 16439
rect 9505 16405 9539 16439
rect 12541 16405 12575 16439
rect 12909 16405 12943 16439
rect 14197 16405 14231 16439
rect 17601 16405 17635 16439
rect 18889 16405 18923 16439
rect 22937 16405 22971 16439
rect 31401 16405 31435 16439
rect 7665 16201 7699 16235
rect 8493 16201 8527 16235
rect 15209 16201 15243 16235
rect 30113 16201 30147 16235
rect 34345 16201 34379 16235
rect 1501 16133 1535 16167
rect 4721 16133 4755 16167
rect 13921 16133 13955 16167
rect 16957 16133 16991 16167
rect 20821 16133 20855 16167
rect 29377 16133 29411 16167
rect 30389 16133 30423 16167
rect 3985 16065 4019 16099
rect 4077 16065 4111 16099
rect 4353 16065 4387 16099
rect 4537 16065 4571 16099
rect 4629 16065 4663 16099
rect 4813 16065 4847 16099
rect 7849 16065 7883 16099
rect 8401 16065 8435 16099
rect 9321 16065 9355 16099
rect 9413 16065 9447 16099
rect 9505 16065 9539 16099
rect 9689 16065 9723 16099
rect 13001 16065 13035 16099
rect 16129 16065 16163 16099
rect 17233 16065 17267 16099
rect 17325 16065 17359 16099
rect 17417 16065 17451 16099
rect 17601 16065 17635 16099
rect 17785 16065 17819 16099
rect 18981 16065 19015 16099
rect 19901 16065 19935 16099
rect 24317 16065 24351 16099
rect 24869 16065 24903 16099
rect 25605 16065 25639 16099
rect 25881 16065 25915 16099
rect 26065 16065 26099 16099
rect 26525 16065 26559 16099
rect 29193 16065 29227 16099
rect 29653 16065 29687 16099
rect 29837 16065 29871 16099
rect 30021 16065 30055 16099
rect 30205 16065 30239 16099
rect 30573 16065 30607 16099
rect 30757 16065 30791 16099
rect 30849 16065 30883 16099
rect 33977 16065 34011 16099
rect 37657 16065 37691 16099
rect 4261 15997 4295 16031
rect 8677 15997 8711 16031
rect 13093 15997 13127 16031
rect 13185 15997 13219 16031
rect 16221 15997 16255 16031
rect 25421 15997 25455 16031
rect 26341 15997 26375 16031
rect 26709 15997 26743 16031
rect 33885 15997 33919 16031
rect 4353 15929 4387 15963
rect 8033 15929 8067 15963
rect 9045 15929 9079 15963
rect 12633 15929 12667 15963
rect 16497 15929 16531 15963
rect 25789 15929 25823 15963
rect 1593 15861 1627 15895
rect 16221 15861 16255 15895
rect 17877 15861 17911 15895
rect 24409 15861 24443 15895
rect 25973 15861 26007 15895
rect 29561 15861 29595 15895
rect 29745 15861 29779 15895
rect 37841 15861 37875 15895
rect 3157 15657 3191 15691
rect 13829 15657 13863 15691
rect 16405 15657 16439 15691
rect 17325 15657 17359 15691
rect 17509 15657 17543 15691
rect 19349 15657 19383 15691
rect 26341 15657 26375 15691
rect 33333 15657 33367 15691
rect 12817 15589 12851 15623
rect 26801 15589 26835 15623
rect 26893 15589 26927 15623
rect 30389 15589 30423 15623
rect 32505 15589 32539 15623
rect 1409 15521 1443 15555
rect 4261 15521 4295 15555
rect 4445 15521 4479 15555
rect 8953 15521 8987 15555
rect 14473 15521 14507 15555
rect 15025 15521 15059 15555
rect 15485 15521 15519 15555
rect 27629 15521 27663 15555
rect 29745 15521 29779 15555
rect 30941 15521 30975 15555
rect 32045 15521 32079 15555
rect 32965 15521 32999 15555
rect 4169 15453 4203 15487
rect 8769 15453 8803 15487
rect 11069 15453 11103 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 14381 15453 14415 15487
rect 14657 15453 14691 15487
rect 15669 15453 15703 15487
rect 15853 15453 15887 15487
rect 15945 15453 15979 15487
rect 16681 15453 16715 15487
rect 16773 15453 16807 15487
rect 19349 15453 19383 15487
rect 20453 15453 20487 15487
rect 20913 15453 20947 15487
rect 21097 15453 21131 15487
rect 21189 15453 21223 15487
rect 22017 15453 22051 15487
rect 22385 15453 22419 15487
rect 22661 15453 22695 15487
rect 22937 15453 22971 15487
rect 23213 15453 23247 15487
rect 23397 15453 23431 15487
rect 23489 15453 23523 15487
rect 24869 15453 24903 15487
rect 25513 15453 25547 15487
rect 26709 15453 26743 15487
rect 26985 15453 27019 15487
rect 27537 15453 27571 15487
rect 28641 15453 28675 15487
rect 29929 15453 29963 15487
rect 30297 15453 30331 15487
rect 30481 15453 30515 15487
rect 31217 15453 31251 15487
rect 31401 15453 31435 15487
rect 32137 15453 32171 15487
rect 33057 15453 33091 15487
rect 1685 15385 1719 15419
rect 9229 15385 9263 15419
rect 10977 15385 11011 15419
rect 11345 15385 11379 15419
rect 16129 15385 16163 15419
rect 17141 15385 17175 15419
rect 22201 15385 22235 15419
rect 22293 15385 22327 15419
rect 30573 15385 30607 15419
rect 30757 15385 30791 15419
rect 3801 15317 3835 15351
rect 8585 15317 8619 15351
rect 16957 15317 16991 15351
rect 17341 15317 17375 15351
rect 20729 15317 20763 15351
rect 22569 15317 22603 15351
rect 26525 15317 26559 15351
rect 27905 15317 27939 15351
rect 28733 15317 28767 15351
rect 30113 15317 30147 15351
rect 31585 15317 31619 15351
rect 1961 15113 1995 15147
rect 2605 15113 2639 15147
rect 2973 15113 3007 15147
rect 3065 15113 3099 15147
rect 4721 15113 4755 15147
rect 8125 15113 8159 15147
rect 9505 15113 9539 15147
rect 9965 15113 9999 15147
rect 10885 15113 10919 15147
rect 11529 15113 11563 15147
rect 11897 15113 11931 15147
rect 11989 15113 12023 15147
rect 13369 15113 13403 15147
rect 16221 15113 16255 15147
rect 20177 15113 20211 15147
rect 26433 15113 26467 15147
rect 27629 15113 27663 15147
rect 33425 15113 33459 15147
rect 16037 15045 16071 15079
rect 19809 15045 19843 15079
rect 26065 15045 26099 15079
rect 26249 15045 26283 15079
rect 26617 15045 26651 15079
rect 29009 15045 29043 15079
rect 33057 15045 33091 15079
rect 33257 15045 33291 15079
rect 33793 15045 33827 15079
rect 2145 14977 2179 15011
rect 4353 14977 4387 15011
rect 4537 14977 4571 15011
rect 6377 14977 6411 15011
rect 9873 14977 9907 15011
rect 11069 14977 11103 15011
rect 13001 14977 13035 15011
rect 13185 14977 13219 15011
rect 13645 14977 13679 15011
rect 14565 14977 14599 15011
rect 15209 14977 15243 15011
rect 17693 14977 17727 15011
rect 17969 14977 18003 15011
rect 18153 14977 18187 15011
rect 18797 14977 18831 15011
rect 19165 14977 19199 15011
rect 20085 14977 20119 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 21005 14977 21039 15011
rect 21189 14977 21223 15011
rect 21281 14977 21315 15011
rect 23397 14977 23431 15011
rect 24593 14977 24627 15011
rect 24777 14977 24811 15011
rect 25513 14977 25547 15011
rect 25697 14977 25731 15011
rect 25789 14977 25823 15011
rect 25973 14977 26007 15011
rect 27813 14977 27847 15011
rect 27905 14977 27939 15011
rect 28089 14977 28123 15011
rect 28273 14977 28307 15011
rect 28457 14979 28491 15013
rect 28825 14977 28859 15011
rect 29193 14977 29227 15011
rect 29377 14977 29411 15011
rect 30849 14977 30883 15011
rect 31033 14977 31067 15011
rect 33517 14977 33551 15011
rect 3157 14909 3191 14943
rect 6653 14909 6687 14943
rect 10149 14909 10183 14943
rect 12081 14909 12115 14943
rect 14289 14909 14323 14943
rect 17509 14909 17543 14943
rect 23949 14909 23983 14943
rect 24961 14909 24995 14943
rect 28549 14909 28583 14943
rect 28641 14909 28675 14943
rect 30205 14909 30239 14943
rect 33793 14909 33827 14943
rect 15669 14841 15703 14875
rect 17877 14841 17911 14875
rect 27997 14841 28031 14875
rect 15025 14773 15059 14807
rect 16037 14773 16071 14807
rect 18245 14773 18279 14807
rect 20545 14773 20579 14807
rect 21373 14773 21407 14807
rect 25605 14773 25639 14807
rect 25789 14773 25823 14807
rect 26709 14773 26743 14807
rect 30849 14773 30883 14807
rect 33241 14773 33275 14807
rect 33609 14773 33643 14807
rect 6377 14569 6411 14603
rect 6561 14569 6595 14603
rect 13277 14569 13311 14603
rect 14381 14569 14415 14603
rect 16773 14569 16807 14603
rect 18889 14569 18923 14603
rect 19625 14569 19659 14603
rect 20085 14569 20119 14603
rect 22293 14569 22327 14603
rect 23489 14569 23523 14603
rect 27353 14569 27387 14603
rect 28181 14569 28215 14603
rect 31953 14569 31987 14603
rect 33333 14569 33367 14603
rect 15761 14501 15795 14535
rect 31125 14501 31159 14535
rect 33517 14501 33551 14535
rect 4629 14433 4663 14467
rect 7389 14433 7423 14467
rect 7573 14433 7607 14467
rect 15117 14433 15151 14467
rect 15393 14433 15427 14467
rect 17509 14433 17543 14467
rect 21189 14433 21223 14467
rect 21833 14433 21867 14467
rect 30573 14433 30607 14467
rect 33241 14433 33275 14467
rect 3893 14365 3927 14399
rect 4077 14365 4111 14399
rect 6745 14365 6779 14399
rect 11529 14365 11563 14399
rect 14289 14365 14323 14399
rect 14657 14365 14691 14399
rect 15301 14365 15335 14399
rect 15485 14365 15519 14399
rect 15577 14365 15611 14399
rect 15945 14365 15979 14399
rect 16037 14365 16071 14399
rect 16129 14365 16163 14399
rect 16405 14365 16439 14399
rect 16681 14365 16715 14399
rect 17785 14365 17819 14399
rect 18245 14365 18279 14399
rect 19901 14365 19935 14399
rect 19993 14365 20027 14399
rect 20453 14365 20487 14399
rect 20729 14365 20763 14399
rect 21465 14365 21499 14399
rect 22017 14365 22051 14399
rect 22109 14365 22143 14399
rect 22477 14365 22511 14399
rect 23305 14365 23339 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 27537 14365 27571 14399
rect 27721 14365 27755 14399
rect 27813 14365 27847 14399
rect 28365 14365 28399 14399
rect 28549 14365 28583 14399
rect 28641 14365 28675 14399
rect 30481 14365 30515 14399
rect 30665 14365 30699 14399
rect 31217 14365 31251 14399
rect 31401 14365 31435 14399
rect 31493 14365 31527 14399
rect 31585 14365 31619 14399
rect 31769 14365 31803 14399
rect 33149 14365 33183 14399
rect 4905 14297 4939 14331
rect 11805 14297 11839 14331
rect 18521 14297 18555 14331
rect 18613 14297 18647 14331
rect 18797 14297 18831 14331
rect 19257 14297 19291 14331
rect 19634 14297 19668 14331
rect 24961 14297 24995 14331
rect 30757 14297 30791 14331
rect 30941 14297 30975 14331
rect 3985 14229 4019 14263
rect 6929 14229 6963 14263
rect 7297 14229 7331 14263
rect 14841 14229 14875 14263
rect 16313 14229 16347 14263
rect 16957 14229 16991 14263
rect 4077 14025 4111 14059
rect 4645 14025 4679 14059
rect 4813 14025 4847 14059
rect 5273 14025 5307 14059
rect 6377 14025 6411 14059
rect 11621 14025 11655 14059
rect 12449 14025 12483 14059
rect 14197 14025 14231 14059
rect 14939 14025 14973 14059
rect 15485 14025 15519 14059
rect 16221 14025 16255 14059
rect 18797 14025 18831 14059
rect 20637 14025 20671 14059
rect 23305 14025 23339 14059
rect 25053 14025 25087 14059
rect 28549 14025 28583 14059
rect 31217 14025 31251 14059
rect 33609 14025 33643 14059
rect 4445 13957 4479 13991
rect 6837 13957 6871 13991
rect 10241 13957 10275 13991
rect 12081 13957 12115 13991
rect 14105 13957 14139 13991
rect 22845 13957 22879 13991
rect 3985 13889 4019 13923
rect 5457 13889 5491 13923
rect 6745 13889 6779 13923
rect 7757 13889 7791 13923
rect 10057 13889 10091 13923
rect 11989 13889 12023 13923
rect 12633 13889 12667 13923
rect 14841 13889 14875 13923
rect 15025 13889 15059 13923
rect 15117 13889 15151 13923
rect 15393 13889 15427 13923
rect 15577 13889 15611 13923
rect 16129 13889 16163 13923
rect 16313 13889 16347 13923
rect 17601 13889 17635 13923
rect 17785 13889 17819 13923
rect 18245 13889 18279 13923
rect 18337 13889 18371 13923
rect 18521 13889 18555 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 20545 13889 20579 13923
rect 21097 13889 21131 13923
rect 22661 13889 22695 13923
rect 23489 13889 23523 13923
rect 24225 13889 24259 13923
rect 24777 13889 24811 13923
rect 25237 13889 25271 13923
rect 25329 13889 25363 13923
rect 25513 13889 25547 13923
rect 25605 13889 25639 13923
rect 25697 13889 25731 13923
rect 25881 13889 25915 13923
rect 26249 13889 26283 13923
rect 26433 13889 26467 13923
rect 26985 13889 27019 13923
rect 27169 13889 27203 13923
rect 28457 13889 28491 13923
rect 28641 13889 28675 13923
rect 31033 13889 31067 13923
rect 33149 13889 33183 13923
rect 33517 13889 33551 13923
rect 33701 13889 33735 13923
rect 1409 13821 1443 13855
rect 1685 13821 1719 13855
rect 4261 13821 4295 13855
rect 7021 13821 7055 13855
rect 9873 13821 9907 13855
rect 12173 13821 12207 13855
rect 17233 13821 17267 13855
rect 21373 13821 21407 13855
rect 22477 13821 22511 13855
rect 23765 13821 23799 13855
rect 24041 13821 24075 13855
rect 30849 13821 30883 13855
rect 33425 13821 33459 13855
rect 3617 13753 3651 13787
rect 24685 13753 24719 13787
rect 33241 13753 33275 13787
rect 3157 13685 3191 13719
rect 4629 13685 4663 13719
rect 8020 13685 8054 13719
rect 9505 13685 9539 13719
rect 23673 13685 23707 13719
rect 25789 13685 25823 13719
rect 26249 13685 26283 13719
rect 27077 13685 27111 13719
rect 33333 13685 33367 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 3801 13481 3835 13515
rect 6561 13481 6595 13515
rect 8217 13481 8251 13515
rect 12449 13481 12483 13515
rect 14933 13481 14967 13515
rect 17417 13481 17451 13515
rect 21189 13481 21223 13515
rect 22201 13481 22235 13515
rect 24685 13481 24719 13515
rect 28273 13481 28307 13515
rect 29193 13481 29227 13515
rect 31953 13481 31987 13515
rect 32137 13481 32171 13515
rect 33793 13481 33827 13515
rect 2513 13413 2547 13447
rect 8953 13413 8987 13447
rect 32689 13413 32723 13447
rect 2973 13345 3007 13379
rect 3065 13345 3099 13379
rect 9597 13345 9631 13379
rect 9781 13345 9815 13379
rect 12909 13345 12943 13379
rect 13093 13345 13127 13379
rect 18797 13345 18831 13379
rect 23121 13345 23155 13379
rect 25697 13345 25731 13379
rect 29377 13345 29411 13379
rect 31861 13345 31895 13379
rect 32873 13345 32907 13379
rect 2145 13277 2179 13311
rect 2881 13277 2915 13311
rect 3801 13277 3835 13311
rect 4077 13277 4111 13311
rect 8401 13277 8435 13311
rect 9965 13277 9999 13311
rect 15117 13277 15151 13311
rect 15209 13277 15243 13311
rect 15393 13277 15427 13311
rect 15485 13277 15519 13311
rect 17417 13277 17451 13311
rect 17601 13277 17635 13311
rect 20269 13277 20303 13311
rect 20453 13277 20487 13311
rect 20545 13277 20579 13311
rect 20638 13277 20672 13311
rect 20913 13277 20947 13311
rect 21833 13277 21867 13311
rect 22017 13277 22051 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 23306 13277 23340 13311
rect 23397 13277 23431 13311
rect 23489 13277 23523 13311
rect 23581 13277 23615 13311
rect 24869 13277 24903 13311
rect 24961 13277 24995 13311
rect 25145 13277 25179 13311
rect 25237 13277 25271 13311
rect 25605 13277 25639 13311
rect 25789 13277 25823 13311
rect 26065 13277 26099 13311
rect 26249 13277 26283 13311
rect 26341 13277 26375 13311
rect 26433 13277 26467 13311
rect 26617 13277 26651 13311
rect 27077 13277 27111 13311
rect 27169 13277 27203 13311
rect 27353 13277 27387 13311
rect 27445 13277 27479 13311
rect 28457 13277 28491 13311
rect 28549 13277 28583 13311
rect 28641 13277 28675 13311
rect 28733 13277 28767 13311
rect 29101 13277 29135 13311
rect 30481 13277 30515 13311
rect 30665 13277 30699 13311
rect 30757 13277 30791 13311
rect 30849 13277 30883 13311
rect 31033 13277 31067 13311
rect 31217 13277 31251 13311
rect 31585 13277 31619 13311
rect 32965 13277 32999 13311
rect 33517 13277 33551 13311
rect 33609 13277 33643 13311
rect 33885 13277 33919 13311
rect 34069 13277 34103 13311
rect 1501 13209 1535 13243
rect 3985 13209 4019 13243
rect 5273 13209 5307 13243
rect 9413 13209 9447 13243
rect 18613 13209 18647 13243
rect 18705 13209 18739 13243
rect 21005 13209 21039 13243
rect 21205 13209 21239 13243
rect 22753 13209 22787 13243
rect 26801 13209 26835 13243
rect 33241 13209 33275 13243
rect 33333 13209 33367 13243
rect 9321 13141 9355 13175
rect 10149 13141 10183 13175
rect 12817 13141 12851 13175
rect 18245 13141 18279 13175
rect 21373 13141 21407 13175
rect 26893 13141 26927 13175
rect 28825 13141 28859 13175
rect 29377 13141 29411 13175
rect 34253 13141 34287 13175
rect 4261 12937 4295 12971
rect 6377 12937 6411 12971
rect 6837 12937 6871 12971
rect 9321 12937 9355 12971
rect 10609 12937 10643 12971
rect 11069 12937 11103 12971
rect 16221 12937 16255 12971
rect 20453 12937 20487 12971
rect 23397 12937 23431 12971
rect 29193 12937 29227 12971
rect 31125 12937 31159 12971
rect 32505 12937 32539 12971
rect 33057 12937 33091 12971
rect 33885 12937 33919 12971
rect 8769 12869 8803 12903
rect 16037 12869 16071 12903
rect 20913 12869 20947 12903
rect 21113 12869 21147 12903
rect 23581 12869 23615 12903
rect 31401 12869 31435 12903
rect 31585 12869 31619 12903
rect 31801 12869 31835 12903
rect 32321 12869 32355 12903
rect 2237 12801 2271 12835
rect 3433 12801 3467 12835
rect 5917 12801 5951 12835
rect 6745 12801 6779 12835
rect 10517 12801 10551 12835
rect 10977 12801 11011 12835
rect 13185 12801 13219 12835
rect 13277 12801 13311 12835
rect 18245 12801 18279 12835
rect 18429 12801 18463 12835
rect 20269 12801 20303 12835
rect 22661 12801 22695 12835
rect 22845 12801 22879 12835
rect 23213 12801 23247 12835
rect 23305 12801 23339 12835
rect 23765 12801 23799 12835
rect 26341 12801 26375 12835
rect 26525 12801 26559 12835
rect 27261 12801 27295 12835
rect 27353 12801 27387 12835
rect 27445 12801 27479 12835
rect 27629 12801 27663 12835
rect 28825 12801 28859 12835
rect 29285 12801 29319 12835
rect 29469 12801 29503 12835
rect 30757 12801 30791 12835
rect 31309 12801 31343 12835
rect 31493 12801 31527 12835
rect 32137 12801 32171 12835
rect 32965 12801 32999 12835
rect 33425 12801 33459 12835
rect 33793 12801 33827 12835
rect 33977 12801 34011 12835
rect 2881 12733 2915 12767
rect 3525 12733 3559 12767
rect 3801 12733 3835 12767
rect 4353 12733 4387 12767
rect 4445 12733 4479 12767
rect 7021 12733 7055 12767
rect 9229 12733 9263 12767
rect 11253 12733 11287 12767
rect 13369 12733 13403 12767
rect 20637 12733 20671 12767
rect 21833 12733 21867 12767
rect 22109 12733 22143 12767
rect 22293 12733 22327 12767
rect 22385 12733 22419 12767
rect 28917 12733 28951 12767
rect 30665 12733 30699 12767
rect 8769 12665 8803 12699
rect 22937 12665 22971 12699
rect 26433 12665 26467 12699
rect 29285 12665 29319 12699
rect 31953 12665 31987 12699
rect 3893 12597 3927 12631
rect 5733 12597 5767 12631
rect 9505 12597 9539 12631
rect 10333 12597 10367 12631
rect 12817 12597 12851 12631
rect 16221 12597 16255 12631
rect 16405 12597 16439 12631
rect 20729 12597 20763 12631
rect 21097 12597 21131 12631
rect 21281 12597 21315 12631
rect 23857 12597 23891 12631
rect 26985 12597 27019 12631
rect 31769 12597 31803 12631
rect 8585 12393 8619 12427
rect 19441 12393 19475 12427
rect 19901 12393 19935 12427
rect 21373 12393 21407 12427
rect 21833 12393 21867 12427
rect 24409 12393 24443 12427
rect 26249 12393 26283 12427
rect 28641 12393 28675 12427
rect 29561 12393 29595 12427
rect 8953 12325 8987 12359
rect 9321 12325 9355 12359
rect 19625 12325 19659 12359
rect 23397 12325 23431 12359
rect 23489 12325 23523 12359
rect 25237 12325 25271 12359
rect 2881 12257 2915 12291
rect 5181 12257 5215 12291
rect 10241 12257 10275 12291
rect 12265 12257 12299 12291
rect 15393 12257 15427 12291
rect 15577 12257 15611 12291
rect 18429 12257 18463 12291
rect 22845 12257 22879 12291
rect 22937 12257 22971 12291
rect 23121 12257 23155 12291
rect 23581 12257 23615 12291
rect 24869 12257 24903 12291
rect 25145 12257 25179 12291
rect 25329 12257 25363 12291
rect 26801 12257 26835 12291
rect 29745 12257 29779 12291
rect 29837 12257 29871 12291
rect 1961 12189 1995 12223
rect 2697 12189 2731 12223
rect 7205 12189 7239 12223
rect 8309 12189 8343 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9413 12189 9447 12223
rect 9597 12189 9631 12223
rect 9781 12189 9815 12223
rect 10057 12189 10091 12223
rect 13093 12189 13127 12223
rect 15945 12189 15979 12223
rect 17969 12189 18003 12223
rect 18153 12189 18187 12223
rect 21005 12189 21039 12223
rect 21373 12189 21407 12223
rect 23029 12189 23063 12223
rect 23305 12189 23339 12223
rect 24593 12189 24627 12223
rect 24685 12189 24719 12223
rect 24777 12189 24811 12223
rect 25053 12189 25087 12223
rect 28917 12189 28951 12223
rect 29285 12189 29319 12223
rect 29377 12189 29411 12223
rect 30205 12189 30239 12223
rect 30573 12189 30607 12223
rect 30757 12189 30791 12223
rect 2605 12121 2639 12155
rect 5457 12121 5491 12155
rect 10517 12121 10551 12155
rect 16221 12121 16255 12155
rect 19257 12121 19291 12155
rect 19462 12121 19496 12155
rect 19717 12121 19751 12155
rect 21649 12121 21683 12155
rect 29009 12121 29043 12155
rect 1777 12053 1811 12087
rect 2237 12053 2271 12087
rect 8769 12053 8803 12087
rect 9965 12053 9999 12087
rect 12909 12053 12943 12087
rect 14933 12053 14967 12087
rect 15301 12053 15335 12087
rect 19917 12053 19951 12087
rect 20085 12053 20119 12087
rect 21557 12053 21591 12087
rect 21849 12053 21883 12087
rect 22017 12053 22051 12087
rect 22661 12053 22695 12087
rect 26617 12053 26651 12087
rect 26709 12053 26743 12087
rect 29101 12053 29135 12087
rect 30021 12053 30055 12087
rect 30113 12053 30147 12087
rect 30665 12053 30699 12087
rect 3157 11849 3191 11883
rect 6009 11849 6043 11883
rect 15485 11849 15519 11883
rect 24225 11849 24259 11883
rect 25053 11849 25087 11883
rect 25513 11849 25547 11883
rect 29377 11849 29411 11883
rect 30021 11849 30055 11883
rect 32965 11849 32999 11883
rect 1685 11781 1719 11815
rect 6653 11781 6687 11815
rect 12357 11781 12391 11815
rect 13185 11781 13219 11815
rect 14933 11781 14967 11815
rect 26985 11781 27019 11815
rect 27201 11781 27235 11815
rect 30665 11781 30699 11815
rect 1409 11713 1443 11747
rect 6193 11713 6227 11747
rect 8493 11713 8527 11747
rect 9137 11713 9171 11747
rect 15669 11713 15703 11747
rect 17877 11713 17911 11747
rect 19533 11713 19567 11747
rect 19625 11713 19659 11747
rect 19717 11713 19751 11747
rect 19901 11713 19935 11747
rect 21189 11713 21223 11747
rect 22661 11713 22695 11747
rect 22937 11713 22971 11747
rect 24041 11713 24075 11747
rect 24317 11713 24351 11747
rect 24409 11713 24443 11747
rect 24593 11713 24627 11747
rect 25421 11713 25455 11747
rect 29101 11713 29135 11747
rect 29193 11713 29227 11747
rect 30481 11713 30515 11747
rect 31309 11713 31343 11747
rect 32873 11713 32907 11747
rect 33057 11713 33091 11747
rect 33333 11713 33367 11747
rect 33609 11713 33643 11747
rect 33793 11713 33827 11747
rect 6377 11645 6411 11679
rect 8401 11645 8435 11679
rect 8769 11645 8803 11679
rect 12449 11645 12483 11679
rect 12541 11645 12575 11679
rect 12909 11645 12943 11679
rect 24501 11645 24535 11679
rect 25605 11645 25639 11679
rect 29377 11645 29411 11679
rect 30205 11645 30239 11679
rect 30297 11645 30331 11679
rect 30389 11645 30423 11679
rect 31033 11645 31067 11679
rect 31125 11645 31159 11679
rect 33149 11645 33183 11679
rect 9597 11577 9631 11611
rect 19257 11577 19291 11611
rect 21373 11577 21407 11611
rect 27353 11577 27387 11611
rect 33885 11577 33919 11611
rect 8769 11509 8803 11543
rect 9045 11509 9079 11543
rect 9413 11509 9447 11543
rect 11989 11509 12023 11543
rect 17969 11509 18003 11543
rect 22753 11509 22787 11543
rect 24041 11509 24075 11543
rect 27169 11509 27203 11543
rect 33517 11509 33551 11543
rect 6653 11305 6687 11339
rect 10057 11305 10091 11339
rect 13277 11305 13311 11339
rect 14197 11305 14231 11339
rect 24501 11305 24535 11339
rect 25513 11305 25547 11339
rect 27629 11305 27663 11339
rect 29561 11305 29595 11339
rect 31861 11305 31895 11339
rect 32597 11305 32631 11339
rect 1685 11237 1719 11271
rect 3801 11237 3835 11271
rect 9597 11237 9631 11271
rect 14565 11237 14599 11271
rect 4353 11169 4387 11203
rect 7113 11169 7147 11203
rect 7205 11169 7239 11203
rect 13737 11169 13771 11203
rect 15209 11169 15243 11203
rect 26801 11169 26835 11203
rect 1501 11101 1535 11135
rect 2513 11101 2547 11135
rect 3433 11101 3467 11135
rect 4629 11101 4663 11135
rect 4813 11101 4847 11135
rect 8953 11101 8987 11135
rect 9438 11101 9472 11135
rect 9689 11101 9723 11135
rect 9873 11101 9907 11135
rect 10425 11101 10459 11135
rect 10517 11101 10551 11135
rect 11529 11101 11563 11135
rect 13461 11101 13495 11135
rect 14105 11101 14139 11135
rect 15025 11101 15059 11135
rect 15577 11101 15611 11135
rect 17325 11101 17359 11135
rect 17693 11101 17727 11135
rect 18245 11101 18279 11135
rect 18521 11101 18555 11135
rect 18705 11101 18739 11135
rect 20269 11101 20303 11135
rect 24409 11101 24443 11135
rect 24593 11101 24627 11135
rect 25421 11101 25455 11135
rect 25605 11101 25639 11135
rect 25697 11101 25731 11135
rect 25881 11101 25915 11135
rect 26617 11101 26651 11135
rect 27261 11101 27295 11135
rect 27445 11101 27479 11135
rect 27537 11101 27571 11135
rect 27813 11101 27847 11135
rect 28089 11101 28123 11135
rect 28181 11101 28215 11135
rect 28365 11101 28399 11135
rect 29745 11101 29779 11135
rect 29929 11101 29963 11135
rect 30021 11101 30055 11135
rect 32045 11101 32079 11135
rect 32321 11101 32355 11135
rect 32505 11101 32539 11135
rect 32781 11101 32815 11135
rect 33057 11101 33091 11135
rect 33241 11101 33275 11135
rect 37565 11101 37599 11135
rect 2329 11033 2363 11067
rect 2697 11033 2731 11067
rect 4169 11033 4203 11067
rect 7021 11033 7055 11067
rect 9321 11033 9355 11067
rect 11805 11033 11839 11067
rect 18429 11033 18463 11067
rect 18889 11033 18923 11067
rect 19257 11033 19291 11067
rect 19993 11033 20027 11067
rect 27077 11033 27111 11067
rect 27997 11033 28031 11067
rect 28273 11033 28307 11067
rect 37933 11033 37967 11067
rect 3249 10965 3283 10999
rect 4261 10965 4295 10999
rect 4721 10965 4755 10999
rect 9229 10965 9263 10999
rect 10701 10965 10735 10999
rect 14933 10965 14967 10999
rect 15393 10965 15427 10999
rect 20453 10965 20487 10999
rect 25881 10965 25915 10999
rect 26249 10965 26283 10999
rect 26709 10965 26743 10999
rect 4629 10761 4663 10795
rect 5089 10761 5123 10795
rect 11805 10761 11839 10795
rect 14289 10761 14323 10795
rect 21373 10761 21407 10795
rect 22845 10761 22879 10795
rect 34897 10761 34931 10795
rect 3065 10693 3099 10727
rect 6101 10693 6135 10727
rect 13553 10693 13587 10727
rect 15025 10693 15059 10727
rect 17601 10693 17635 10727
rect 22017 10693 22051 10727
rect 4997 10625 5031 10659
rect 5733 10625 5767 10659
rect 5917 10625 5951 10659
rect 6561 10625 6595 10659
rect 7849 10625 7883 10659
rect 10425 10625 10459 10659
rect 11989 10625 12023 10659
rect 13461 10625 13495 10659
rect 14749 10625 14783 10659
rect 16865 10625 16899 10659
rect 18061 10625 18095 10659
rect 18705 10625 18739 10659
rect 20085 10625 20119 10659
rect 20177 10625 20211 10659
rect 20269 10625 20303 10659
rect 21189 10625 21223 10659
rect 21465 10625 21499 10659
rect 21833 10625 21867 10659
rect 22109 10625 22143 10659
rect 22201 10625 22235 10659
rect 22477 10625 22511 10659
rect 22661 10625 22695 10659
rect 22937 10625 22971 10659
rect 23489 10625 23523 10659
rect 23581 10625 23615 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 27353 10625 27387 10659
rect 27537 10625 27571 10659
rect 28549 10625 28583 10659
rect 28641 10625 28675 10659
rect 28917 10625 28951 10659
rect 29101 10625 29135 10659
rect 30757 10625 30791 10659
rect 30941 10625 30975 10659
rect 32689 10625 32723 10659
rect 33149 10625 33183 10659
rect 34529 10625 34563 10659
rect 36553 10625 36587 10659
rect 36737 10625 36771 10659
rect 2789 10557 2823 10591
rect 5181 10557 5215 10591
rect 10241 10557 10275 10591
rect 13737 10557 13771 10591
rect 14381 10557 14415 10591
rect 14473 10557 14507 10591
rect 16497 10557 16531 10591
rect 27261 10557 27295 10591
rect 30849 10557 30883 10591
rect 32597 10557 32631 10591
rect 34621 10557 34655 10591
rect 4537 10489 4571 10523
rect 9137 10489 9171 10523
rect 13093 10489 13127 10523
rect 19073 10489 19107 10523
rect 20453 10489 20487 10523
rect 28733 10489 28767 10523
rect 29193 10489 29227 10523
rect 33057 10489 33091 10523
rect 6377 10421 6411 10455
rect 10609 10421 10643 10455
rect 13921 10421 13955 10455
rect 21189 10421 21223 10455
rect 22385 10421 22419 10455
rect 23765 10421 23799 10455
rect 27721 10421 27755 10455
rect 33241 10421 33275 10455
rect 36921 10421 36955 10455
rect 4629 10217 4663 10251
rect 4721 10217 4755 10251
rect 5996 10217 6030 10251
rect 8033 10217 8067 10251
rect 9413 10217 9447 10251
rect 16957 10217 16991 10251
rect 35173 10217 35207 10251
rect 14105 10149 14139 10183
rect 19073 10149 19107 10183
rect 21097 10149 21131 10183
rect 22201 10149 22235 10183
rect 24409 10149 24443 10183
rect 34253 10149 34287 10183
rect 4261 10081 4295 10115
rect 5733 10081 5767 10115
rect 8125 10081 8159 10115
rect 8401 10081 8435 10115
rect 8493 10081 8527 10115
rect 8677 10081 8711 10115
rect 10333 10081 10367 10115
rect 15209 10081 15243 10115
rect 17417 10081 17451 10115
rect 17877 10081 17911 10115
rect 19257 10081 19291 10115
rect 20637 10081 20671 10115
rect 21373 10081 21407 10115
rect 21465 10081 21499 10115
rect 21557 10081 21591 10115
rect 24869 10081 24903 10115
rect 24961 10081 24995 10115
rect 34805 10081 34839 10115
rect 2789 10013 2823 10047
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 3157 10013 3191 10047
rect 4445 10013 4479 10047
rect 4721 10013 4755 10047
rect 4905 10013 4939 10047
rect 7849 10013 7883 10047
rect 7941 10013 7975 10047
rect 8585 10013 8619 10047
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 10241 10013 10275 10047
rect 14289 10013 14323 10047
rect 14565 10013 14599 10047
rect 15025 10013 15059 10047
rect 17785 10013 17819 10047
rect 18153 10013 18187 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 18613 10013 18647 10047
rect 18705 10013 18739 10047
rect 18798 10013 18832 10047
rect 19441 10013 19475 10047
rect 20085 10013 20119 10047
rect 20361 10013 20395 10047
rect 20545 10013 20579 10047
rect 20821 10013 20855 10047
rect 21281 10013 21315 10047
rect 21741 10013 21775 10047
rect 22385 10013 22419 10047
rect 22477 10013 22511 10047
rect 22661 10013 22695 10047
rect 22753 10013 22787 10047
rect 23029 10013 23063 10047
rect 23121 10013 23155 10047
rect 23213 10013 23247 10047
rect 23489 10013 23523 10047
rect 26985 10013 27019 10047
rect 27077 10013 27111 10047
rect 27169 10013 27203 10047
rect 27353 10013 27387 10047
rect 28549 10013 28583 10047
rect 28733 10013 28767 10047
rect 29009 10013 29043 10047
rect 29193 10013 29227 10047
rect 29653 10023 29687 10057
rect 29837 10013 29871 10047
rect 30205 10013 30239 10047
rect 30389 10013 30423 10047
rect 30481 10013 30515 10047
rect 30573 10013 30607 10047
rect 30757 10013 30791 10047
rect 31217 10013 31251 10047
rect 31585 10013 31619 10047
rect 33793 10013 33827 10047
rect 33885 10013 33919 10047
rect 33977 10013 34011 10047
rect 34161 10013 34195 10047
rect 34529 10013 34563 10047
rect 34897 10013 34931 10047
rect 7757 9945 7791 9979
rect 10609 9945 10643 9979
rect 14473 9945 14507 9979
rect 15485 9945 15519 9979
rect 21005 9945 21039 9979
rect 23351 9945 23385 9979
rect 33517 9945 33551 9979
rect 34253 9945 34287 9979
rect 2513 9877 2547 9911
rect 8217 9877 8251 9911
rect 9597 9877 9631 9911
rect 10057 9877 10091 9911
rect 12081 9877 12115 9911
rect 14841 9877 14875 9911
rect 19625 9877 19659 9911
rect 20177 9877 20211 9911
rect 20453 9877 20487 9911
rect 22845 9877 22879 9911
rect 24777 9877 24811 9911
rect 26709 9877 26743 9911
rect 28917 9877 28951 9911
rect 29101 9877 29135 9911
rect 29837 9877 29871 9911
rect 30941 9877 30975 9911
rect 32229 9877 32263 9911
rect 34437 9877 34471 9911
rect 6469 9673 6503 9707
rect 6929 9673 6963 9707
rect 10609 9673 10643 9707
rect 11069 9673 11103 9707
rect 22937 9673 22971 9707
rect 25053 9673 25087 9707
rect 29837 9673 29871 9707
rect 4537 9605 4571 9639
rect 6837 9605 6871 9639
rect 10977 9605 11011 9639
rect 19533 9605 19567 9639
rect 21097 9605 21131 9639
rect 21297 9605 21331 9639
rect 24777 9605 24811 9639
rect 32689 9605 32723 9639
rect 32873 9605 32907 9639
rect 33057 9605 33091 9639
rect 1409 9537 1443 9571
rect 4169 9537 4203 9571
rect 4353 9537 4387 9571
rect 4445 9537 4479 9571
rect 4793 9537 4827 9571
rect 4905 9537 4939 9571
rect 4997 9537 5031 9571
rect 5181 9537 5215 9571
rect 8401 9537 8435 9571
rect 8493 9537 8527 9571
rect 8677 9537 8711 9571
rect 8769 9537 8803 9571
rect 8867 9537 8901 9571
rect 9045 9537 9079 9571
rect 12265 9537 12299 9571
rect 12725 9537 12759 9571
rect 14197 9537 14231 9571
rect 17877 9537 17911 9571
rect 20637 9537 20671 9571
rect 20821 9537 20855 9571
rect 20913 9537 20947 9571
rect 22569 9537 22603 9571
rect 22753 9537 22787 9571
rect 24547 9537 24581 9571
rect 24685 9537 24719 9571
rect 24869 9537 24903 9571
rect 25605 9537 25639 9571
rect 25881 9537 25915 9571
rect 26249 9537 26283 9571
rect 27169 9537 27203 9571
rect 27445 9537 27479 9571
rect 27629 9537 27663 9571
rect 28917 9537 28951 9571
rect 29101 9537 29135 9571
rect 29745 9537 29779 9571
rect 29929 9537 29963 9571
rect 30849 9537 30883 9571
rect 31217 9537 31251 9571
rect 31677 9537 31711 9571
rect 1685 9469 1719 9503
rect 7113 9469 7147 9503
rect 8953 9469 8987 9503
rect 11161 9469 11195 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 14289 9469 14323 9503
rect 14473 9469 14507 9503
rect 18153 9469 18187 9503
rect 26065 9469 26099 9503
rect 26433 9469 26467 9503
rect 30665 9469 30699 9503
rect 4169 9401 4203 9435
rect 12357 9401 12391 9435
rect 19809 9401 19843 9435
rect 31217 9401 31251 9435
rect 3157 9333 3191 9367
rect 8217 9333 8251 9367
rect 12081 9333 12115 9367
rect 13829 9333 13863 9367
rect 20637 9333 20671 9367
rect 21281 9333 21315 9367
rect 21465 9333 21499 9367
rect 22753 9333 22787 9367
rect 25697 9333 25731 9367
rect 26985 9333 27019 9367
rect 29285 9333 29319 9367
rect 1961 9129 1995 9163
rect 5181 9129 5215 9163
rect 8033 9129 8067 9163
rect 12246 9129 12280 9163
rect 17693 9129 17727 9163
rect 22753 9129 22787 9163
rect 23765 9129 23799 9163
rect 27629 9129 27663 9163
rect 29745 9129 29779 9163
rect 31861 9129 31895 9163
rect 32597 9129 32631 9163
rect 33057 9129 33091 9163
rect 33517 9129 33551 9163
rect 2329 9061 2363 9095
rect 3985 9061 4019 9095
rect 5273 9061 5307 9095
rect 32229 9061 32263 9095
rect 2789 8993 2823 9027
rect 2973 8993 3007 9027
rect 4445 8993 4479 9027
rect 4537 8993 4571 9027
rect 8217 8993 8251 9027
rect 15485 8993 15519 9027
rect 17785 8993 17819 9027
rect 21189 8993 21223 9027
rect 22937 8993 22971 9027
rect 23305 8993 23339 9027
rect 25789 8993 25823 9027
rect 29653 8993 29687 9027
rect 37657 8993 37691 9027
rect 1501 8925 1535 8959
rect 2145 8925 2179 8959
rect 2697 8925 2731 8959
rect 3341 8925 3375 8959
rect 5273 8925 5307 8959
rect 5457 8925 5491 8959
rect 7941 8925 7975 8959
rect 8309 8925 8343 8959
rect 9873 8925 9907 8959
rect 9965 8925 9999 8959
rect 10057 8925 10091 8959
rect 10241 8925 10275 8959
rect 11989 8925 12023 8959
rect 15301 8925 15335 8959
rect 17325 8925 17359 8959
rect 17509 8925 17543 8959
rect 17969 8925 18003 8959
rect 19349 8925 19383 8959
rect 20177 8925 20211 8959
rect 20545 8925 20579 8959
rect 21097 8925 21131 8959
rect 23029 8925 23063 8959
rect 23397 8925 23431 8959
rect 23673 8925 23707 8959
rect 24041 8925 24075 8959
rect 24133 8925 24167 8959
rect 24225 8925 24259 8959
rect 24409 8925 24443 8959
rect 24502 8925 24536 8959
rect 24874 8925 24908 8959
rect 25513 8925 25547 8959
rect 25605 8925 25639 8959
rect 25881 8925 25915 8959
rect 26249 8925 26283 8959
rect 26341 8925 26375 8959
rect 26433 8925 26467 8959
rect 26617 8925 26651 8959
rect 26893 8925 26927 8959
rect 27077 8925 27111 8959
rect 27169 8925 27203 8959
rect 27261 8925 27295 8959
rect 27445 8925 27479 8959
rect 28437 8925 28471 8959
rect 28549 8925 28583 8959
rect 28641 8925 28675 8959
rect 28825 8925 28859 8959
rect 29561 8925 29595 8959
rect 31585 8925 31619 8959
rect 31677 8925 31711 8959
rect 31953 8925 31987 8959
rect 32137 8925 32171 8959
rect 32781 8925 32815 8959
rect 32873 8925 32907 8959
rect 33149 8925 33183 8959
rect 33241 8925 33275 8959
rect 33517 8925 33551 8959
rect 33701 8925 33735 8959
rect 37473 8925 37507 8959
rect 3157 8857 3191 8891
rect 4813 8857 4847 8891
rect 4997 8857 5031 8891
rect 8401 8857 8435 8891
rect 18153 8857 18187 8891
rect 24685 8857 24719 8891
rect 24777 8857 24811 8891
rect 25329 8857 25363 8891
rect 1593 8789 1627 8823
rect 3525 8789 3559 8823
rect 4353 8789 4387 8823
rect 9597 8789 9631 8823
rect 13737 8789 13771 8823
rect 14933 8789 14967 8823
rect 15393 8789 15427 8823
rect 20729 8789 20763 8823
rect 21373 8789 21407 8823
rect 25053 8789 25087 8823
rect 25973 8789 26007 8823
rect 28181 8789 28215 8823
rect 29929 8789 29963 8823
rect 31217 8789 31251 8823
rect 4553 8585 4587 8619
rect 4721 8585 4755 8619
rect 7113 8585 7147 8619
rect 7665 8585 7699 8619
rect 8033 8585 8067 8619
rect 8861 8585 8895 8619
rect 20821 8585 20855 8619
rect 25145 8585 25179 8619
rect 27353 8585 27387 8619
rect 28917 8585 28951 8619
rect 31401 8585 31435 8619
rect 4353 8517 4387 8551
rect 19257 8517 19291 8551
rect 19625 8517 19659 8551
rect 23305 8517 23339 8551
rect 27169 8517 27203 8551
rect 2329 8449 2363 8483
rect 2881 8449 2915 8483
rect 2973 8449 3007 8483
rect 3065 8449 3099 8483
rect 3249 8449 3283 8483
rect 7021 8449 7055 8483
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 12357 8449 12391 8483
rect 14289 8449 14323 8483
rect 14381 8449 14415 8483
rect 16405 8449 16439 8483
rect 16681 8449 16715 8483
rect 18521 8449 18555 8483
rect 19533 8449 19567 8483
rect 19717 8449 19751 8483
rect 20085 8449 20119 8483
rect 20177 8449 20211 8483
rect 20269 8449 20303 8483
rect 20637 8449 20671 8483
rect 20913 8449 20947 8483
rect 22385 8449 22419 8483
rect 22477 8449 22511 8483
rect 22845 8449 22879 8483
rect 22937 8449 22971 8483
rect 23085 8449 23119 8483
rect 23213 8449 23247 8483
rect 23443 8449 23477 8483
rect 26985 8449 27019 8483
rect 28365 8449 28399 8483
rect 28549 8449 28583 8483
rect 28825 8449 28859 8483
rect 29009 8449 29043 8483
rect 29929 8449 29963 8483
rect 30113 8449 30147 8483
rect 31401 8449 31435 8483
rect 31585 8449 31619 8483
rect 33057 8449 33091 8483
rect 7205 8381 7239 8415
rect 8125 8381 8159 8415
rect 8217 8381 8251 8415
rect 14657 8381 14691 8415
rect 16129 8381 16163 8415
rect 16957 8381 16991 8415
rect 18429 8381 18463 8415
rect 19993 8381 20027 8415
rect 22753 8381 22787 8415
rect 25237 8381 25271 8415
rect 25329 8381 25363 8415
rect 30297 8381 30331 8415
rect 31769 8381 31803 8415
rect 32965 8381 32999 8415
rect 2605 8313 2639 8347
rect 14105 8313 14139 8347
rect 16221 8313 16255 8347
rect 19809 8313 19843 8347
rect 22201 8313 22235 8347
rect 24777 8313 24811 8347
rect 33425 8313 33459 8347
rect 4537 8245 4571 8279
rect 6653 8245 6687 8279
rect 12633 8245 12667 8279
rect 20453 8245 20487 8279
rect 23581 8245 23615 8279
rect 28365 8245 28399 8279
rect 7481 8041 7515 8075
rect 7941 8041 7975 8075
rect 10885 8041 10919 8075
rect 11989 8041 12023 8075
rect 14289 8041 14323 8075
rect 28825 8041 28859 8075
rect 29193 8041 29227 8075
rect 31953 8041 31987 8075
rect 12725 7973 12759 8007
rect 19717 7973 19751 8007
rect 4721 7905 4755 7939
rect 4997 7905 5031 7939
rect 5733 7905 5767 7939
rect 10701 7905 10735 7939
rect 11897 7905 11931 7939
rect 13185 7905 13219 7939
rect 13277 7905 13311 7939
rect 14749 7905 14783 7939
rect 14841 7905 14875 7939
rect 27077 7905 27111 7939
rect 30481 7905 30515 7939
rect 4629 7837 4663 7871
rect 7849 7837 7883 7871
rect 8953 7837 8987 7871
rect 10977 7837 11011 7871
rect 11345 7837 11379 7871
rect 11621 7837 11655 7871
rect 13093 7837 13127 7871
rect 13737 7837 13771 7871
rect 14657 7837 14691 7871
rect 19717 7837 19751 7871
rect 19993 7837 20027 7871
rect 23213 7837 23247 7871
rect 23489 7837 23523 7871
rect 23673 7837 23707 7871
rect 26801 7837 26835 7871
rect 26985 7837 27019 7871
rect 27169 7837 27203 7871
rect 27353 7837 27387 7871
rect 28825 7837 28859 7871
rect 28917 7837 28951 7871
rect 29561 7837 29595 7871
rect 29745 7837 29779 7871
rect 30205 7837 30239 7871
rect 30389 7837 30423 7871
rect 30573 7837 30607 7871
rect 30757 7837 30791 7871
rect 31033 7837 31067 7871
rect 31401 7837 31435 7871
rect 31493 7837 31527 7871
rect 31585 7837 31619 7871
rect 6009 7769 6043 7803
rect 9229 7769 9263 7803
rect 19901 7769 19935 7803
rect 29653 7769 29687 7803
rect 31769 7769 31803 7803
rect 12173 7701 12207 7735
rect 13553 7701 13587 7735
rect 23029 7701 23063 7735
rect 27537 7701 27571 7735
rect 30941 7701 30975 7735
rect 31309 7701 31343 7735
rect 4445 7497 4479 7531
rect 4905 7497 4939 7531
rect 5365 7497 5399 7531
rect 6377 7497 6411 7531
rect 9321 7497 9355 7531
rect 15301 7497 15335 7531
rect 17693 7497 17727 7531
rect 20545 7497 20579 7531
rect 26801 7497 26835 7531
rect 33701 7497 33735 7531
rect 13001 7429 13035 7463
rect 17233 7429 17267 7463
rect 19625 7429 19659 7463
rect 22937 7429 22971 7463
rect 24041 7429 24075 7463
rect 25053 7429 25087 7463
rect 25881 7429 25915 7463
rect 30757 7429 30791 7463
rect 1501 7361 1535 7395
rect 4353 7361 4387 7395
rect 5273 7361 5307 7395
rect 6561 7361 6595 7395
rect 9229 7361 9263 7395
rect 9413 7361 9447 7395
rect 11621 7361 11655 7395
rect 15393 7361 15427 7395
rect 17417 7361 17451 7395
rect 17509 7361 17543 7395
rect 17601 7361 17635 7395
rect 17785 7361 17819 7395
rect 19533 7361 19567 7395
rect 19717 7361 19751 7395
rect 19993 7361 20027 7395
rect 20177 7361 20211 7395
rect 20269 7361 20303 7395
rect 20361 7361 20395 7395
rect 20545 7361 20579 7395
rect 20821 7361 20855 7395
rect 22017 7361 22051 7395
rect 22109 7361 22143 7395
rect 22339 7361 22373 7395
rect 22477 7361 22511 7395
rect 22845 7361 22879 7395
rect 23949 7361 23983 7395
rect 24133 7361 24167 7395
rect 24225 7361 24259 7395
rect 24409 7361 24443 7395
rect 24593 7361 24627 7395
rect 24777 7361 24811 7395
rect 25513 7361 25547 7395
rect 25789 7361 25823 7395
rect 25973 7361 26007 7395
rect 26617 7351 26651 7385
rect 26801 7361 26835 7395
rect 27261 7361 27295 7395
rect 27353 7361 27387 7395
rect 27445 7361 27479 7395
rect 27629 7361 27663 7395
rect 28457 7361 28491 7395
rect 29193 7361 29227 7395
rect 29285 7361 29319 7395
rect 29561 7361 29595 7395
rect 29837 7361 29871 7395
rect 31401 7361 31435 7395
rect 31769 7361 31803 7395
rect 31953 7361 31987 7395
rect 33333 7361 33367 7395
rect 4629 7293 4663 7327
rect 5457 7293 5491 7327
rect 9597 7293 9631 7327
rect 9873 7293 9907 7327
rect 11345 7293 11379 7327
rect 12725 7293 12759 7327
rect 14749 7293 14783 7327
rect 15485 7293 15519 7327
rect 20913 7293 20947 7327
rect 21833 7293 21867 7327
rect 22753 7293 22787 7327
rect 24501 7293 24535 7327
rect 25421 7293 25455 7327
rect 26985 7293 27019 7327
rect 29101 7293 29135 7327
rect 31309 7293 31343 7327
rect 33241 7293 33275 7327
rect 1685 7225 1719 7259
rect 19809 7225 19843 7259
rect 21189 7225 21223 7259
rect 22569 7225 22603 7259
rect 3985 7157 4019 7191
rect 12173 7157 12207 7191
rect 14933 7157 14967 7191
rect 17233 7157 17267 7191
rect 22293 7157 22327 7191
rect 24961 7157 24995 7191
rect 25145 7157 25179 7191
rect 25697 7157 25731 7191
rect 11253 6953 11287 6987
rect 11529 6953 11563 6987
rect 17785 6953 17819 6987
rect 20085 6953 20119 6987
rect 25605 6953 25639 6987
rect 33149 6953 33183 6987
rect 17049 6885 17083 6919
rect 18153 6885 18187 6919
rect 21741 6885 21775 6919
rect 23673 6885 23707 6919
rect 28549 6885 28583 6919
rect 30941 6885 30975 6919
rect 3801 6817 3835 6851
rect 6193 6817 6227 6851
rect 8493 6817 8527 6851
rect 8585 6817 8619 6851
rect 11621 6817 11655 6851
rect 17509 6817 17543 6851
rect 17969 6817 18003 6851
rect 19257 6817 19291 6851
rect 25053 6817 25087 6851
rect 27445 6817 27479 6851
rect 30481 6817 30515 6851
rect 32505 6817 32539 6851
rect 32781 6817 32815 6851
rect 32873 6817 32907 6851
rect 3617 6749 3651 6783
rect 11253 6749 11287 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 12081 6749 12115 6783
rect 13185 6749 13219 6783
rect 15209 6749 15243 6783
rect 15301 6749 15335 6783
rect 17417 6739 17451 6773
rect 17601 6749 17635 6783
rect 17693 6749 17727 6783
rect 18061 6749 18095 6783
rect 18521 6749 18555 6783
rect 18613 6749 18647 6783
rect 18705 6749 18739 6783
rect 18889 6749 18923 6783
rect 19441 6749 19475 6783
rect 21557 6749 21591 6783
rect 21833 6749 21867 6783
rect 22201 6749 22235 6783
rect 22385 6749 22419 6783
rect 22477 6749 22511 6783
rect 22753 6749 22787 6783
rect 22845 6749 22879 6783
rect 25145 6749 25179 6783
rect 25605 6749 25639 6783
rect 25881 6749 25915 6783
rect 27169 6749 27203 6783
rect 27261 6749 27295 6783
rect 27721 6749 27755 6783
rect 27869 6749 27903 6783
rect 27997 6749 28031 6783
rect 28186 6749 28220 6783
rect 28733 6749 28767 6783
rect 28917 6749 28951 6783
rect 29009 6749 29043 6783
rect 30205 6749 30239 6783
rect 30665 6749 30699 6783
rect 31033 6749 31067 6783
rect 31125 6749 31159 6783
rect 32689 6749 32723 6783
rect 32965 6749 32999 6783
rect 33149 6749 33183 6783
rect 33333 6749 33367 6783
rect 33425 6749 33459 6783
rect 4077 6681 4111 6715
rect 6469 6681 6503 6715
rect 15577 6681 15611 6715
rect 18245 6681 18279 6715
rect 19625 6681 19659 6715
rect 19993 6681 20027 6715
rect 22017 6681 22051 6715
rect 23213 6681 23247 6715
rect 25789 6681 25823 6715
rect 27445 6681 27479 6715
rect 28089 6681 28123 6715
rect 3433 6613 3467 6647
rect 5549 6613 5583 6647
rect 7941 6613 7975 6647
rect 8033 6613 8067 6647
rect 8401 6613 8435 6647
rect 11897 6613 11931 6647
rect 12081 6613 12115 6647
rect 15025 6613 15059 6647
rect 21373 6613 21407 6647
rect 25513 6613 25547 6647
rect 28365 6613 28399 6647
rect 6837 6409 6871 6443
rect 9229 6409 9263 6443
rect 13185 6409 13219 6443
rect 18889 6409 18923 6443
rect 23121 6409 23155 6443
rect 24691 6409 24725 6443
rect 28181 6409 28215 6443
rect 31953 6409 31987 6443
rect 32137 6409 32171 6443
rect 11897 6341 11931 6375
rect 12265 6341 12299 6375
rect 12633 6341 12667 6375
rect 19073 6341 19107 6375
rect 24777 6341 24811 6375
rect 31585 6341 31619 6375
rect 31769 6341 31803 6375
rect 7021 6273 7055 6307
rect 7941 6273 7975 6307
rect 8125 6273 8159 6307
rect 8217 6273 8251 6307
rect 8585 6273 8619 6307
rect 9321 6273 9355 6307
rect 9505 6273 9539 6307
rect 9689 6273 9723 6307
rect 11621 6273 11655 6307
rect 13461 6273 13495 6307
rect 18245 6273 18279 6307
rect 18429 6273 18463 6307
rect 18521 6273 18555 6307
rect 18705 6273 18739 6307
rect 19257 6273 19291 6307
rect 22201 6273 22235 6307
rect 22385 6273 22419 6307
rect 22477 6273 22511 6307
rect 22625 6273 22659 6307
rect 22753 6273 22787 6307
rect 22845 6273 22879 6307
rect 22983 6273 23017 6307
rect 24593 6273 24627 6307
rect 24869 6273 24903 6307
rect 27813 6273 27847 6307
rect 27997 6273 28031 6307
rect 28089 6273 28123 6307
rect 30113 6273 30147 6307
rect 30297 6273 30331 6307
rect 32413 6273 32447 6307
rect 32505 6273 32539 6307
rect 32597 6273 32631 6307
rect 32781 6273 32815 6307
rect 8033 6205 8067 6239
rect 8493 6205 8527 6239
rect 13093 6205 13127 6239
rect 13645 6205 13679 6239
rect 8309 6137 8343 6171
rect 27813 6137 27847 6171
rect 30297 6137 30331 6171
rect 8401 6069 8435 6103
rect 9321 6069 9355 6103
rect 9781 6069 9815 6103
rect 18337 6069 18371 6103
rect 18705 6069 18739 6103
rect 19441 6069 19475 6103
rect 22293 6069 22327 6103
rect 12633 5865 12667 5899
rect 13093 5865 13127 5899
rect 20637 5865 20671 5899
rect 24225 5865 24259 5899
rect 27721 5865 27755 5899
rect 28365 5865 28399 5899
rect 30113 5865 30147 5899
rect 31125 5865 31159 5899
rect 32045 5865 32079 5899
rect 7665 5797 7699 5831
rect 9597 5797 9631 5831
rect 13369 5797 13403 5831
rect 15209 5797 15243 5831
rect 29929 5797 29963 5831
rect 30481 5797 30515 5831
rect 7757 5729 7791 5763
rect 8677 5729 8711 5763
rect 9689 5729 9723 5763
rect 13553 5729 13587 5763
rect 15761 5729 15795 5763
rect 19901 5729 19935 5763
rect 20177 5729 20211 5763
rect 22661 5729 22695 5763
rect 7481 5661 7515 5695
rect 8125 5661 8159 5695
rect 8953 5661 8987 5695
rect 9046 5661 9080 5695
rect 9321 5661 9355 5695
rect 9418 5661 9452 5695
rect 10425 5661 10459 5695
rect 12265 5661 12299 5695
rect 12449 5661 12483 5695
rect 13001 5661 13035 5695
rect 13185 5661 13219 5695
rect 13737 5661 13771 5695
rect 14657 5661 14691 5695
rect 15025 5661 15059 5695
rect 15301 5661 15335 5695
rect 19809 5661 19843 5695
rect 19993 5661 20027 5695
rect 20269 5661 20303 5695
rect 22569 5661 22603 5695
rect 22753 5661 22787 5695
rect 23213 5661 23247 5695
rect 23305 5661 23339 5695
rect 23673 5661 23707 5695
rect 23857 5661 23891 5695
rect 23949 5661 23983 5695
rect 24041 5661 24075 5695
rect 24869 5661 24903 5695
rect 25145 5661 25179 5695
rect 25329 5661 25363 5695
rect 27905 5661 27939 5695
rect 28089 5661 28123 5695
rect 28181 5661 28215 5695
rect 28273 5661 28307 5695
rect 28457 5661 28491 5695
rect 29653 5661 29687 5695
rect 30205 5661 30239 5695
rect 30941 5661 30975 5695
rect 31953 5661 31987 5695
rect 32137 5661 32171 5695
rect 9229 5593 9263 5627
rect 13921 5593 13955 5627
rect 14841 5593 14875 5627
rect 14933 5593 14967 5627
rect 15393 5593 15427 5627
rect 30757 5593 30791 5627
rect 7297 5525 7331 5559
rect 10333 5525 10367 5559
rect 11713 5525 11747 5559
rect 16405 5525 16439 5559
rect 22845 5525 22879 5559
rect 23489 5525 23523 5559
rect 24685 5525 24719 5559
rect 30665 5525 30699 5559
rect 8125 5321 8159 5355
rect 9413 5321 9447 5355
rect 12173 5321 12207 5355
rect 12449 5321 12483 5355
rect 13737 5321 13771 5355
rect 14473 5321 14507 5355
rect 16451 5321 16485 5355
rect 30113 5321 30147 5355
rect 31585 5321 31619 5355
rect 6653 5253 6687 5287
rect 9137 5253 9171 5287
rect 9781 5253 9815 5287
rect 19717 5253 19751 5287
rect 20821 5253 20855 5287
rect 21465 5253 21499 5287
rect 24317 5253 24351 5287
rect 6377 5185 6411 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 8677 5185 8711 5219
rect 8769 5185 8803 5219
rect 8917 5185 8951 5219
rect 9045 5185 9079 5219
rect 9275 5185 9309 5219
rect 9505 5185 9539 5219
rect 12265 5185 12299 5219
rect 12449 5185 12483 5219
rect 12725 5185 12759 5219
rect 13829 5185 13863 5219
rect 14381 5185 14415 5219
rect 14657 5185 14691 5219
rect 19349 5185 19383 5219
rect 19441 5185 19475 5219
rect 19901 5185 19935 5219
rect 20085 5185 20119 5219
rect 20269 5185 20303 5219
rect 20545 5185 20579 5219
rect 21281 5185 21315 5219
rect 22753 5185 22787 5219
rect 22937 5185 22971 5219
rect 23213 5185 23247 5219
rect 23765 5185 23799 5219
rect 23949 5185 23983 5219
rect 29653 5185 29687 5219
rect 29745 5185 29779 5219
rect 29929 5185 29963 5219
rect 30297 5185 30331 5219
rect 30573 5185 30607 5219
rect 30757 5185 30791 5219
rect 31217 5185 31251 5219
rect 11529 5117 11563 5151
rect 14013 5117 14047 5151
rect 15025 5117 15059 5151
rect 19809 5117 19843 5151
rect 20361 5117 20395 5151
rect 20913 5117 20947 5151
rect 22845 5117 22879 5151
rect 23029 5117 23063 5151
rect 29837 5117 29871 5151
rect 31125 5117 31159 5151
rect 30389 5049 30423 5083
rect 30481 5049 30515 5083
rect 8217 4981 8251 5015
rect 11253 4981 11287 5015
rect 13277 4981 13311 5015
rect 13369 4981 13403 5015
rect 19165 4981 19199 5015
rect 21649 4981 21683 5015
rect 29469 4981 29503 5015
rect 6732 4777 6766 4811
rect 9321 4777 9355 4811
rect 9762 4777 9796 4811
rect 13645 4777 13679 4811
rect 16589 4777 16623 4811
rect 19993 4777 20027 4811
rect 20361 4777 20395 4811
rect 20545 4777 20579 4811
rect 24593 4777 24627 4811
rect 26065 4777 26099 4811
rect 26433 4777 26467 4811
rect 30021 4777 30055 4811
rect 30297 4777 30331 4811
rect 30389 4777 30423 4811
rect 13737 4709 13771 4743
rect 15853 4709 15887 4743
rect 23949 4709 23983 4743
rect 27169 4709 27203 4743
rect 6469 4641 6503 4675
rect 9505 4641 9539 4675
rect 11897 4641 11931 4675
rect 14381 4641 14415 4675
rect 15945 4641 15979 4675
rect 19625 4641 19659 4675
rect 23305 4641 23339 4675
rect 24685 4641 24719 4675
rect 24777 4641 24811 4675
rect 26893 4641 26927 4675
rect 28549 4641 28583 4675
rect 29285 4641 29319 4675
rect 1501 4573 1535 4607
rect 8953 4573 8987 4607
rect 13921 4573 13955 4607
rect 14105 4573 14139 4607
rect 19257 4573 19291 4607
rect 19441 4573 19475 4607
rect 19717 4573 19751 4607
rect 22661 4573 22695 4607
rect 22937 4573 22971 4607
rect 24225 4573 24259 4607
rect 24409 4573 24443 4607
rect 24501 4573 24535 4607
rect 24961 4573 24995 4607
rect 25053 4573 25087 4607
rect 25145 4573 25179 4607
rect 25237 4573 25271 4607
rect 25605 4573 25639 4607
rect 25881 4573 25915 4607
rect 25973 4573 26007 4607
rect 26801 4573 26835 4607
rect 27629 4573 27663 4607
rect 28641 4573 28675 4607
rect 29837 4573 29871 4607
rect 30389 4573 30423 4607
rect 30573 4573 30607 4607
rect 9137 4505 9171 4539
rect 12173 4505 12207 4539
rect 20177 4505 20211 4539
rect 20377 4505 20411 4539
rect 23949 4505 23983 4539
rect 25421 4505 25455 4539
rect 27445 4505 27479 4539
rect 1593 4437 1627 4471
rect 8217 4437 8251 4471
rect 11253 4437 11287 4471
rect 19441 4437 19475 4471
rect 24133 4437 24167 4471
rect 25789 4437 25823 4471
rect 27813 4437 27847 4471
rect 9045 4233 9079 4267
rect 12633 4233 12667 4267
rect 13001 4233 13035 4267
rect 25421 4233 25455 4267
rect 25789 4233 25823 4267
rect 26341 4233 26375 4267
rect 26985 4233 27019 4267
rect 28549 4233 28583 4267
rect 26709 4165 26743 4199
rect 27813 4165 27847 4199
rect 8401 4097 8435 4131
rect 12817 4097 12851 4131
rect 13090 4119 13124 4153
rect 21925 4097 21959 4131
rect 22477 4097 22511 4131
rect 25329 4097 25363 4131
rect 25507 4097 25541 4131
rect 25605 4097 25639 4131
rect 25797 4087 25831 4121
rect 26065 4097 26099 4131
rect 26617 4097 26651 4131
rect 26801 4097 26835 4131
rect 27353 4097 27387 4131
rect 27629 4097 27663 4131
rect 27997 4097 28031 4131
rect 28089 4097 28123 4131
rect 28457 4097 28491 4131
rect 28641 4097 28675 4131
rect 26341 4029 26375 4063
rect 27445 4029 27479 4063
rect 26157 3893 26191 3927
rect 27813 3893 27847 3927
rect 11805 3009 11839 3043
rect 13185 3009 13219 3043
rect 16405 3009 16439 3043
rect 17601 3009 17635 3043
rect 24593 3009 24627 3043
rect 37105 3009 37139 3043
rect 37565 3009 37599 3043
rect 36921 2873 36955 2907
rect 11621 2805 11655 2839
rect 13001 2805 13035 2839
rect 16221 2805 16255 2839
rect 17417 2805 17451 2839
rect 24409 2805 24443 2839
rect 37657 2805 37691 2839
rect 8677 2601 8711 2635
rect 11253 2601 11287 2635
rect 37657 2533 37691 2567
rect 1501 2397 1535 2431
rect 2145 2397 2179 2431
rect 4077 2397 4111 2431
rect 6653 2397 6687 2431
rect 8493 2397 8527 2431
rect 13093 2397 13127 2431
rect 15025 2397 15059 2431
rect 17601 2397 17635 2431
rect 19533 2397 19567 2431
rect 37473 2397 37507 2431
rect 11161 2329 11195 2363
rect 27077 2329 27111 2363
rect 1593 2261 1627 2295
rect 2237 2261 2271 2295
rect 4169 2261 4203 2295
rect 6929 2261 6963 2295
rect 13185 2261 13219 2295
rect 15301 2261 15335 2295
rect 17693 2261 17727 2295
rect 19625 2261 19659 2295
rect 27169 2261 27203 2295
<< metal1 >>
rect 1104 39194 38272 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38272 39194
rect 1104 39120 38272 39142
rect 14 39040 20 39092
rect 72 39080 78 39092
rect 1581 39083 1639 39089
rect 1581 39080 1593 39083
rect 72 39052 1593 39080
rect 72 39040 78 39052
rect 1581 39049 1593 39052
rect 1627 39049 1639 39083
rect 1581 39043 1639 39049
rect 4522 39040 4528 39092
rect 4580 39080 4586 39092
rect 4985 39083 5043 39089
rect 4985 39080 4997 39083
rect 4580 39052 4997 39080
rect 4580 39040 4586 39052
rect 4985 39049 4997 39052
rect 5031 39049 5043 39083
rect 4985 39043 5043 39049
rect 9030 39040 9036 39092
rect 9088 39080 9094 39092
rect 9493 39083 9551 39089
rect 9493 39080 9505 39083
rect 9088 39052 9505 39080
rect 9088 39040 9094 39052
rect 9493 39049 9505 39052
rect 9539 39049 9551 39083
rect 9493 39043 9551 39049
rect 11054 39040 11060 39092
rect 11112 39080 11118 39092
rect 11701 39083 11759 39089
rect 11701 39080 11713 39083
rect 11112 39052 11713 39080
rect 11112 39040 11118 39052
rect 11701 39049 11713 39052
rect 11747 39049 11759 39083
rect 11701 39043 11759 39049
rect 12894 39040 12900 39092
rect 12952 39080 12958 39092
rect 13173 39083 13231 39089
rect 13173 39080 13185 39083
rect 12952 39052 13185 39080
rect 12952 39040 12958 39052
rect 13173 39049 13185 39052
rect 13219 39049 13231 39083
rect 13173 39043 13231 39049
rect 14476 39052 16068 39080
rect 9122 38972 9128 39024
rect 9180 39012 9186 39024
rect 14476 39012 14504 39052
rect 16040 39024 16068 39052
rect 17402 39040 17408 39092
rect 17460 39080 17466 39092
rect 17865 39083 17923 39089
rect 17865 39080 17877 39083
rect 17460 39052 17877 39080
rect 17460 39040 17466 39052
rect 17865 39049 17877 39052
rect 17911 39049 17923 39083
rect 17865 39043 17923 39049
rect 21910 39040 21916 39092
rect 21968 39080 21974 39092
rect 22189 39083 22247 39089
rect 22189 39080 22201 39083
rect 21968 39052 22201 39080
rect 21968 39040 21974 39052
rect 22189 39049 22201 39052
rect 22235 39049 22247 39083
rect 22189 39043 22247 39049
rect 26418 39040 26424 39092
rect 26476 39080 26482 39092
rect 27157 39083 27215 39089
rect 27157 39080 27169 39083
rect 26476 39052 27169 39080
rect 26476 39040 26482 39052
rect 27157 39049 27169 39052
rect 27203 39049 27215 39083
rect 27157 39043 27215 39049
rect 32858 39040 32864 39092
rect 32916 39080 32922 39092
rect 33137 39083 33195 39089
rect 33137 39080 33149 39083
rect 32916 39052 33149 39080
rect 32916 39040 32922 39052
rect 33137 39049 33149 39052
rect 33183 39049 33195 39083
rect 33137 39043 33195 39049
rect 9180 38984 14504 39012
rect 9180 38972 9186 38984
rect 15470 38972 15476 39024
rect 15528 39012 15534 39024
rect 15657 39015 15715 39021
rect 15657 39012 15669 39015
rect 15528 38984 15669 39012
rect 15528 38972 15534 38984
rect 15657 38981 15669 38984
rect 15703 38981 15715 39015
rect 15657 38975 15715 38981
rect 16022 38972 16028 39024
rect 16080 38972 16086 39024
rect 24394 39012 24400 39024
rect 17696 38984 24400 39012
rect 1489 38947 1547 38953
rect 1489 38913 1501 38947
rect 1535 38944 1547 38947
rect 3786 38944 3792 38956
rect 1535 38916 3792 38944
rect 1535 38913 1547 38916
rect 1489 38907 1547 38913
rect 3786 38904 3792 38916
rect 3844 38904 3850 38956
rect 4798 38904 4804 38956
rect 4856 38904 4862 38956
rect 9306 38904 9312 38956
rect 9364 38904 9370 38956
rect 11606 38904 11612 38956
rect 11664 38904 11670 38956
rect 11974 38904 11980 38956
rect 12032 38944 12038 38956
rect 12253 38947 12311 38953
rect 12253 38944 12265 38947
rect 12032 38916 12265 38944
rect 12032 38904 12038 38916
rect 12253 38913 12265 38916
rect 12299 38913 12311 38947
rect 12253 38907 12311 38913
rect 12710 38904 12716 38956
rect 12768 38904 12774 38956
rect 12986 38904 12992 38956
rect 13044 38904 13050 38956
rect 17696 38953 17724 38984
rect 24394 38972 24400 38984
rect 24452 38972 24458 39024
rect 30926 38972 30932 39024
rect 30984 39012 30990 39024
rect 31113 39015 31171 39021
rect 31113 39012 31125 39015
rect 30984 38984 31125 39012
rect 30984 38972 30990 38984
rect 31113 38981 31125 38984
rect 31159 38981 31171 39015
rect 31113 38975 31171 38981
rect 35894 38972 35900 39024
rect 35952 39012 35958 39024
rect 35989 39015 36047 39021
rect 35989 39012 36001 39015
rect 35952 38984 36001 39012
rect 35952 38972 35958 38984
rect 35989 38981 36001 38984
rect 36035 38981 36047 39015
rect 35989 38975 36047 38981
rect 17681 38947 17739 38953
rect 17681 38913 17693 38947
rect 17727 38913 17739 38947
rect 17681 38907 17739 38913
rect 19978 38904 19984 38956
rect 20036 38944 20042 38956
rect 20073 38947 20131 38953
rect 20073 38944 20085 38947
rect 20036 38916 20085 38944
rect 20036 38904 20042 38916
rect 20073 38913 20085 38916
rect 20119 38913 20131 38947
rect 20073 38907 20131 38913
rect 22094 38904 22100 38956
rect 22152 38904 22158 38956
rect 24762 38904 24768 38956
rect 24820 38904 24826 38956
rect 25038 38904 25044 38956
rect 25096 38944 25102 38956
rect 25869 38947 25927 38953
rect 25869 38944 25881 38947
rect 25096 38916 25881 38944
rect 25096 38904 25102 38916
rect 25869 38913 25881 38916
rect 25915 38913 25927 38947
rect 25869 38907 25927 38913
rect 27062 38904 27068 38956
rect 27120 38904 27126 38956
rect 33042 38904 33048 38956
rect 33100 38904 33106 38956
rect 35618 38904 35624 38956
rect 35676 38904 35682 38956
rect 37366 38904 37372 38956
rect 37424 38944 37430 38956
rect 37461 38947 37519 38953
rect 37461 38944 37473 38947
rect 37424 38916 37473 38944
rect 37424 38904 37430 38916
rect 37461 38913 37473 38916
rect 37507 38913 37519 38947
rect 37461 38907 37519 38913
rect 11238 38836 11244 38888
rect 11296 38876 11302 38888
rect 20349 38879 20407 38885
rect 20349 38876 20361 38879
rect 11296 38848 20361 38876
rect 11296 38836 11302 38848
rect 20349 38845 20361 38848
rect 20395 38845 20407 38879
rect 20349 38839 20407 38845
rect 26142 38836 26148 38888
rect 26200 38836 26206 38888
rect 10226 38768 10232 38820
rect 10284 38808 10290 38820
rect 10284 38780 15792 38808
rect 10284 38768 10290 38780
rect 12342 38700 12348 38752
rect 12400 38700 12406 38752
rect 12434 38700 12440 38752
rect 12492 38740 12498 38752
rect 15764 38749 15792 38780
rect 16022 38768 16028 38820
rect 16080 38808 16086 38820
rect 37645 38811 37703 38817
rect 37645 38808 37657 38811
rect 16080 38780 37657 38808
rect 16080 38768 16086 38780
rect 37645 38777 37657 38780
rect 37691 38777 37703 38811
rect 37645 38771 37703 38777
rect 12529 38743 12587 38749
rect 12529 38740 12541 38743
rect 12492 38712 12541 38740
rect 12492 38700 12498 38712
rect 12529 38709 12541 38712
rect 12575 38709 12587 38743
rect 12529 38703 12587 38709
rect 15749 38743 15807 38749
rect 15749 38709 15761 38743
rect 15795 38709 15807 38743
rect 15749 38703 15807 38709
rect 24857 38743 24915 38749
rect 24857 38709 24869 38743
rect 24903 38740 24915 38743
rect 24946 38740 24952 38752
rect 24903 38712 24952 38740
rect 24903 38709 24915 38712
rect 24857 38703 24915 38709
rect 24946 38700 24952 38712
rect 25004 38700 25010 38752
rect 31202 38700 31208 38752
rect 31260 38700 31266 38752
rect 1104 38650 38272 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38272 38650
rect 1104 38576 38272 38598
rect 4798 38496 4804 38548
rect 4856 38536 4862 38548
rect 4985 38539 5043 38545
rect 4985 38536 4997 38539
rect 4856 38508 4997 38536
rect 4856 38496 4862 38508
rect 4985 38505 4997 38508
rect 5031 38505 5043 38539
rect 4985 38499 5043 38505
rect 9306 38496 9312 38548
rect 9364 38496 9370 38548
rect 12332 38539 12390 38545
rect 12332 38505 12344 38539
rect 12378 38536 12390 38539
rect 12434 38536 12440 38548
rect 12378 38508 12440 38536
rect 12378 38505 12390 38508
rect 12332 38499 12390 38505
rect 12434 38496 12440 38508
rect 12492 38496 12498 38548
rect 17494 38496 17500 38548
rect 17552 38536 17558 38548
rect 22646 38536 22652 38548
rect 17552 38508 22652 38536
rect 17552 38496 17558 38508
rect 22646 38496 22652 38508
rect 22704 38496 22710 38548
rect 24394 38496 24400 38548
rect 24452 38496 24458 38548
rect 25038 38536 25044 38548
rect 24504 38508 25044 38536
rect 12069 38403 12127 38409
rect 12069 38369 12081 38403
rect 12115 38400 12127 38403
rect 12342 38400 12348 38412
rect 12115 38372 12348 38400
rect 12115 38369 12127 38372
rect 12069 38363 12127 38369
rect 12342 38360 12348 38372
rect 12400 38360 12406 38412
rect 14458 38360 14464 38412
rect 14516 38400 14522 38412
rect 20898 38400 20904 38412
rect 14516 38372 20904 38400
rect 14516 38360 14522 38372
rect 20898 38360 20904 38372
rect 20956 38360 20962 38412
rect 22741 38403 22799 38409
rect 22741 38400 22753 38403
rect 21928 38372 22753 38400
rect 5166 38292 5172 38344
rect 5224 38292 5230 38344
rect 8481 38335 8539 38341
rect 8481 38332 8493 38335
rect 7116 38304 8493 38332
rect 7116 38208 7144 38304
rect 8481 38301 8493 38304
rect 8527 38301 8539 38335
rect 8481 38295 8539 38301
rect 8496 38264 8524 38295
rect 9490 38292 9496 38344
rect 9548 38292 9554 38344
rect 9861 38335 9919 38341
rect 9861 38332 9873 38335
rect 9646 38304 9873 38332
rect 9646 38264 9674 38304
rect 9861 38301 9873 38304
rect 9907 38301 9919 38335
rect 9861 38295 9919 38301
rect 9953 38335 10011 38341
rect 9953 38301 9965 38335
rect 9999 38332 10011 38335
rect 10137 38335 10195 38341
rect 10137 38332 10149 38335
rect 9999 38304 10149 38332
rect 9999 38301 10011 38304
rect 9953 38295 10011 38301
rect 10137 38301 10149 38304
rect 10183 38301 10195 38335
rect 10137 38295 10195 38301
rect 20162 38292 20168 38344
rect 20220 38292 20226 38344
rect 20257 38335 20315 38341
rect 20257 38301 20269 38335
rect 20303 38301 20315 38335
rect 20257 38295 20315 38301
rect 20349 38335 20407 38341
rect 20349 38301 20361 38335
rect 20395 38332 20407 38335
rect 20533 38335 20591 38341
rect 20533 38332 20545 38335
rect 20395 38304 20545 38332
rect 20395 38301 20407 38304
rect 20349 38295 20407 38301
rect 20533 38301 20545 38304
rect 20579 38301 20591 38335
rect 21928 38318 21956 38372
rect 22741 38369 22753 38372
rect 22787 38400 22799 38403
rect 24394 38400 24400 38412
rect 22787 38372 24400 38400
rect 22787 38369 22799 38372
rect 22741 38363 22799 38369
rect 24394 38360 24400 38372
rect 24452 38360 24458 38412
rect 20533 38295 20591 38301
rect 8496 38236 9674 38264
rect 10410 38224 10416 38276
rect 10468 38224 10474 38276
rect 13998 38264 14004 38276
rect 11638 38236 12834 38264
rect 13648 38236 14004 38264
rect 7098 38156 7104 38208
rect 7156 38156 7162 38208
rect 8570 38156 8576 38208
rect 8628 38156 8634 38208
rect 10594 38156 10600 38208
rect 10652 38196 10658 38208
rect 11716 38196 11744 38236
rect 10652 38168 11744 38196
rect 10652 38156 10658 38168
rect 11882 38156 11888 38208
rect 11940 38156 11946 38208
rect 11974 38156 11980 38208
rect 12032 38196 12038 38208
rect 13648 38196 13676 38236
rect 13998 38224 14004 38236
rect 14056 38264 14062 38276
rect 20272 38264 20300 38295
rect 22554 38292 22560 38344
rect 22612 38332 22618 38344
rect 24504 38332 24532 38508
rect 25038 38496 25044 38508
rect 25096 38496 25102 38548
rect 27890 38536 27896 38548
rect 27080 38508 27896 38536
rect 24673 38403 24731 38409
rect 24673 38369 24685 38403
rect 24719 38400 24731 38403
rect 24946 38400 24952 38412
rect 24719 38372 24952 38400
rect 24719 38369 24731 38372
rect 24673 38363 24731 38369
rect 24946 38360 24952 38372
rect 25004 38360 25010 38412
rect 26142 38360 26148 38412
rect 26200 38400 26206 38412
rect 27080 38400 27108 38508
rect 27890 38496 27896 38508
rect 27948 38536 27954 38548
rect 30282 38536 30288 38548
rect 27948 38508 30288 38536
rect 27948 38496 27954 38508
rect 30282 38496 30288 38508
rect 30340 38496 30346 38548
rect 32125 38539 32183 38545
rect 32125 38505 32137 38539
rect 32171 38536 32183 38539
rect 33042 38536 33048 38548
rect 32171 38508 33048 38536
rect 32171 38505 32183 38508
rect 32125 38499 32183 38505
rect 33042 38496 33048 38508
rect 33100 38496 33106 38548
rect 34701 38539 34759 38545
rect 34701 38505 34713 38539
rect 34747 38536 34759 38539
rect 35618 38536 35624 38548
rect 34747 38508 35624 38536
rect 34747 38505 34759 38508
rect 34701 38499 34759 38505
rect 35618 38496 35624 38508
rect 35676 38496 35682 38548
rect 37829 38539 37887 38545
rect 37829 38505 37841 38539
rect 37875 38536 37887 38539
rect 37918 38536 37924 38548
rect 37875 38508 37924 38536
rect 37875 38505 37887 38508
rect 37829 38499 37887 38505
rect 37918 38496 37924 38508
rect 37976 38496 37982 38548
rect 27338 38400 27344 38412
rect 26200 38372 27344 38400
rect 26200 38360 26206 38372
rect 27338 38360 27344 38372
rect 27396 38360 27402 38412
rect 27614 38360 27620 38412
rect 27672 38400 27678 38412
rect 28721 38403 28779 38409
rect 28721 38400 28733 38403
rect 27672 38372 28733 38400
rect 27672 38360 27678 38372
rect 28721 38369 28733 38372
rect 28767 38369 28779 38403
rect 28721 38363 28779 38369
rect 29196 38372 31892 38400
rect 22612 38304 24532 38332
rect 24581 38335 24639 38341
rect 22612 38292 22618 38304
rect 24581 38301 24593 38335
rect 24627 38301 24639 38335
rect 26160 38332 26188 38360
rect 29196 38341 29224 38372
rect 26082 38304 26188 38332
rect 26697 38335 26755 38341
rect 24581 38295 24639 38301
rect 26697 38301 26709 38335
rect 26743 38301 26755 38335
rect 26697 38295 26755 38301
rect 26789 38335 26847 38341
rect 26789 38301 26801 38335
rect 26835 38332 26847 38335
rect 26973 38335 27031 38341
rect 26973 38332 26985 38335
rect 26835 38304 26985 38332
rect 26835 38301 26847 38304
rect 26789 38295 26847 38301
rect 26973 38301 26985 38304
rect 27019 38301 27031 38335
rect 26973 38295 27031 38301
rect 29181 38335 29239 38341
rect 29181 38301 29193 38335
rect 29227 38301 29239 38335
rect 29181 38295 29239 38301
rect 29273 38335 29331 38341
rect 29273 38301 29285 38335
rect 29319 38332 29331 38335
rect 29549 38335 29607 38341
rect 29549 38332 29561 38335
rect 29319 38304 29561 38332
rect 29319 38301 29331 38304
rect 29273 38295 29331 38301
rect 29549 38301 29561 38304
rect 29595 38301 29607 38335
rect 29549 38295 29607 38301
rect 14056 38236 20300 38264
rect 20809 38267 20867 38273
rect 14056 38224 14062 38236
rect 20809 38233 20821 38267
rect 20855 38233 20867 38267
rect 24596 38264 24624 38295
rect 24854 38264 24860 38276
rect 24596 38236 24860 38264
rect 20809 38227 20867 38233
rect 12032 38168 13676 38196
rect 12032 38156 12038 38168
rect 13722 38156 13728 38208
rect 13780 38196 13786 38208
rect 13817 38199 13875 38205
rect 13817 38196 13829 38199
rect 13780 38168 13829 38196
rect 13780 38156 13786 38168
rect 13817 38165 13829 38168
rect 13863 38196 13875 38199
rect 16206 38196 16212 38208
rect 13863 38168 16212 38196
rect 13863 38165 13875 38168
rect 13817 38159 13875 38165
rect 16206 38156 16212 38168
rect 16264 38156 16270 38208
rect 18690 38156 18696 38208
rect 18748 38196 18754 38208
rect 19886 38196 19892 38208
rect 18748 38168 19892 38196
rect 18748 38156 18754 38168
rect 19886 38156 19892 38168
rect 19944 38156 19950 38208
rect 19981 38199 20039 38205
rect 19981 38165 19993 38199
rect 20027 38196 20039 38199
rect 20824 38196 20852 38227
rect 24854 38224 24860 38236
rect 24912 38224 24918 38276
rect 24946 38224 24952 38276
rect 25004 38224 25010 38276
rect 26712 38264 26740 38295
rect 26252 38236 26740 38264
rect 20027 38168 20852 38196
rect 20027 38165 20039 38168
rect 19981 38159 20039 38165
rect 22278 38156 22284 38208
rect 22336 38156 22342 38208
rect 24762 38156 24768 38208
rect 24820 38196 24826 38208
rect 26252 38196 26280 38236
rect 24820 38168 26280 38196
rect 24820 38156 24826 38168
rect 26418 38156 26424 38208
rect 26476 38156 26482 38208
rect 26712 38196 26740 38236
rect 27246 38224 27252 38276
rect 27304 38224 27310 38276
rect 27338 38224 27344 38276
rect 27396 38264 27402 38276
rect 27396 38236 27738 38264
rect 27396 38224 27402 38236
rect 27614 38196 27620 38208
rect 26712 38168 27620 38196
rect 27614 38156 27620 38168
rect 27672 38196 27678 38208
rect 29196 38196 29224 38295
rect 31202 38292 31208 38344
rect 31260 38332 31266 38344
rect 31864 38341 31892 38372
rect 31849 38335 31907 38341
rect 31260 38304 31800 38332
rect 31260 38292 31266 38304
rect 29822 38224 29828 38276
rect 29880 38224 29886 38276
rect 30282 38224 30288 38276
rect 30340 38224 30346 38276
rect 31772 38264 31800 38304
rect 31849 38301 31861 38335
rect 31895 38301 31907 38335
rect 31849 38295 31907 38301
rect 32030 38292 32036 38344
rect 32088 38332 32094 38344
rect 32309 38335 32367 38341
rect 32309 38332 32321 38335
rect 32088 38304 32321 38332
rect 32088 38292 32094 38304
rect 32309 38301 32321 38304
rect 32355 38301 32367 38335
rect 32309 38295 32367 38301
rect 34514 38292 34520 38344
rect 34572 38332 34578 38344
rect 34885 38335 34943 38341
rect 34885 38332 34897 38335
rect 34572 38304 34897 38332
rect 34572 38292 34578 38304
rect 34885 38301 34897 38304
rect 34931 38301 34943 38335
rect 34885 38295 34943 38301
rect 37553 38267 37611 38273
rect 37553 38264 37565 38267
rect 31772 38236 37565 38264
rect 37553 38233 37565 38236
rect 37599 38233 37611 38267
rect 37553 38227 37611 38233
rect 27672 38168 29224 38196
rect 27672 38156 27678 38168
rect 29270 38156 29276 38208
rect 29328 38196 29334 38208
rect 31297 38199 31355 38205
rect 31297 38196 31309 38199
rect 29328 38168 31309 38196
rect 29328 38156 29334 38168
rect 31297 38165 31309 38168
rect 31343 38165 31355 38199
rect 31297 38159 31355 38165
rect 31938 38156 31944 38208
rect 31996 38156 32002 38208
rect 1104 38106 38272 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38272 38106
rect 1104 38032 38272 38054
rect 8570 37952 8576 38004
rect 8628 37952 8634 38004
rect 10321 37995 10379 38001
rect 10321 37961 10333 37995
rect 10367 37992 10379 37995
rect 10410 37992 10416 38004
rect 10367 37964 10416 37992
rect 10367 37961 10379 37964
rect 10321 37955 10379 37961
rect 10410 37952 10416 37964
rect 10468 37952 10474 38004
rect 10778 37952 10784 38004
rect 10836 37992 10842 38004
rect 11057 37995 11115 38001
rect 11057 37992 11069 37995
rect 10836 37964 11069 37992
rect 10836 37952 10842 37964
rect 11057 37961 11069 37964
rect 11103 37992 11115 37995
rect 11517 37995 11575 38001
rect 11103 37964 11284 37992
rect 11103 37961 11115 37964
rect 11057 37955 11115 37961
rect 8588 37924 8616 37952
rect 10594 37924 10600 37936
rect 8404 37896 8616 37924
rect 9890 37896 10600 37924
rect 8404 37865 8432 37896
rect 10594 37884 10600 37896
rect 10652 37884 10658 37936
rect 8389 37859 8447 37865
rect 8389 37825 8401 37859
rect 8435 37825 8447 37859
rect 8389 37819 8447 37825
rect 10505 37859 10563 37865
rect 10505 37825 10517 37859
rect 10551 37856 10563 37859
rect 10965 37859 11023 37865
rect 10551 37828 10640 37856
rect 10551 37825 10563 37828
rect 10505 37819 10563 37825
rect 8662 37748 8668 37800
rect 8720 37748 8726 37800
rect 10612 37729 10640 37828
rect 10965 37825 10977 37859
rect 11011 37825 11023 37859
rect 10965 37819 11023 37825
rect 10597 37723 10655 37729
rect 10597 37689 10609 37723
rect 10643 37689 10655 37723
rect 10980 37720 11008 37819
rect 11146 37748 11152 37800
rect 11204 37748 11210 37800
rect 11256 37788 11284 37964
rect 11517 37961 11529 37995
rect 11563 37992 11575 37995
rect 11606 37992 11612 38004
rect 11563 37964 11612 37992
rect 11563 37961 11575 37964
rect 11517 37955 11575 37961
rect 11606 37952 11612 37964
rect 11664 37952 11670 38004
rect 12253 37995 12311 38001
rect 12253 37961 12265 37995
rect 12299 37992 12311 37995
rect 12710 37992 12716 38004
rect 12299 37964 12716 37992
rect 12299 37961 12311 37964
rect 12253 37955 12311 37961
rect 12710 37952 12716 37964
rect 12768 37952 12774 38004
rect 13722 37952 13728 38004
rect 13780 37952 13786 38004
rect 14458 37992 14464 38004
rect 13832 37964 14464 37992
rect 12621 37927 12679 37933
rect 12621 37893 12633 37927
rect 12667 37924 12679 37927
rect 13078 37924 13084 37936
rect 12667 37896 13084 37924
rect 12667 37893 12679 37896
rect 12621 37887 12679 37893
rect 13078 37884 13084 37896
rect 13136 37924 13142 37936
rect 13740 37924 13768 37952
rect 13136 37896 13768 37924
rect 13136 37884 13142 37896
rect 11698 37816 11704 37868
rect 11756 37816 11762 37868
rect 12713 37791 12771 37797
rect 12713 37788 12725 37791
rect 11256 37760 12725 37788
rect 12713 37757 12725 37760
rect 12759 37757 12771 37791
rect 12713 37751 12771 37757
rect 12897 37791 12955 37797
rect 12897 37757 12909 37791
rect 12943 37788 12955 37791
rect 13832 37788 13860 37964
rect 14458 37952 14464 37964
rect 14516 37952 14522 38004
rect 14550 37952 14556 38004
rect 14608 37992 14614 38004
rect 14645 37995 14703 38001
rect 14645 37992 14657 37995
rect 14608 37964 14657 37992
rect 14608 37952 14614 37964
rect 14645 37961 14657 37964
rect 14691 37961 14703 37995
rect 17678 37992 17684 38004
rect 14645 37955 14703 37961
rect 17420 37964 17684 37992
rect 14568 37924 14596 37952
rect 17420 37924 17448 37964
rect 14108 37896 14596 37924
rect 14660 37896 17448 37924
rect 14108 37865 14136 37896
rect 14093 37859 14151 37865
rect 14093 37825 14105 37859
rect 14139 37825 14151 37859
rect 14093 37819 14151 37825
rect 14274 37816 14280 37868
rect 14332 37816 14338 37868
rect 14366 37816 14372 37868
rect 14424 37856 14430 37868
rect 14553 37859 14611 37865
rect 14553 37856 14565 37859
rect 14424 37828 14565 37856
rect 14424 37816 14430 37828
rect 14553 37825 14565 37828
rect 14599 37825 14611 37859
rect 14553 37819 14611 37825
rect 12943 37760 13860 37788
rect 13909 37791 13967 37797
rect 12943 37757 12955 37760
rect 12897 37751 12955 37757
rect 13909 37757 13921 37791
rect 13955 37788 13967 37791
rect 14384 37788 14412 37816
rect 13955 37760 14412 37788
rect 13955 37757 13967 37760
rect 13909 37751 13967 37757
rect 11882 37720 11888 37732
rect 10980 37692 11888 37720
rect 10597 37683 10655 37689
rect 11882 37680 11888 37692
rect 11940 37720 11946 37732
rect 12342 37720 12348 37732
rect 11940 37692 12348 37720
rect 11940 37680 11946 37692
rect 12342 37680 12348 37692
rect 12400 37720 12406 37732
rect 14369 37723 14427 37729
rect 14369 37720 14381 37723
rect 12400 37692 14381 37720
rect 12400 37680 12406 37692
rect 14369 37689 14381 37692
rect 14415 37720 14427 37723
rect 14660 37720 14688 37896
rect 17494 37884 17500 37936
rect 17552 37884 17558 37936
rect 17604 37933 17632 37964
rect 17678 37952 17684 37964
rect 17736 37952 17742 38004
rect 17862 37952 17868 38004
rect 17920 37952 17926 38004
rect 18690 37992 18696 38004
rect 18248 37964 18696 37992
rect 18248 37933 18276 37964
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 18782 37952 18788 38004
rect 18840 37992 18846 38004
rect 18840 37964 19472 37992
rect 18840 37952 18846 37964
rect 17589 37927 17647 37933
rect 17589 37893 17601 37927
rect 17635 37893 17647 37927
rect 18233 37927 18291 37933
rect 17589 37887 17647 37893
rect 17696 37896 18184 37924
rect 14737 37859 14795 37865
rect 14737 37825 14749 37859
rect 14783 37856 14795 37859
rect 14826 37856 14832 37868
rect 14783 37828 14832 37856
rect 14783 37825 14795 37828
rect 14737 37819 14795 37825
rect 14826 37816 14832 37828
rect 14884 37816 14890 37868
rect 14921 37859 14979 37865
rect 14921 37825 14933 37859
rect 14967 37856 14979 37859
rect 15565 37859 15623 37865
rect 15565 37856 15577 37859
rect 14967 37828 15577 37856
rect 14967 37825 14979 37828
rect 14921 37819 14979 37825
rect 15565 37825 15577 37828
rect 15611 37825 15623 37859
rect 15565 37819 15623 37825
rect 15657 37859 15715 37865
rect 15657 37825 15669 37859
rect 15703 37825 15715 37859
rect 15657 37819 15715 37825
rect 14415 37692 14688 37720
rect 15672 37720 15700 37819
rect 15746 37816 15752 37868
rect 15804 37856 15810 37868
rect 15841 37859 15899 37865
rect 15841 37856 15853 37859
rect 15804 37828 15853 37856
rect 15804 37816 15810 37828
rect 15841 37825 15853 37828
rect 15887 37825 15899 37859
rect 15841 37819 15899 37825
rect 15930 37816 15936 37868
rect 15988 37816 15994 37868
rect 16022 37816 16028 37868
rect 16080 37816 16086 37868
rect 17696 37865 17724 37896
rect 18156 37868 18184 37896
rect 18233 37893 18245 37927
rect 18279 37893 18291 37927
rect 18233 37887 18291 37893
rect 18601 37927 18659 37933
rect 18601 37893 18613 37927
rect 18647 37924 18659 37927
rect 18969 37927 19027 37933
rect 18969 37924 18981 37927
rect 18647 37896 18981 37924
rect 18647 37893 18659 37896
rect 18601 37887 18659 37893
rect 18969 37893 18981 37896
rect 19015 37893 19027 37927
rect 18969 37887 19027 37893
rect 17313 37859 17371 37865
rect 17313 37825 17325 37859
rect 17359 37825 17371 37859
rect 17313 37819 17371 37825
rect 17681 37859 17739 37865
rect 17681 37825 17693 37859
rect 17727 37825 17739 37859
rect 17681 37819 17739 37825
rect 17328 37720 17356 37819
rect 18138 37816 18144 37868
rect 18196 37816 18202 37868
rect 18417 37859 18475 37865
rect 18417 37825 18429 37859
rect 18463 37856 18475 37859
rect 18506 37856 18512 37868
rect 18463 37828 18512 37856
rect 18463 37825 18475 37828
rect 18417 37819 18475 37825
rect 18506 37816 18512 37828
rect 18564 37816 18570 37868
rect 18785 37859 18843 37865
rect 18785 37825 18797 37859
rect 18831 37856 18843 37859
rect 18874 37856 18880 37868
rect 18831 37828 18880 37856
rect 18831 37825 18843 37828
rect 18785 37819 18843 37825
rect 18874 37816 18880 37828
rect 18932 37816 18938 37868
rect 19058 37816 19064 37868
rect 19116 37816 19122 37868
rect 19150 37816 19156 37868
rect 19208 37816 19214 37868
rect 19444 37865 19472 37964
rect 20162 37952 20168 38004
rect 20220 37992 20226 38004
rect 20441 37995 20499 38001
rect 20441 37992 20453 37995
rect 20220 37964 20453 37992
rect 20220 37952 20226 37964
rect 20441 37961 20453 37964
rect 20487 37961 20499 37995
rect 20441 37955 20499 37961
rect 22097 37995 22155 38001
rect 22097 37961 22109 37995
rect 22143 37992 22155 37995
rect 22186 37992 22192 38004
rect 22143 37964 22192 37992
rect 22143 37961 22155 37964
rect 22097 37955 22155 37961
rect 22186 37952 22192 37964
rect 22244 37952 22250 38004
rect 22646 37952 22652 38004
rect 22704 37992 22710 38004
rect 23934 37992 23940 38004
rect 22704 37964 23940 37992
rect 22704 37952 22710 37964
rect 23934 37952 23940 37964
rect 23992 37952 23998 38004
rect 24946 37952 24952 38004
rect 25004 37992 25010 38004
rect 25501 37995 25559 38001
rect 25501 37992 25513 37995
rect 25004 37964 25513 37992
rect 25004 37952 25010 37964
rect 25501 37961 25513 37964
rect 25547 37961 25559 37995
rect 26418 37992 26424 38004
rect 25501 37955 25559 37961
rect 26160 37964 26424 37992
rect 19978 37884 19984 37936
rect 20036 37924 20042 37936
rect 20809 37927 20867 37933
rect 20036 37896 20300 37924
rect 20036 37884 20042 37896
rect 19429 37859 19487 37865
rect 19429 37825 19441 37859
rect 19475 37825 19487 37859
rect 19429 37819 19487 37825
rect 19613 37859 19671 37865
rect 19613 37825 19625 37859
rect 19659 37856 19671 37859
rect 20162 37856 20168 37868
rect 19659 37828 20168 37856
rect 19659 37825 19671 37828
rect 19613 37819 19671 37825
rect 20162 37816 20168 37828
rect 20220 37816 20226 37868
rect 20272 37856 20300 37896
rect 20809 37893 20821 37927
rect 20855 37924 20867 37927
rect 21453 37927 21511 37933
rect 21453 37924 21465 37927
rect 20855 37896 21465 37924
rect 20855 37893 20867 37896
rect 20809 37887 20867 37893
rect 21453 37893 21465 37896
rect 21499 37924 21511 37927
rect 22278 37924 22284 37936
rect 21499 37896 22284 37924
rect 21499 37893 21511 37896
rect 21453 37887 21511 37893
rect 22278 37884 22284 37896
rect 22336 37884 22342 37936
rect 22664 37924 22692 37952
rect 26160 37933 26188 37964
rect 26418 37952 26424 37964
rect 26476 37952 26482 38004
rect 26605 37995 26663 38001
rect 26605 37961 26617 37995
rect 26651 37992 26663 37995
rect 27246 37992 27252 38004
rect 26651 37964 27252 37992
rect 26651 37961 26663 37964
rect 26605 37955 26663 37961
rect 27246 37952 27252 37964
rect 27304 37952 27310 38004
rect 28813 37995 28871 38001
rect 28813 37961 28825 37995
rect 28859 37961 28871 37995
rect 28813 37955 28871 37961
rect 26145 37927 26203 37933
rect 26145 37924 26157 37927
rect 22664 37896 22784 37924
rect 21269 37859 21327 37865
rect 21269 37856 21281 37859
rect 20272 37828 21281 37856
rect 21269 37825 21281 37828
rect 21315 37825 21327 37859
rect 21269 37819 21327 37825
rect 22002 37816 22008 37868
rect 22060 37816 22066 37868
rect 22189 37859 22247 37865
rect 22189 37825 22201 37859
rect 22235 37856 22247 37859
rect 22462 37856 22468 37868
rect 22235 37828 22468 37856
rect 22235 37825 22247 37828
rect 22189 37819 22247 37825
rect 22462 37816 22468 37828
rect 22520 37816 22526 37868
rect 22557 37859 22615 37865
rect 22557 37825 22569 37859
rect 22603 37856 22615 37859
rect 22646 37856 22652 37868
rect 22603 37828 22652 37856
rect 22603 37825 22615 37828
rect 22557 37819 22615 37825
rect 22646 37816 22652 37828
rect 22704 37816 22710 37868
rect 22756 37865 22784 37896
rect 24504 37896 26157 37924
rect 22741 37859 22799 37865
rect 22741 37825 22753 37859
rect 22787 37825 22799 37859
rect 22741 37819 22799 37825
rect 22830 37816 22836 37868
rect 22888 37816 22894 37868
rect 22922 37816 22928 37868
rect 22980 37816 22986 37868
rect 20898 37748 20904 37800
rect 20956 37748 20962 37800
rect 20990 37748 20996 37800
rect 21048 37748 21054 37800
rect 24504 37788 24532 37896
rect 26145 37893 26157 37896
rect 26191 37893 26203 37927
rect 26145 37887 26203 37893
rect 26237 37927 26295 37933
rect 26237 37893 26249 37927
rect 26283 37924 26295 37927
rect 28828 37924 28856 37955
rect 29270 37952 29276 38004
rect 29328 37952 29334 38004
rect 29641 37995 29699 38001
rect 29641 37961 29653 37995
rect 29687 37992 29699 37995
rect 29822 37992 29828 38004
rect 29687 37964 29828 37992
rect 29687 37961 29699 37964
rect 29641 37955 29699 37961
rect 29822 37952 29828 37964
rect 29880 37952 29886 38004
rect 31938 37992 31944 38004
rect 30024 37964 31944 37992
rect 26283 37896 27384 37924
rect 28828 37896 29868 37924
rect 26283 37893 26295 37896
rect 26237 37887 26295 37893
rect 27356 37868 27384 37896
rect 24765 37859 24823 37865
rect 24765 37825 24777 37859
rect 24811 37856 24823 37859
rect 24811 37828 24900 37856
rect 24811 37825 24823 37828
rect 24765 37819 24823 37825
rect 21473 37760 24532 37788
rect 24581 37791 24639 37797
rect 21473 37720 21501 37760
rect 24581 37757 24593 37791
rect 24627 37788 24639 37791
rect 24627 37760 24808 37788
rect 24627 37757 24639 37760
rect 24581 37751 24639 37757
rect 15672 37692 21501 37720
rect 14415 37689 14427 37692
rect 14369 37683 14427 37689
rect 21542 37680 21548 37732
rect 21600 37720 21606 37732
rect 21821 37723 21879 37729
rect 21821 37720 21833 37723
rect 21600 37692 21833 37720
rect 21600 37680 21606 37692
rect 21821 37689 21833 37692
rect 21867 37720 21879 37723
rect 22830 37720 22836 37732
rect 21867 37692 22836 37720
rect 21867 37689 21879 37692
rect 21821 37683 21879 37689
rect 22830 37680 22836 37692
rect 22888 37680 22894 37732
rect 24780 37664 24808 37760
rect 24872 37720 24900 37828
rect 24946 37816 24952 37868
rect 25004 37816 25010 37868
rect 25222 37816 25228 37868
rect 25280 37816 25286 37868
rect 25406 37816 25412 37868
rect 25464 37816 25470 37868
rect 25685 37859 25743 37865
rect 25685 37825 25697 37859
rect 25731 37856 25743 37859
rect 26789 37859 26847 37865
rect 25731 37828 25820 37856
rect 25731 37825 25743 37828
rect 25685 37819 25743 37825
rect 25041 37791 25099 37797
rect 25041 37757 25053 37791
rect 25087 37788 25099 37791
rect 25087 37760 25452 37788
rect 25087 37757 25099 37760
rect 25041 37751 25099 37757
rect 25222 37720 25228 37732
rect 24872 37692 25228 37720
rect 25222 37680 25228 37692
rect 25280 37680 25286 37732
rect 25424 37664 25452 37760
rect 25792 37729 25820 37828
rect 26789 37825 26801 37859
rect 26835 37856 26847 37859
rect 26835 37828 27108 37856
rect 26835 37825 26847 37828
rect 26789 37819 26847 37825
rect 26421 37791 26479 37797
rect 26421 37757 26433 37791
rect 26467 37788 26479 37791
rect 26970 37788 26976 37800
rect 26467 37760 26976 37788
rect 26467 37757 26479 37760
rect 26421 37751 26479 37757
rect 26970 37748 26976 37760
rect 27028 37748 27034 37800
rect 27080 37729 27108 37828
rect 27338 37816 27344 37868
rect 27396 37856 27402 37868
rect 27433 37859 27491 37865
rect 27433 37856 27445 37859
rect 27396 37828 27445 37856
rect 27396 37816 27402 37828
rect 27433 37825 27445 37828
rect 27479 37825 27491 37859
rect 27433 37819 27491 37825
rect 27982 37816 27988 37868
rect 28040 37816 28046 37868
rect 28077 37859 28135 37865
rect 28077 37825 28089 37859
rect 28123 37825 28135 37859
rect 28077 37819 28135 37825
rect 27522 37788 27528 37800
rect 27172 37760 27528 37788
rect 25777 37723 25835 37729
rect 25777 37689 25789 37723
rect 25823 37689 25835 37723
rect 25777 37683 25835 37689
rect 27065 37723 27123 37729
rect 27065 37689 27077 37723
rect 27111 37689 27123 37723
rect 27065 37683 27123 37689
rect 10134 37612 10140 37664
rect 10192 37612 10198 37664
rect 15194 37612 15200 37664
rect 15252 37652 15258 37664
rect 15565 37655 15623 37661
rect 15565 37652 15577 37655
rect 15252 37624 15577 37652
rect 15252 37612 15258 37624
rect 15565 37621 15577 37624
rect 15611 37621 15623 37655
rect 15565 37615 15623 37621
rect 19334 37612 19340 37664
rect 19392 37612 19398 37664
rect 19794 37612 19800 37664
rect 19852 37612 19858 37664
rect 21637 37655 21695 37661
rect 21637 37621 21649 37655
rect 21683 37652 21695 37655
rect 22094 37652 22100 37664
rect 21683 37624 22100 37652
rect 21683 37621 21695 37624
rect 21637 37615 21695 37621
rect 22094 37612 22100 37624
rect 22152 37612 22158 37664
rect 22370 37612 22376 37664
rect 22428 37612 22434 37664
rect 23106 37612 23112 37664
rect 23164 37612 23170 37664
rect 24762 37612 24768 37664
rect 24820 37612 24826 37664
rect 25406 37612 25412 37664
rect 25464 37612 25470 37664
rect 26234 37612 26240 37664
rect 26292 37652 26298 37664
rect 27172 37652 27200 37760
rect 27522 37748 27528 37760
rect 27580 37748 27586 37800
rect 27617 37791 27675 37797
rect 27617 37757 27629 37791
rect 27663 37757 27675 37791
rect 27617 37751 27675 37757
rect 27632 37720 27660 37751
rect 27798 37748 27804 37800
rect 27856 37788 27862 37800
rect 28092 37788 28120 37819
rect 29178 37816 29184 37868
rect 29236 37816 29242 37868
rect 29840 37865 29868 37896
rect 30024 37865 30052 37964
rect 31938 37952 31944 37964
rect 31996 37952 32002 38004
rect 30282 37884 30288 37936
rect 30340 37924 30346 37936
rect 30340 37896 30774 37924
rect 30340 37884 30346 37896
rect 29825 37859 29883 37865
rect 29825 37825 29837 37859
rect 29871 37825 29883 37859
rect 29825 37819 29883 37825
rect 30009 37859 30067 37865
rect 30009 37825 30021 37859
rect 30055 37825 30067 37859
rect 30009 37819 30067 37825
rect 32306 37816 32312 37868
rect 32364 37816 32370 37868
rect 29365 37791 29423 37797
rect 29365 37788 29377 37791
rect 27856 37760 28120 37788
rect 28184 37760 29377 37788
rect 27856 37748 27862 37760
rect 28184 37720 28212 37760
rect 29365 37757 29377 37760
rect 29411 37757 29423 37791
rect 29365 37751 29423 37757
rect 30285 37791 30343 37797
rect 30285 37757 30297 37791
rect 30331 37788 30343 37791
rect 30331 37760 32168 37788
rect 30331 37757 30343 37760
rect 30285 37751 30343 37757
rect 27540 37692 28212 37720
rect 28261 37723 28319 37729
rect 27540 37664 27568 37692
rect 28261 37689 28273 37723
rect 28307 37720 28319 37723
rect 32030 37720 32036 37732
rect 28307 37692 30144 37720
rect 28307 37689 28319 37692
rect 28261 37683 28319 37689
rect 26292 37624 27200 37652
rect 26292 37612 26298 37624
rect 27522 37612 27528 37664
rect 27580 37612 27586 37664
rect 30116 37652 30144 37692
rect 31312 37692 32036 37720
rect 31312 37652 31340 37692
rect 32030 37680 32036 37692
rect 32088 37680 32094 37732
rect 32140 37729 32168 37760
rect 32125 37723 32183 37729
rect 32125 37689 32137 37723
rect 32171 37689 32183 37723
rect 32125 37683 32183 37689
rect 30116 37624 31340 37652
rect 31754 37612 31760 37664
rect 31812 37612 31818 37664
rect 1104 37562 38272 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38272 37562
rect 1104 37488 38272 37510
rect 8662 37408 8668 37460
rect 8720 37448 8726 37460
rect 8941 37451 8999 37457
rect 8941 37448 8953 37451
rect 8720 37420 8953 37448
rect 8720 37408 8726 37420
rect 8941 37417 8953 37420
rect 8987 37417 8999 37451
rect 8941 37411 8999 37417
rect 16022 37408 16028 37460
rect 16080 37408 16086 37460
rect 17862 37408 17868 37460
rect 17920 37448 17926 37460
rect 19429 37451 19487 37457
rect 19429 37448 19441 37451
rect 17920 37420 19441 37448
rect 17920 37408 17926 37420
rect 19429 37417 19441 37420
rect 19475 37417 19487 37451
rect 19429 37411 19487 37417
rect 23106 37408 23112 37460
rect 23164 37448 23170 37460
rect 23569 37451 23627 37457
rect 23569 37448 23581 37451
rect 23164 37420 23581 37448
rect 23164 37408 23170 37420
rect 23569 37417 23581 37420
rect 23615 37417 23627 37451
rect 23569 37411 23627 37417
rect 24854 37408 24860 37460
rect 24912 37448 24918 37460
rect 25133 37451 25191 37457
rect 25133 37448 25145 37451
rect 24912 37420 25145 37448
rect 24912 37408 24918 37420
rect 25133 37417 25145 37420
rect 25179 37417 25191 37451
rect 25133 37411 25191 37417
rect 11146 37380 11152 37392
rect 10060 37352 11152 37380
rect 10060 37324 10088 37352
rect 11146 37340 11152 37352
rect 11204 37340 11210 37392
rect 13262 37340 13268 37392
rect 13320 37380 13326 37392
rect 15930 37380 15936 37392
rect 13320 37352 15936 37380
rect 13320 37340 13326 37352
rect 15930 37340 15936 37352
rect 15988 37340 15994 37392
rect 1765 37315 1823 37321
rect 1765 37281 1777 37315
rect 1811 37312 1823 37315
rect 6454 37312 6460 37324
rect 1811 37284 6460 37312
rect 1811 37281 1823 37284
rect 1765 37275 1823 37281
rect 6454 37272 6460 37284
rect 6512 37272 6518 37324
rect 10042 37272 10048 37324
rect 10100 37272 10106 37324
rect 10134 37272 10140 37324
rect 10192 37312 10198 37324
rect 16040 37312 16068 37408
rect 18230 37340 18236 37392
rect 18288 37380 18294 37392
rect 19058 37380 19064 37392
rect 18288 37352 19064 37380
rect 18288 37340 18294 37352
rect 19058 37340 19064 37352
rect 19116 37380 19122 37392
rect 25038 37380 25044 37392
rect 19116 37352 25044 37380
rect 19116 37340 19122 37352
rect 25038 37340 25044 37352
rect 25096 37340 25102 37392
rect 27062 37340 27068 37392
rect 27120 37380 27126 37392
rect 27120 37352 31340 37380
rect 27120 37340 27126 37352
rect 31312 37324 31340 37352
rect 18046 37312 18052 37324
rect 10192 37284 15976 37312
rect 16040 37284 18052 37312
rect 10192 37272 10198 37284
rect 9125 37247 9183 37253
rect 9125 37213 9137 37247
rect 9171 37244 9183 37247
rect 9861 37247 9919 37253
rect 9171 37216 9536 37244
rect 9171 37213 9183 37216
rect 9125 37207 9183 37213
rect 934 37136 940 37188
rect 992 37176 998 37188
rect 1489 37179 1547 37185
rect 1489 37176 1501 37179
rect 992 37148 1501 37176
rect 992 37136 998 37148
rect 1489 37145 1501 37148
rect 1535 37145 1547 37179
rect 1489 37139 1547 37145
rect 9508 37117 9536 37216
rect 9861 37213 9873 37247
rect 9907 37244 9919 37247
rect 10152 37244 10180 37272
rect 9907 37216 10180 37244
rect 9907 37213 9919 37216
rect 9861 37207 9919 37213
rect 14274 37204 14280 37256
rect 14332 37204 14338 37256
rect 15948 37244 15976 37284
rect 18046 37272 18052 37284
rect 18104 37272 18110 37324
rect 18156 37284 19288 37312
rect 18156 37244 18184 37284
rect 15948 37216 18184 37244
rect 19260 37244 19288 37284
rect 19334 37272 19340 37324
rect 19392 37312 19398 37324
rect 19521 37315 19579 37321
rect 19521 37312 19533 37315
rect 19392 37284 19533 37312
rect 19392 37272 19398 37284
rect 19521 37281 19533 37284
rect 19567 37281 19579 37315
rect 19521 37275 19579 37281
rect 19628 37284 21588 37312
rect 19628 37244 19656 37284
rect 21560 37256 21588 37284
rect 21836 37284 22232 37312
rect 21836 37256 21864 37284
rect 19260 37216 19656 37244
rect 19705 37247 19763 37253
rect 19705 37213 19717 37247
rect 19751 37244 19763 37247
rect 19794 37244 19800 37256
rect 19751 37216 19800 37244
rect 19751 37213 19763 37216
rect 19705 37207 19763 37213
rect 19794 37204 19800 37216
rect 19852 37204 19858 37256
rect 21542 37204 21548 37256
rect 21600 37204 21606 37256
rect 21818 37204 21824 37256
rect 21876 37204 21882 37256
rect 21910 37204 21916 37256
rect 21968 37204 21974 37256
rect 22094 37204 22100 37256
rect 22152 37204 22158 37256
rect 22204 37253 22232 37284
rect 24670 37272 24676 37324
rect 24728 37312 24734 37324
rect 24765 37315 24823 37321
rect 24765 37312 24777 37315
rect 24728 37284 24777 37312
rect 24728 37272 24734 37284
rect 24765 37281 24777 37284
rect 24811 37281 24823 37315
rect 24765 37275 24823 37281
rect 26970 37272 26976 37324
rect 27028 37272 27034 37324
rect 27798 37312 27804 37324
rect 27172 37284 27804 37312
rect 22189 37247 22247 37253
rect 22189 37213 22201 37247
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22281 37247 22339 37253
rect 22281 37213 22293 37247
rect 22327 37213 22339 37247
rect 22281 37207 22339 37213
rect 15102 37136 15108 37188
rect 15160 37136 15166 37188
rect 19426 37136 19432 37188
rect 19484 37136 19490 37188
rect 22296 37176 22324 37207
rect 22370 37204 22376 37256
rect 22428 37244 22434 37256
rect 22557 37247 22615 37253
rect 22557 37244 22569 37247
rect 22428 37216 22569 37244
rect 22428 37204 22434 37216
rect 22557 37213 22569 37216
rect 22603 37213 22615 37247
rect 22557 37207 22615 37213
rect 22646 37204 22652 37256
rect 22704 37244 22710 37256
rect 23106 37253 23112 37256
rect 23063 37247 23112 37253
rect 22704 37216 22749 37244
rect 22704 37204 22710 37216
rect 23063 37213 23075 37247
rect 23109 37213 23112 37247
rect 23063 37207 23112 37213
rect 23106 37204 23112 37207
rect 23164 37204 23170 37256
rect 23753 37247 23811 37253
rect 23753 37244 23765 37247
rect 23216 37216 23765 37244
rect 19812 37148 22324 37176
rect 9493 37111 9551 37117
rect 9493 37077 9505 37111
rect 9539 37077 9551 37111
rect 9493 37071 9551 37077
rect 9953 37111 10011 37117
rect 9953 37077 9965 37111
rect 9999 37108 10011 37111
rect 11790 37108 11796 37120
rect 9999 37080 11796 37108
rect 9999 37077 10011 37080
rect 9953 37071 10011 37077
rect 11790 37068 11796 37080
rect 11848 37068 11854 37120
rect 15930 37068 15936 37120
rect 15988 37108 15994 37120
rect 18782 37108 18788 37120
rect 15988 37080 18788 37108
rect 15988 37068 15994 37080
rect 18782 37068 18788 37080
rect 18840 37068 18846 37120
rect 19150 37068 19156 37120
rect 19208 37108 19214 37120
rect 19812 37108 19840 37148
rect 22830 37136 22836 37188
rect 22888 37136 22894 37188
rect 22922 37136 22928 37188
rect 22980 37136 22986 37188
rect 23216 37176 23244 37216
rect 23753 37213 23765 37216
rect 23799 37213 23811 37247
rect 23753 37207 23811 37213
rect 23842 37204 23848 37256
rect 23900 37204 23906 37256
rect 24949 37247 25007 37253
rect 24949 37213 24961 37247
rect 24995 37244 25007 37247
rect 25222 37244 25228 37256
rect 24995 37216 25228 37244
rect 24995 37213 25007 37216
rect 24949 37207 25007 37213
rect 25222 37204 25228 37216
rect 25280 37244 25286 37256
rect 27172 37253 27200 37284
rect 27798 37272 27804 37284
rect 27856 37272 27862 37324
rect 29178 37272 29184 37324
rect 29236 37312 29242 37324
rect 31202 37312 31208 37324
rect 29236 37284 31208 37312
rect 29236 37272 29242 37284
rect 31202 37272 31208 37284
rect 31260 37272 31266 37324
rect 31294 37272 31300 37324
rect 31352 37272 31358 37324
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 25280 37216 27169 37244
rect 25280 37204 25286 37216
rect 23124 37148 23244 37176
rect 19208 37080 19840 37108
rect 19889 37111 19947 37117
rect 19208 37068 19214 37080
rect 19889 37077 19901 37111
rect 19935 37108 19947 37111
rect 20070 37108 20076 37120
rect 19935 37080 20076 37108
rect 19935 37077 19947 37080
rect 19889 37071 19947 37077
rect 20070 37068 20076 37080
rect 20128 37068 20134 37120
rect 22465 37111 22523 37117
rect 22465 37077 22477 37111
rect 22511 37108 22523 37111
rect 23124 37108 23152 37148
rect 23566 37136 23572 37188
rect 23624 37136 23630 37188
rect 25884 37120 25912 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 27341 37247 27399 37253
rect 27341 37213 27353 37247
rect 27387 37244 27399 37247
rect 34514 37244 34520 37256
rect 27387 37216 34520 37244
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 34514 37204 34520 37216
rect 34572 37204 34578 37256
rect 37645 37247 37703 37253
rect 37645 37213 37657 37247
rect 37691 37213 37703 37247
rect 37645 37207 37703 37213
rect 32306 37176 32312 37188
rect 30760 37148 32312 37176
rect 22511 37080 23152 37108
rect 22511 37077 22523 37080
rect 22465 37071 22523 37077
rect 23198 37068 23204 37120
rect 23256 37068 23262 37120
rect 23658 37068 23664 37120
rect 23716 37108 23722 37120
rect 24029 37111 24087 37117
rect 24029 37108 24041 37111
rect 23716 37080 24041 37108
rect 23716 37068 23722 37080
rect 24029 37077 24041 37080
rect 24075 37077 24087 37111
rect 24029 37071 24087 37077
rect 25866 37068 25872 37120
rect 25924 37068 25930 37120
rect 30760 37117 30788 37148
rect 32306 37136 32312 37148
rect 32364 37136 32370 37188
rect 37274 37136 37280 37188
rect 37332 37176 37338 37188
rect 37660 37176 37688 37207
rect 37332 37148 37688 37176
rect 37332 37136 37338 37148
rect 30745 37111 30803 37117
rect 30745 37077 30757 37111
rect 30791 37077 30803 37111
rect 30745 37071 30803 37077
rect 31110 37068 31116 37120
rect 31168 37068 31174 37120
rect 31202 37068 31208 37120
rect 31260 37108 31266 37120
rect 33134 37108 33140 37120
rect 31260 37080 33140 37108
rect 31260 37068 31266 37080
rect 33134 37068 33140 37080
rect 33192 37068 33198 37120
rect 37826 37068 37832 37120
rect 37884 37068 37890 37120
rect 1104 37018 38272 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38272 37018
rect 1104 36944 38272 36966
rect 18230 36904 18236 36916
rect 15948 36876 18236 36904
rect 15948 36845 15976 36876
rect 18230 36864 18236 36876
rect 18288 36864 18294 36916
rect 22646 36864 22652 36916
rect 22704 36864 22710 36916
rect 23109 36907 23167 36913
rect 23109 36873 23121 36907
rect 23155 36904 23167 36907
rect 23842 36904 23848 36916
rect 23155 36876 23848 36904
rect 23155 36873 23167 36876
rect 23109 36867 23167 36873
rect 23842 36864 23848 36876
rect 23900 36864 23906 36916
rect 24394 36864 24400 36916
rect 24452 36904 24458 36916
rect 28258 36904 28264 36916
rect 24452 36876 28264 36904
rect 24452 36864 24458 36876
rect 28258 36864 28264 36876
rect 28316 36864 28322 36916
rect 31754 36904 31760 36916
rect 31726 36864 31760 36904
rect 31812 36864 31818 36916
rect 15933 36839 15991 36845
rect 15933 36805 15945 36839
rect 15979 36805 15991 36839
rect 15933 36799 15991 36805
rect 18874 36796 18880 36848
rect 18932 36836 18938 36848
rect 21450 36836 21456 36848
rect 18932 36808 21456 36836
rect 18932 36796 18938 36808
rect 21450 36796 21456 36808
rect 21508 36836 21514 36848
rect 21910 36836 21916 36848
rect 21508 36808 21916 36836
rect 21508 36796 21514 36808
rect 21910 36796 21916 36808
rect 21968 36796 21974 36848
rect 22664 36836 22692 36864
rect 22664 36808 23336 36836
rect 7009 36771 7067 36777
rect 7009 36737 7021 36771
rect 7055 36737 7067 36771
rect 7009 36731 7067 36737
rect 7024 36700 7052 36731
rect 15838 36728 15844 36780
rect 15896 36768 15902 36780
rect 16117 36771 16175 36777
rect 16117 36768 16129 36771
rect 15896 36740 16129 36768
rect 15896 36728 15902 36740
rect 16117 36737 16129 36740
rect 16163 36737 16175 36771
rect 16117 36731 16175 36737
rect 16206 36728 16212 36780
rect 16264 36728 16270 36780
rect 16298 36728 16304 36780
rect 16356 36777 16362 36780
rect 16356 36768 16364 36777
rect 16356 36740 16401 36768
rect 16356 36731 16364 36740
rect 16356 36728 16362 36731
rect 20162 36728 20168 36780
rect 20220 36768 20226 36780
rect 22925 36771 22983 36777
rect 22925 36768 22937 36771
rect 20220 36740 22937 36768
rect 20220 36728 20226 36740
rect 22925 36737 22937 36740
rect 22971 36737 22983 36771
rect 23308 36768 23336 36808
rect 24946 36796 24952 36848
rect 25004 36836 25010 36848
rect 25501 36839 25559 36845
rect 25501 36836 25513 36839
rect 25004 36808 25513 36836
rect 25004 36796 25010 36808
rect 25501 36805 25513 36808
rect 25547 36836 25559 36839
rect 29730 36836 29736 36848
rect 25547 36808 26188 36836
rect 25547 36805 25559 36808
rect 25501 36799 25559 36805
rect 26160 36780 26188 36808
rect 27540 36808 29736 36836
rect 25225 36771 25283 36777
rect 25225 36768 25237 36771
rect 23308 36740 25237 36768
rect 22925 36731 22983 36737
rect 25225 36737 25237 36740
rect 25271 36737 25283 36771
rect 25225 36731 25283 36737
rect 7098 36700 7104 36712
rect 7024 36672 7104 36700
rect 7098 36660 7104 36672
rect 7156 36660 7162 36712
rect 17218 36660 17224 36712
rect 17276 36700 17282 36712
rect 20438 36700 20444 36712
rect 17276 36672 20444 36700
rect 17276 36660 17282 36672
rect 20438 36660 20444 36672
rect 20496 36660 20502 36712
rect 22741 36703 22799 36709
rect 22741 36669 22753 36703
rect 22787 36700 22799 36703
rect 25240 36700 25268 36731
rect 25314 36728 25320 36780
rect 25372 36768 25378 36780
rect 25409 36771 25467 36777
rect 25409 36768 25421 36771
rect 25372 36740 25421 36768
rect 25372 36728 25378 36740
rect 25409 36737 25421 36740
rect 25455 36737 25467 36771
rect 25409 36731 25467 36737
rect 25593 36771 25651 36777
rect 25593 36737 25605 36771
rect 25639 36768 25651 36771
rect 25958 36768 25964 36780
rect 25639 36740 25964 36768
rect 25639 36737 25651 36740
rect 25593 36731 25651 36737
rect 25958 36728 25964 36740
rect 26016 36728 26022 36780
rect 26142 36728 26148 36780
rect 26200 36728 26206 36780
rect 27540 36700 27568 36808
rect 29730 36796 29736 36808
rect 29788 36836 29794 36848
rect 31110 36836 31116 36848
rect 29788 36808 31116 36836
rect 29788 36796 29794 36808
rect 31110 36796 31116 36808
rect 31168 36836 31174 36848
rect 31726 36836 31754 36864
rect 31168 36808 31754 36836
rect 31168 36796 31174 36808
rect 27617 36771 27675 36777
rect 27617 36737 27629 36771
rect 27663 36768 27675 36771
rect 27663 36740 28764 36768
rect 27663 36737 27675 36740
rect 27617 36731 27675 36737
rect 28736 36712 28764 36740
rect 32950 36728 32956 36780
rect 33008 36728 33014 36780
rect 22787 36672 22968 36700
rect 25240 36672 27568 36700
rect 22787 36669 22799 36672
rect 22741 36663 22799 36669
rect 22940 36644 22968 36672
rect 28718 36660 28724 36712
rect 28776 36660 28782 36712
rect 11790 36592 11796 36644
rect 11848 36632 11854 36644
rect 11848 36604 20944 36632
rect 11848 36592 11854 36604
rect 20916 36576 20944 36604
rect 22922 36592 22928 36644
rect 22980 36592 22986 36644
rect 24578 36592 24584 36644
rect 24636 36632 24642 36644
rect 26786 36632 26792 36644
rect 24636 36604 26792 36632
rect 24636 36592 24642 36604
rect 26786 36592 26792 36604
rect 26844 36632 26850 36644
rect 30006 36632 30012 36644
rect 26844 36604 30012 36632
rect 26844 36592 26850 36604
rect 30006 36592 30012 36604
rect 30064 36592 30070 36644
rect 7006 36524 7012 36576
rect 7064 36564 7070 36576
rect 7101 36567 7159 36573
rect 7101 36564 7113 36567
rect 7064 36536 7113 36564
rect 7064 36524 7070 36536
rect 7101 36533 7113 36536
rect 7147 36533 7159 36567
rect 7101 36527 7159 36533
rect 15286 36524 15292 36576
rect 15344 36564 15350 36576
rect 15933 36567 15991 36573
rect 15933 36564 15945 36567
rect 15344 36536 15945 36564
rect 15344 36524 15350 36536
rect 15933 36533 15945 36536
rect 15979 36533 15991 36567
rect 15933 36527 15991 36533
rect 16206 36524 16212 36576
rect 16264 36564 16270 36576
rect 18506 36564 18512 36576
rect 16264 36536 18512 36564
rect 16264 36524 16270 36536
rect 18506 36524 18512 36536
rect 18564 36524 18570 36576
rect 19886 36524 19892 36576
rect 19944 36564 19950 36576
rect 20346 36564 20352 36576
rect 19944 36536 20352 36564
rect 19944 36524 19950 36536
rect 20346 36524 20352 36536
rect 20404 36524 20410 36576
rect 20898 36524 20904 36576
rect 20956 36524 20962 36576
rect 21910 36524 21916 36576
rect 21968 36564 21974 36576
rect 25682 36564 25688 36576
rect 21968 36536 25688 36564
rect 21968 36524 21974 36536
rect 25682 36524 25688 36536
rect 25740 36524 25746 36576
rect 25774 36524 25780 36576
rect 25832 36524 25838 36576
rect 27430 36524 27436 36576
rect 27488 36564 27494 36576
rect 27709 36567 27767 36573
rect 27709 36564 27721 36567
rect 27488 36536 27721 36564
rect 27488 36524 27494 36536
rect 27709 36533 27721 36536
rect 27755 36533 27767 36567
rect 27709 36527 27767 36533
rect 32766 36524 32772 36576
rect 32824 36524 32830 36576
rect 1104 36474 38272 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38272 36474
rect 1104 36400 38272 36422
rect 7006 36320 7012 36372
rect 7064 36320 7070 36372
rect 17494 36320 17500 36372
rect 17552 36360 17558 36372
rect 18322 36360 18328 36372
rect 17552 36332 18328 36360
rect 17552 36320 17558 36332
rect 18322 36320 18328 36332
rect 18380 36320 18386 36372
rect 18414 36320 18420 36372
rect 18472 36360 18478 36372
rect 19061 36363 19119 36369
rect 19061 36360 19073 36363
rect 18472 36332 19073 36360
rect 18472 36320 18478 36332
rect 19061 36329 19073 36332
rect 19107 36329 19119 36363
rect 19061 36323 19119 36329
rect 19426 36320 19432 36372
rect 19484 36360 19490 36372
rect 20901 36363 20959 36369
rect 20901 36360 20913 36363
rect 19484 36332 20913 36360
rect 19484 36320 19490 36332
rect 20901 36329 20913 36332
rect 20947 36329 20959 36363
rect 20901 36323 20959 36329
rect 22462 36320 22468 36372
rect 22520 36360 22526 36372
rect 23290 36360 23296 36372
rect 22520 36332 23296 36360
rect 22520 36320 22526 36332
rect 23290 36320 23296 36332
rect 23348 36320 23354 36372
rect 23477 36363 23535 36369
rect 23477 36329 23489 36363
rect 23523 36360 23535 36363
rect 23566 36360 23572 36372
rect 23523 36332 23572 36360
rect 23523 36329 23535 36332
rect 23477 36323 23535 36329
rect 23566 36320 23572 36332
rect 23624 36320 23630 36372
rect 25038 36320 25044 36372
rect 25096 36360 25102 36372
rect 26234 36360 26240 36372
rect 25096 36332 26240 36360
rect 25096 36320 25102 36332
rect 26234 36320 26240 36332
rect 26292 36320 26298 36372
rect 26418 36320 26424 36372
rect 26476 36320 26482 36372
rect 26786 36320 26792 36372
rect 26844 36320 26850 36372
rect 29086 36360 29092 36372
rect 26896 36332 29092 36360
rect 6917 36227 6975 36233
rect 6917 36193 6929 36227
rect 6963 36224 6975 36227
rect 7024 36224 7052 36320
rect 12805 36295 12863 36301
rect 12805 36261 12817 36295
rect 12851 36292 12863 36295
rect 13541 36295 13599 36301
rect 13541 36292 13553 36295
rect 12851 36264 13553 36292
rect 12851 36261 12863 36264
rect 12805 36255 12863 36261
rect 13541 36261 13553 36264
rect 13587 36261 13599 36295
rect 17770 36292 17776 36304
rect 13541 36255 13599 36261
rect 13648 36264 17776 36292
rect 6963 36196 7052 36224
rect 6963 36193 6975 36196
rect 6917 36187 6975 36193
rect 10686 36184 10692 36236
rect 10744 36224 10750 36236
rect 13648 36224 13676 36264
rect 17126 36224 17132 36236
rect 10744 36196 13676 36224
rect 15120 36196 17132 36224
rect 10744 36184 10750 36196
rect 4709 36159 4767 36165
rect 4709 36125 4721 36159
rect 4755 36125 4767 36159
rect 4709 36119 4767 36125
rect 4801 36159 4859 36165
rect 4801 36125 4813 36159
rect 4847 36156 4859 36159
rect 4985 36159 5043 36165
rect 4985 36156 4997 36159
rect 4847 36128 4997 36156
rect 4847 36125 4859 36128
rect 4801 36119 4859 36125
rect 4985 36125 4997 36128
rect 5031 36125 5043 36159
rect 4985 36119 5043 36125
rect 4724 36020 4752 36119
rect 8938 36116 8944 36168
rect 8996 36116 9002 36168
rect 10594 36156 10600 36168
rect 10350 36142 10600 36156
rect 10336 36128 10600 36142
rect 5261 36091 5319 36097
rect 5261 36057 5273 36091
rect 5307 36088 5319 36091
rect 5534 36088 5540 36100
rect 5307 36060 5540 36088
rect 5307 36057 5319 36060
rect 5261 36051 5319 36057
rect 5534 36048 5540 36060
rect 5592 36048 5598 36100
rect 6822 36088 6828 36100
rect 6486 36060 6828 36088
rect 6822 36048 6828 36060
rect 6880 36048 6886 36100
rect 7190 36048 7196 36100
rect 7248 36048 7254 36100
rect 8478 36088 8484 36100
rect 8418 36060 8484 36088
rect 8478 36048 8484 36060
rect 8536 36088 8542 36100
rect 8536 36060 8800 36088
rect 8536 36048 8542 36060
rect 5350 36020 5356 36032
rect 4724 35992 5356 36020
rect 5350 35980 5356 35992
rect 5408 35980 5414 36032
rect 6730 35980 6736 36032
rect 6788 35980 6794 36032
rect 8662 35980 8668 36032
rect 8720 35980 8726 36032
rect 8772 36020 8800 36060
rect 9214 36048 9220 36100
rect 9272 36048 9278 36100
rect 10336 36020 10364 36128
rect 10594 36116 10600 36128
rect 10652 36116 10658 36168
rect 12253 36159 12311 36165
rect 12253 36125 12265 36159
rect 12299 36156 12311 36159
rect 12342 36156 12348 36168
rect 12299 36128 12348 36156
rect 12299 36125 12311 36128
rect 12253 36119 12311 36125
rect 12342 36116 12348 36128
rect 12400 36116 12406 36168
rect 12544 36165 12572 36196
rect 12529 36159 12587 36165
rect 12529 36125 12541 36159
rect 12575 36125 12587 36159
rect 12529 36119 12587 36125
rect 12618 36116 12624 36168
rect 12676 36116 12682 36168
rect 12802 36116 12808 36168
rect 12860 36156 12866 36168
rect 13111 36159 13169 36165
rect 13111 36156 13123 36159
rect 12860 36128 13123 36156
rect 12860 36116 12866 36128
rect 13111 36125 13123 36128
rect 13157 36125 13169 36159
rect 13111 36119 13169 36125
rect 13630 36116 13636 36168
rect 13688 36116 13694 36168
rect 15120 36165 15148 36196
rect 17126 36184 17132 36196
rect 17184 36184 17190 36236
rect 15105 36159 15163 36165
rect 15105 36125 15117 36159
rect 15151 36125 15163 36159
rect 15105 36119 15163 36125
rect 15194 36116 15200 36168
rect 15252 36116 15258 36168
rect 15286 36116 15292 36168
rect 15344 36116 15350 36168
rect 15562 36116 15568 36168
rect 15620 36116 15626 36168
rect 17420 36165 17448 36264
rect 17770 36252 17776 36264
rect 17828 36252 17834 36304
rect 18598 36252 18604 36304
rect 18656 36292 18662 36304
rect 18656 36264 19656 36292
rect 18656 36252 18662 36264
rect 18322 36184 18328 36236
rect 18380 36184 18386 36236
rect 18690 36184 18696 36236
rect 18748 36224 18754 36236
rect 18748 36196 19472 36224
rect 18748 36184 18754 36196
rect 17405 36159 17463 36165
rect 17405 36125 17417 36159
rect 17451 36125 17463 36159
rect 17405 36119 17463 36125
rect 17678 36116 17684 36168
rect 17736 36116 17742 36168
rect 17770 36116 17776 36168
rect 17828 36116 17834 36168
rect 18049 36159 18107 36165
rect 18049 36125 18061 36159
rect 18095 36156 18107 36159
rect 18138 36156 18144 36168
rect 18095 36128 18144 36156
rect 18095 36125 18107 36128
rect 18049 36119 18107 36125
rect 18138 36116 18144 36128
rect 18196 36116 18202 36168
rect 18233 36159 18291 36165
rect 18233 36125 18245 36159
rect 18279 36156 18291 36159
rect 18340 36156 18368 36184
rect 18279 36128 18368 36156
rect 18417 36159 18475 36165
rect 18279 36125 18291 36128
rect 18233 36119 18291 36125
rect 18417 36125 18429 36159
rect 18463 36125 18475 36159
rect 18417 36119 18475 36125
rect 12434 36048 12440 36100
rect 12492 36048 12498 36100
rect 14734 36048 14740 36100
rect 14792 36088 14798 36100
rect 15407 36091 15465 36097
rect 15407 36088 15419 36091
rect 14792 36060 15419 36088
rect 14792 36048 14798 36060
rect 15407 36057 15419 36060
rect 15453 36057 15465 36091
rect 15407 36051 15465 36057
rect 17589 36091 17647 36097
rect 17589 36057 17601 36091
rect 17635 36057 17647 36091
rect 18432 36088 18460 36119
rect 18506 36116 18512 36168
rect 18564 36116 18570 36168
rect 18782 36116 18788 36168
rect 18840 36116 18846 36168
rect 18874 36116 18880 36168
rect 18932 36165 18938 36168
rect 18932 36156 18940 36165
rect 18932 36128 18977 36156
rect 18932 36119 18940 36128
rect 18932 36116 18938 36119
rect 17589 36051 17647 36057
rect 17972 36060 18460 36088
rect 8772 35992 10364 36020
rect 12986 35980 12992 36032
rect 13044 35980 13050 36032
rect 13173 36023 13231 36029
rect 13173 35989 13185 36023
rect 13219 36020 13231 36023
rect 14921 36023 14979 36029
rect 14921 36020 14933 36023
rect 13219 35992 14933 36020
rect 13219 35989 13231 35992
rect 13173 35983 13231 35989
rect 14921 35989 14933 35992
rect 14967 35989 14979 36023
rect 14921 35983 14979 35989
rect 17402 35980 17408 36032
rect 17460 36020 17466 36032
rect 17604 36020 17632 36051
rect 17972 36029 18000 36060
rect 18598 36048 18604 36100
rect 18656 36088 18662 36100
rect 18693 36091 18751 36097
rect 18693 36088 18705 36091
rect 18656 36060 18705 36088
rect 18656 36048 18662 36060
rect 18693 36057 18705 36060
rect 18739 36057 18751 36091
rect 19334 36088 19340 36100
rect 18693 36051 18751 36057
rect 18984 36060 19340 36088
rect 17460 35992 17632 36020
rect 17957 36023 18015 36029
rect 17460 35980 17466 35992
rect 17957 35989 17969 36023
rect 18003 35989 18015 36023
rect 17957 35983 18015 35989
rect 18233 36023 18291 36029
rect 18233 35989 18245 36023
rect 18279 36020 18291 36023
rect 18984 36020 19012 36060
rect 19334 36048 19340 36060
rect 19392 36048 19398 36100
rect 18279 35992 19012 36020
rect 19444 36020 19472 36196
rect 19628 36088 19656 36264
rect 19720 36264 22508 36292
rect 19720 36165 19748 36264
rect 22094 36224 22100 36236
rect 19812 36196 22100 36224
rect 19812 36165 19840 36196
rect 19705 36159 19763 36165
rect 19705 36125 19717 36159
rect 19751 36125 19763 36159
rect 19705 36119 19763 36125
rect 19797 36159 19855 36165
rect 19797 36125 19809 36159
rect 19843 36125 19855 36159
rect 19797 36119 19855 36125
rect 19886 36116 19892 36168
rect 19944 36156 19950 36168
rect 20073 36159 20131 36165
rect 20073 36156 20085 36159
rect 19944 36128 20085 36156
rect 19944 36116 19950 36128
rect 20073 36125 20085 36128
rect 20119 36125 20131 36159
rect 20073 36119 20131 36125
rect 20165 36159 20223 36165
rect 20165 36125 20177 36159
rect 20211 36156 20223 36159
rect 20211 36128 20300 36156
rect 20211 36125 20223 36128
rect 20165 36119 20223 36125
rect 19904 36088 19932 36116
rect 19628 36060 19932 36088
rect 19981 36091 20039 36097
rect 19981 36057 19993 36091
rect 20027 36057 20039 36091
rect 20272 36088 20300 36128
rect 20346 36116 20352 36168
rect 20404 36116 20410 36168
rect 20438 36116 20444 36168
rect 20496 36156 20502 36168
rect 20640 36165 20668 36196
rect 22094 36184 22100 36196
rect 22152 36184 22158 36236
rect 22480 36168 22508 36264
rect 22572 36264 23336 36292
rect 20625 36159 20683 36165
rect 20496 36128 20576 36156
rect 20496 36116 20502 36128
rect 20548 36097 20576 36128
rect 20625 36125 20637 36159
rect 20671 36125 20683 36159
rect 20625 36119 20683 36125
rect 20714 36116 20720 36168
rect 20772 36156 20778 36168
rect 20772 36128 22012 36156
rect 20772 36116 20778 36128
rect 20533 36091 20591 36097
rect 20272 36060 20484 36088
rect 19981 36051 20039 36057
rect 19705 36023 19763 36029
rect 19705 36020 19717 36023
rect 19444 35992 19717 36020
rect 18279 35989 18291 35992
rect 18233 35983 18291 35989
rect 19705 35989 19717 35992
rect 19751 35989 19763 36023
rect 19996 36020 20024 36051
rect 20346 36020 20352 36032
rect 19996 35992 20352 36020
rect 19705 35983 19763 35989
rect 20346 35980 20352 35992
rect 20404 35980 20410 36032
rect 20456 36020 20484 36060
rect 20533 36057 20545 36091
rect 20579 36088 20591 36091
rect 21984 36088 22012 36128
rect 22462 36116 22468 36168
rect 22520 36116 22526 36168
rect 22572 36088 22600 36264
rect 22646 36184 22652 36236
rect 22704 36224 22710 36236
rect 22704 36196 23244 36224
rect 22704 36184 22710 36196
rect 22738 36116 22744 36168
rect 22796 36156 22802 36168
rect 23216 36165 23244 36196
rect 23308 36165 23336 36264
rect 25056 36224 25084 36320
rect 26050 36252 26056 36304
rect 26108 36292 26114 36304
rect 26145 36295 26203 36301
rect 26145 36292 26157 36295
rect 26108 36264 26157 36292
rect 26108 36252 26114 36264
rect 26145 36261 26157 36264
rect 26191 36261 26203 36295
rect 26145 36255 26203 36261
rect 25056 36196 25268 36224
rect 22925 36159 22983 36165
rect 22796 36152 22876 36156
rect 22925 36152 22937 36159
rect 22796 36128 22937 36152
rect 22796 36116 22802 36128
rect 22848 36125 22937 36128
rect 22971 36125 22983 36159
rect 22848 36124 22983 36125
rect 22925 36119 22983 36124
rect 23109 36159 23167 36165
rect 23109 36125 23121 36159
rect 23155 36125 23167 36159
rect 23109 36119 23167 36125
rect 23201 36159 23259 36165
rect 23201 36125 23213 36159
rect 23247 36125 23259 36159
rect 23201 36119 23259 36125
rect 23293 36159 23351 36165
rect 23293 36125 23305 36159
rect 23339 36156 23351 36159
rect 24118 36156 24124 36168
rect 23339 36128 24124 36156
rect 23339 36125 23351 36128
rect 23293 36119 23351 36125
rect 20579 36060 21772 36088
rect 21984 36060 22600 36088
rect 20579 36057 20591 36060
rect 20533 36051 20591 36057
rect 21634 36020 21640 36032
rect 20456 35992 21640 36020
rect 21634 35980 21640 35992
rect 21692 35980 21698 36032
rect 21744 36020 21772 36060
rect 23124 36020 23152 36119
rect 23216 36088 23244 36119
rect 24118 36116 24124 36128
rect 24176 36116 24182 36168
rect 24946 36116 24952 36168
rect 25004 36116 25010 36168
rect 25240 36165 25268 36196
rect 25314 36184 25320 36236
rect 25372 36224 25378 36236
rect 26436 36224 26464 36320
rect 25372 36196 25437 36224
rect 25372 36184 25378 36196
rect 25409 36165 25437 36196
rect 25884 36196 26740 36224
rect 25133 36159 25191 36165
rect 25133 36125 25145 36159
rect 25179 36125 25191 36159
rect 25133 36119 25191 36125
rect 25225 36159 25283 36165
rect 25225 36125 25237 36159
rect 25271 36125 25283 36159
rect 25225 36119 25283 36125
rect 25409 36159 25467 36165
rect 25409 36125 25421 36159
rect 25455 36125 25467 36159
rect 25409 36119 25467 36125
rect 24964 36088 24992 36116
rect 23216 36060 24992 36088
rect 25148 36088 25176 36119
rect 25498 36116 25504 36168
rect 25556 36116 25562 36168
rect 25593 36159 25651 36165
rect 25593 36125 25605 36159
rect 25639 36158 25651 36159
rect 25639 36156 25820 36158
rect 25884 36156 25912 36196
rect 25639 36130 25912 36156
rect 25639 36125 25651 36130
rect 25792 36128 25912 36130
rect 25593 36119 25651 36125
rect 25958 36116 25964 36168
rect 26016 36116 26022 36168
rect 26326 36116 26332 36168
rect 26384 36116 26390 36168
rect 26418 36116 26424 36168
rect 26476 36156 26482 36168
rect 26712 36165 26740 36196
rect 26804 36165 26832 36320
rect 26697 36159 26755 36165
rect 26476 36128 26521 36156
rect 26476 36116 26482 36128
rect 26697 36125 26709 36159
rect 26743 36125 26755 36159
rect 26697 36119 26755 36125
rect 26794 36159 26852 36165
rect 26794 36125 26806 36159
rect 26840 36125 26852 36159
rect 26794 36119 26852 36125
rect 25314 36088 25320 36100
rect 25148 36060 25320 36088
rect 25314 36048 25320 36060
rect 25372 36048 25378 36100
rect 25777 36091 25835 36097
rect 25777 36057 25789 36091
rect 25823 36057 25835 36091
rect 25777 36051 25835 36057
rect 25869 36091 25927 36097
rect 25869 36057 25881 36091
rect 25915 36088 25927 36091
rect 26050 36088 26056 36100
rect 25915 36060 26056 36088
rect 25915 36057 25927 36060
rect 25869 36051 25927 36057
rect 21744 35992 23152 36020
rect 24949 36023 25007 36029
rect 24949 35989 24961 36023
rect 24995 36020 25007 36023
rect 25130 36020 25136 36032
rect 24995 35992 25136 36020
rect 24995 35989 25007 35992
rect 24949 35983 25007 35989
rect 25130 35980 25136 35992
rect 25188 35980 25194 36032
rect 25590 35980 25596 36032
rect 25648 36020 25654 36032
rect 25792 36020 25820 36051
rect 26050 36048 26056 36060
rect 26108 36088 26114 36100
rect 26234 36088 26240 36100
rect 26108 36060 26240 36088
rect 26108 36048 26114 36060
rect 26234 36048 26240 36060
rect 26292 36048 26298 36100
rect 25648 35992 25820 36020
rect 26344 36020 26372 36116
rect 26510 36048 26516 36100
rect 26568 36088 26574 36100
rect 26605 36091 26663 36097
rect 26605 36088 26617 36091
rect 26568 36060 26617 36088
rect 26568 36048 26574 36060
rect 26605 36057 26617 36060
rect 26651 36057 26663 36091
rect 26605 36051 26663 36057
rect 26896 36020 26924 36332
rect 29086 36320 29092 36332
rect 29144 36360 29150 36372
rect 29362 36360 29368 36372
rect 29144 36332 29368 36360
rect 29144 36320 29150 36332
rect 29362 36320 29368 36332
rect 29420 36320 29426 36372
rect 27430 36252 27436 36304
rect 27488 36252 27494 36304
rect 29273 36295 29331 36301
rect 29273 36292 29285 36295
rect 28966 36264 29285 36292
rect 27448 36224 27476 36252
rect 27525 36227 27583 36233
rect 27525 36224 27537 36227
rect 27448 36196 27537 36224
rect 27525 36193 27537 36196
rect 27571 36193 27583 36227
rect 27525 36187 27583 36193
rect 27798 36184 27804 36236
rect 27856 36224 27862 36236
rect 28966 36224 28994 36264
rect 29273 36261 29285 36264
rect 29319 36261 29331 36295
rect 29273 36255 29331 36261
rect 29454 36252 29460 36304
rect 29512 36292 29518 36304
rect 30193 36295 30251 36301
rect 30193 36292 30205 36295
rect 29512 36264 30205 36292
rect 29512 36252 29518 36264
rect 30193 36261 30205 36264
rect 30239 36261 30251 36295
rect 30193 36255 30251 36261
rect 27856 36196 28994 36224
rect 29197 36196 30328 36224
rect 27856 36184 27862 36196
rect 27430 36116 27436 36168
rect 27488 36116 27494 36168
rect 27801 36091 27859 36097
rect 27801 36088 27813 36091
rect 27264 36060 27813 36088
rect 26344 35992 26924 36020
rect 25648 35980 25654 35992
rect 26970 35980 26976 36032
rect 27028 35980 27034 36032
rect 27264 36029 27292 36060
rect 27801 36057 27813 36060
rect 27847 36057 27859 36091
rect 27801 36051 27859 36057
rect 28258 36048 28264 36100
rect 28316 36048 28322 36100
rect 27249 36023 27307 36029
rect 27249 35989 27261 36023
rect 27295 35989 27307 36023
rect 27249 35983 27307 35989
rect 28718 35980 28724 36032
rect 28776 36020 28782 36032
rect 29197 36020 29225 36196
rect 29270 36116 29276 36168
rect 29328 36116 29334 36168
rect 29362 36116 29368 36168
rect 29420 36156 29426 36168
rect 29549 36159 29607 36165
rect 29549 36156 29561 36159
rect 29420 36128 29561 36156
rect 29420 36116 29426 36128
rect 29549 36125 29561 36128
rect 29595 36125 29607 36159
rect 29549 36119 29607 36125
rect 29642 36159 29700 36165
rect 29642 36125 29654 36159
rect 29688 36125 29700 36159
rect 29642 36119 29700 36125
rect 29288 36088 29316 36116
rect 29657 36088 29685 36119
rect 29730 36116 29736 36168
rect 29788 36156 29794 36168
rect 29917 36159 29975 36165
rect 29917 36156 29929 36159
rect 29788 36128 29929 36156
rect 29788 36116 29794 36128
rect 29917 36125 29929 36128
rect 29963 36125 29975 36159
rect 29917 36119 29975 36125
rect 30006 36116 30012 36168
rect 30064 36165 30070 36168
rect 30300 36165 30328 36196
rect 32766 36184 32772 36236
rect 32824 36184 32830 36236
rect 30064 36156 30072 36165
rect 30285 36159 30343 36165
rect 30064 36128 30109 36156
rect 30064 36119 30072 36128
rect 30285 36125 30297 36159
rect 30331 36125 30343 36159
rect 30285 36119 30343 36125
rect 30064 36116 30070 36119
rect 29288 36060 29685 36088
rect 29825 36091 29883 36097
rect 29825 36057 29837 36091
rect 29871 36057 29883 36091
rect 30300 36088 30328 36119
rect 30926 36116 30932 36168
rect 30984 36116 30990 36168
rect 32217 36159 32275 36165
rect 32217 36125 32229 36159
rect 32263 36125 32275 36159
rect 32217 36119 32275 36125
rect 32309 36159 32367 36165
rect 32309 36125 32321 36159
rect 32355 36156 32367 36159
rect 32493 36159 32551 36165
rect 32493 36156 32505 36159
rect 32355 36128 32505 36156
rect 32355 36125 32367 36128
rect 32309 36119 32367 36125
rect 32493 36125 32505 36128
rect 32539 36125 32551 36159
rect 32493 36119 32551 36125
rect 32232 36088 32260 36119
rect 30300 36060 32260 36088
rect 29825 36051 29883 36057
rect 28776 35992 29225 36020
rect 28776 35980 28782 35992
rect 29362 35980 29368 36032
rect 29420 36020 29426 36032
rect 29840 36020 29868 36051
rect 29420 35992 29868 36020
rect 29420 35980 29426 35992
rect 30374 35980 30380 36032
rect 30432 35980 30438 36032
rect 30742 35980 30748 36032
rect 30800 35980 30806 36032
rect 32232 36020 32260 36060
rect 32674 36048 32680 36100
rect 32732 36088 32738 36100
rect 32732 36060 33258 36088
rect 32732 36048 32738 36060
rect 32766 36020 32772 36032
rect 32232 35992 32772 36020
rect 32766 35980 32772 35992
rect 32824 35980 32830 36032
rect 34238 35980 34244 36032
rect 34296 35980 34302 36032
rect 1104 35930 38272 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38272 35930
rect 1104 35856 38272 35878
rect 5534 35776 5540 35828
rect 5592 35776 5598 35828
rect 7190 35776 7196 35828
rect 7248 35816 7254 35828
rect 7469 35819 7527 35825
rect 7469 35816 7481 35819
rect 7248 35788 7481 35816
rect 7248 35776 7254 35788
rect 7469 35785 7481 35788
rect 7515 35785 7527 35819
rect 7469 35779 7527 35785
rect 7837 35819 7895 35825
rect 7837 35785 7849 35819
rect 7883 35785 7895 35819
rect 7837 35779 7895 35785
rect 8205 35819 8263 35825
rect 8205 35785 8217 35819
rect 8251 35816 8263 35819
rect 8662 35816 8668 35828
rect 8251 35788 8668 35816
rect 8251 35785 8263 35788
rect 8205 35779 8263 35785
rect 5626 35708 5632 35760
rect 5684 35748 5690 35760
rect 6365 35751 6423 35757
rect 6365 35748 6377 35751
rect 5684 35720 6377 35748
rect 5684 35708 5690 35720
rect 6365 35717 6377 35720
rect 6411 35748 6423 35751
rect 6454 35748 6460 35760
rect 6411 35720 6460 35748
rect 6411 35717 6423 35720
rect 6365 35711 6423 35717
rect 6454 35708 6460 35720
rect 6512 35708 6518 35760
rect 5718 35640 5724 35692
rect 5776 35640 5782 35692
rect 7653 35683 7711 35689
rect 7653 35649 7665 35683
rect 7699 35680 7711 35683
rect 7852 35680 7880 35779
rect 8662 35776 8668 35788
rect 8720 35776 8726 35828
rect 8938 35776 8944 35828
rect 8996 35816 9002 35828
rect 9125 35819 9183 35825
rect 9125 35816 9137 35819
rect 8996 35788 9137 35816
rect 8996 35776 9002 35788
rect 9125 35785 9137 35788
rect 9171 35785 9183 35819
rect 9125 35779 9183 35785
rect 9214 35776 9220 35828
rect 9272 35816 9278 35828
rect 9309 35819 9367 35825
rect 9309 35816 9321 35819
rect 9272 35788 9321 35816
rect 9272 35776 9278 35788
rect 9309 35785 9321 35788
rect 9355 35785 9367 35819
rect 9309 35779 9367 35785
rect 10229 35819 10287 35825
rect 10229 35785 10241 35819
rect 10275 35816 10287 35819
rect 10686 35816 10692 35828
rect 10275 35788 10692 35816
rect 10275 35785 10287 35788
rect 10229 35779 10287 35785
rect 10686 35776 10692 35788
rect 10744 35776 10750 35828
rect 13541 35819 13599 35825
rect 13541 35785 13553 35819
rect 13587 35816 13599 35819
rect 13630 35816 13636 35828
rect 13587 35788 13636 35816
rect 13587 35785 13599 35788
rect 13541 35779 13599 35785
rect 13630 35776 13636 35788
rect 13688 35776 13694 35828
rect 14829 35819 14887 35825
rect 14829 35785 14841 35819
rect 14875 35816 14887 35819
rect 15562 35816 15568 35828
rect 14875 35788 15568 35816
rect 14875 35785 14887 35788
rect 14829 35779 14887 35785
rect 15562 35776 15568 35788
rect 15620 35776 15626 35828
rect 17126 35776 17132 35828
rect 17184 35816 17190 35828
rect 18690 35816 18696 35828
rect 17184 35788 18696 35816
rect 17184 35776 17190 35788
rect 18690 35776 18696 35788
rect 18748 35776 18754 35828
rect 22738 35816 22744 35828
rect 21560 35788 22744 35816
rect 8478 35748 8484 35760
rect 7699 35652 7880 35680
rect 8220 35720 8484 35748
rect 7699 35649 7711 35652
rect 7653 35643 7711 35649
rect 6822 35572 6828 35624
rect 6880 35612 6886 35624
rect 7193 35615 7251 35621
rect 7193 35612 7205 35615
rect 6880 35584 7205 35612
rect 6880 35572 6886 35584
rect 7193 35581 7205 35584
rect 7239 35612 7251 35615
rect 8220 35612 8248 35720
rect 8478 35708 8484 35720
rect 8536 35708 8542 35760
rect 9048 35720 9996 35748
rect 9048 35689 9076 35720
rect 9968 35692 9996 35720
rect 11974 35708 11980 35760
rect 12032 35748 12038 35760
rect 20898 35748 20904 35760
rect 12032 35720 20904 35748
rect 12032 35708 12038 35720
rect 20898 35708 20904 35720
rect 20956 35748 20962 35760
rect 21560 35748 21588 35788
rect 22738 35776 22744 35788
rect 22796 35816 22802 35828
rect 22796 35788 23336 35816
rect 22796 35776 22802 35788
rect 20956 35720 21588 35748
rect 20956 35708 20962 35720
rect 21634 35708 21640 35760
rect 21692 35748 21698 35760
rect 21910 35748 21916 35760
rect 21692 35720 21916 35748
rect 21692 35708 21698 35720
rect 21910 35708 21916 35720
rect 21968 35748 21974 35760
rect 21968 35720 23249 35748
rect 21968 35708 21974 35720
rect 8297 35683 8355 35689
rect 8297 35649 8309 35683
rect 8343 35680 8355 35683
rect 9033 35683 9091 35689
rect 8343 35652 8984 35680
rect 8343 35649 8355 35652
rect 8297 35643 8355 35649
rect 8956 35624 8984 35652
rect 9033 35649 9045 35683
rect 9079 35649 9091 35683
rect 9033 35643 9091 35649
rect 9493 35683 9551 35689
rect 9493 35649 9505 35683
rect 9539 35680 9551 35683
rect 9539 35652 9812 35680
rect 9539 35649 9551 35652
rect 9493 35643 9551 35649
rect 7239 35584 8248 35612
rect 8389 35615 8447 35621
rect 7239 35581 7251 35584
rect 7193 35575 7251 35581
rect 8389 35581 8401 35615
rect 8435 35581 8447 35615
rect 8389 35575 8447 35581
rect 8404 35544 8432 35575
rect 8938 35572 8944 35624
rect 8996 35572 9002 35624
rect 9784 35553 9812 35652
rect 9950 35640 9956 35692
rect 10008 35640 10014 35692
rect 10137 35683 10195 35689
rect 10137 35649 10149 35683
rect 10183 35649 10195 35683
rect 10137 35643 10195 35649
rect 10781 35683 10839 35689
rect 10781 35649 10793 35683
rect 10827 35680 10839 35683
rect 10827 35652 11560 35680
rect 10827 35649 10839 35652
rect 10781 35643 10839 35649
rect 8220 35516 8432 35544
rect 9769 35547 9827 35553
rect 8220 35488 8248 35516
rect 9769 35513 9781 35547
rect 9815 35513 9827 35547
rect 10152 35544 10180 35643
rect 10413 35615 10471 35621
rect 10413 35581 10425 35615
rect 10459 35612 10471 35615
rect 10459 35584 11468 35612
rect 10459 35581 10471 35584
rect 10413 35575 10471 35581
rect 10778 35544 10784 35556
rect 10152 35516 10784 35544
rect 9769 35507 9827 35513
rect 10778 35504 10784 35516
rect 10836 35504 10842 35556
rect 8202 35436 8208 35488
rect 8260 35436 8266 35488
rect 10594 35436 10600 35488
rect 10652 35436 10658 35488
rect 11440 35476 11468 35584
rect 11532 35553 11560 35652
rect 11790 35640 11796 35692
rect 11848 35680 11854 35692
rect 11885 35683 11943 35689
rect 11885 35680 11897 35683
rect 11848 35652 11897 35680
rect 11848 35640 11854 35652
rect 11885 35649 11897 35652
rect 11931 35649 11943 35683
rect 11885 35643 11943 35649
rect 12802 35640 12808 35692
rect 12860 35680 12866 35692
rect 12897 35683 12955 35689
rect 12897 35680 12909 35683
rect 12860 35652 12909 35680
rect 12860 35640 12866 35652
rect 12897 35649 12909 35652
rect 12943 35649 12955 35683
rect 12897 35643 12955 35649
rect 12986 35640 12992 35692
rect 13044 35680 13050 35692
rect 13170 35689 13176 35692
rect 13127 35683 13176 35689
rect 13044 35652 13089 35680
rect 13044 35640 13050 35652
rect 13127 35649 13139 35683
rect 13173 35649 13176 35683
rect 13127 35643 13176 35649
rect 13170 35640 13176 35643
rect 13228 35640 13234 35692
rect 13262 35640 13268 35692
rect 13320 35640 13326 35692
rect 13354 35640 13360 35692
rect 13412 35689 13418 35692
rect 13412 35680 13420 35689
rect 13412 35652 13457 35680
rect 13412 35643 13420 35652
rect 13412 35640 13418 35643
rect 14182 35640 14188 35692
rect 14240 35680 14246 35692
rect 14737 35683 14795 35689
rect 14737 35680 14749 35683
rect 14240 35652 14749 35680
rect 14240 35640 14246 35652
rect 14737 35649 14749 35652
rect 14783 35649 14795 35683
rect 14737 35643 14795 35649
rect 18598 35640 18604 35692
rect 18656 35680 18662 35692
rect 21726 35680 21732 35692
rect 18656 35652 21732 35680
rect 18656 35640 18662 35652
rect 21726 35640 21732 35652
rect 21784 35640 21790 35692
rect 21818 35640 21824 35692
rect 21876 35680 21882 35692
rect 22097 35683 22155 35689
rect 22097 35680 22109 35683
rect 21876 35652 22109 35680
rect 21876 35640 21882 35652
rect 22097 35649 22109 35652
rect 22143 35680 22155 35683
rect 22186 35680 22192 35692
rect 22143 35652 22192 35680
rect 22143 35649 22155 35652
rect 22097 35643 22155 35649
rect 22186 35640 22192 35652
rect 22244 35640 22250 35692
rect 22281 35683 22339 35689
rect 22281 35649 22293 35683
rect 22327 35649 22339 35683
rect 22281 35643 22339 35649
rect 12161 35615 12219 35621
rect 12161 35581 12173 35615
rect 12207 35612 12219 35615
rect 12250 35612 12256 35624
rect 12207 35584 12256 35612
rect 12207 35581 12219 35584
rect 12161 35575 12219 35581
rect 11517 35547 11575 35553
rect 11517 35513 11529 35547
rect 11563 35513 11575 35547
rect 11517 35507 11575 35513
rect 12176 35476 12204 35575
rect 12250 35572 12256 35584
rect 12308 35572 12314 35624
rect 22296 35612 22324 35643
rect 22370 35640 22376 35692
rect 22428 35640 22434 35692
rect 22465 35683 22523 35689
rect 22465 35649 22477 35683
rect 22511 35680 22523 35683
rect 22554 35680 22560 35692
rect 22511 35652 22560 35680
rect 22511 35649 22523 35652
rect 22465 35643 22523 35649
rect 22554 35640 22560 35652
rect 22612 35640 22618 35692
rect 22741 35683 22799 35689
rect 22741 35649 22753 35683
rect 22787 35649 22799 35683
rect 22741 35643 22799 35649
rect 22756 35612 22784 35643
rect 22830 35640 22836 35692
rect 22888 35680 22894 35692
rect 23221 35689 23249 35720
rect 23017 35683 23075 35689
rect 22888 35652 22933 35680
rect 22888 35640 22894 35652
rect 23017 35649 23029 35683
rect 23063 35649 23075 35683
rect 23017 35643 23075 35649
rect 23109 35683 23167 35689
rect 23109 35649 23121 35683
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 23206 35683 23264 35689
rect 23206 35649 23218 35683
rect 23252 35649 23264 35683
rect 23206 35643 23264 35649
rect 21836 35584 22324 35612
rect 22388 35584 22784 35612
rect 21836 35488 21864 35584
rect 22388 35488 22416 35584
rect 23032 35544 23060 35643
rect 23124 35612 23152 35643
rect 23308 35612 23336 35788
rect 25774 35776 25780 35828
rect 25832 35776 25838 35828
rect 27249 35819 27307 35825
rect 27249 35785 27261 35819
rect 27295 35816 27307 35819
rect 27430 35816 27436 35828
rect 27295 35788 27436 35816
rect 27295 35785 27307 35788
rect 27249 35779 27307 35785
rect 27430 35776 27436 35788
rect 27488 35776 27494 35828
rect 32674 35816 32680 35828
rect 31496 35788 32680 35816
rect 25225 35751 25283 35757
rect 25225 35717 25237 35751
rect 25271 35748 25283 35751
rect 25590 35748 25596 35760
rect 25271 35720 25596 35748
rect 25271 35717 25283 35720
rect 25225 35711 25283 35717
rect 25590 35708 25596 35720
rect 25648 35708 25654 35760
rect 25792 35748 25820 35776
rect 25700 35720 25820 35748
rect 25700 35689 25728 35720
rect 26142 35708 26148 35760
rect 26200 35748 26206 35760
rect 29641 35751 29699 35757
rect 29641 35748 29653 35751
rect 26200 35720 29653 35748
rect 26200 35708 26206 35720
rect 29641 35717 29653 35720
rect 29687 35748 29699 35751
rect 30374 35748 30380 35760
rect 29687 35720 30057 35748
rect 29687 35717 29699 35720
rect 29641 35711 29699 35717
rect 25409 35683 25467 35689
rect 25409 35680 25421 35683
rect 25332 35652 25421 35680
rect 23566 35612 23572 35624
rect 23124 35584 23572 35612
rect 23566 35572 23572 35584
rect 23624 35572 23630 35624
rect 25332 35556 25360 35652
rect 25409 35649 25421 35652
rect 25455 35649 25467 35683
rect 25409 35643 25467 35649
rect 25501 35683 25559 35689
rect 25501 35649 25513 35683
rect 25547 35649 25559 35683
rect 25501 35643 25559 35649
rect 25685 35683 25743 35689
rect 25685 35649 25697 35683
rect 25731 35649 25743 35683
rect 25685 35643 25743 35649
rect 25516 35556 25544 35643
rect 25774 35640 25780 35692
rect 25832 35680 25838 35692
rect 26050 35680 26056 35692
rect 25832 35652 26056 35680
rect 25832 35640 25838 35652
rect 26050 35640 26056 35652
rect 26108 35640 26114 35692
rect 26234 35640 26240 35692
rect 26292 35640 26298 35692
rect 27338 35640 27344 35692
rect 27396 35680 27402 35692
rect 27617 35683 27675 35689
rect 27617 35680 27629 35683
rect 27396 35652 27629 35680
rect 27396 35640 27402 35652
rect 27617 35649 27629 35652
rect 27663 35649 27675 35683
rect 29178 35680 29184 35692
rect 29104 35670 29184 35680
rect 27617 35643 27675 35649
rect 28966 35652 29184 35670
rect 28966 35642 29132 35652
rect 26252 35612 26280 35640
rect 27430 35612 27436 35624
rect 26252 35584 27436 35612
rect 27430 35572 27436 35584
rect 27488 35612 27494 35624
rect 27709 35615 27767 35621
rect 27709 35612 27721 35615
rect 27488 35584 27721 35612
rect 27488 35572 27494 35584
rect 27709 35581 27721 35584
rect 27755 35612 27767 35615
rect 27798 35612 27804 35624
rect 27755 35584 27804 35612
rect 27755 35581 27767 35584
rect 27709 35575 27767 35581
rect 27798 35572 27804 35584
rect 27856 35572 27862 35624
rect 27893 35615 27951 35621
rect 27893 35581 27905 35615
rect 27939 35612 27951 35615
rect 28966 35612 28994 35642
rect 29178 35640 29184 35652
rect 29236 35640 29242 35692
rect 29454 35640 29460 35692
rect 29512 35640 29518 35692
rect 29546 35640 29552 35692
rect 29604 35680 29610 35692
rect 29733 35683 29791 35689
rect 29733 35680 29745 35683
rect 29604 35652 29745 35680
rect 29604 35640 29610 35652
rect 29733 35649 29745 35652
rect 29779 35649 29791 35683
rect 29733 35643 29791 35649
rect 27939 35584 28994 35612
rect 27939 35581 27951 35584
rect 27893 35575 27951 35581
rect 22756 35516 23060 35544
rect 22756 35488 22784 35516
rect 23106 35504 23112 35556
rect 23164 35544 23170 35556
rect 24026 35544 24032 35556
rect 23164 35516 24032 35544
rect 23164 35504 23170 35516
rect 24026 35504 24032 35516
rect 24084 35504 24090 35556
rect 25314 35504 25320 35556
rect 25372 35504 25378 35556
rect 25498 35504 25504 35556
rect 25556 35544 25562 35556
rect 28994 35544 29000 35556
rect 25556 35516 29000 35544
rect 25556 35504 25562 35516
rect 28994 35504 29000 35516
rect 29052 35504 29058 35556
rect 29197 35516 29408 35544
rect 11440 35448 12204 35476
rect 12710 35436 12716 35488
rect 12768 35476 12774 35488
rect 13354 35476 13360 35488
rect 12768 35448 13360 35476
rect 12768 35436 12774 35448
rect 13354 35436 13360 35448
rect 13412 35436 13418 35488
rect 21818 35436 21824 35488
rect 21876 35436 21882 35488
rect 22370 35436 22376 35488
rect 22428 35436 22434 35488
rect 22646 35436 22652 35488
rect 22704 35436 22710 35488
rect 22738 35436 22744 35488
rect 22796 35436 22802 35488
rect 23382 35436 23388 35488
rect 23440 35436 23446 35488
rect 24578 35436 24584 35488
rect 24636 35476 24642 35488
rect 26510 35476 26516 35488
rect 24636 35448 26516 35476
rect 24636 35436 24642 35448
rect 26510 35436 26516 35448
rect 26568 35476 26574 35488
rect 29197 35476 29225 35516
rect 29380 35488 29408 35516
rect 26568 35448 29225 35476
rect 26568 35436 26574 35448
rect 29270 35436 29276 35488
rect 29328 35436 29334 35488
rect 29362 35436 29368 35488
rect 29420 35436 29426 35488
rect 30029 35476 30057 35720
rect 30116 35720 30380 35748
rect 30116 35689 30144 35720
rect 30374 35708 30380 35720
rect 30432 35708 30438 35760
rect 30466 35708 30472 35760
rect 30524 35748 30530 35760
rect 30834 35748 30840 35760
rect 30524 35720 30840 35748
rect 30524 35708 30530 35720
rect 30834 35708 30840 35720
rect 30892 35708 30898 35760
rect 30101 35683 30159 35689
rect 30101 35649 30113 35683
rect 30147 35649 30159 35683
rect 30101 35643 30159 35649
rect 30377 35615 30435 35621
rect 30377 35581 30389 35615
rect 30423 35612 30435 35615
rect 30742 35612 30748 35624
rect 30423 35584 30748 35612
rect 30423 35581 30435 35584
rect 30377 35575 30435 35581
rect 30742 35572 30748 35584
rect 30800 35572 30806 35624
rect 30834 35572 30840 35624
rect 30892 35612 30898 35624
rect 31496 35612 31524 35788
rect 32674 35776 32680 35788
rect 32732 35776 32738 35828
rect 32769 35819 32827 35825
rect 32769 35785 32781 35819
rect 32815 35816 32827 35819
rect 32950 35816 32956 35828
rect 32815 35788 32956 35816
rect 32815 35785 32827 35788
rect 32769 35779 32827 35785
rect 32950 35776 32956 35788
rect 33008 35776 33014 35828
rect 33134 35776 33140 35828
rect 33192 35776 33198 35828
rect 33229 35819 33287 35825
rect 33229 35785 33241 35819
rect 33275 35816 33287 35819
rect 34238 35816 34244 35828
rect 33275 35788 34244 35816
rect 33275 35785 33287 35788
rect 33229 35779 33287 35785
rect 30892 35584 31524 35612
rect 30892 35572 30898 35584
rect 33244 35544 33272 35779
rect 34238 35776 34244 35788
rect 34296 35776 34302 35828
rect 33318 35572 33324 35624
rect 33376 35572 33382 35624
rect 31404 35516 33272 35544
rect 31404 35476 31432 35516
rect 30029 35448 31432 35476
rect 31846 35436 31852 35488
rect 31904 35436 31910 35488
rect 1104 35386 38272 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38272 35386
rect 1104 35312 38272 35334
rect 5718 35232 5724 35284
rect 5776 35272 5782 35284
rect 5997 35275 6055 35281
rect 5997 35272 6009 35275
rect 5776 35244 6009 35272
rect 5776 35232 5782 35244
rect 5997 35241 6009 35244
rect 6043 35241 6055 35275
rect 5997 35235 6055 35241
rect 8662 35232 8668 35284
rect 8720 35272 8726 35284
rect 11882 35272 11888 35284
rect 8720 35244 11888 35272
rect 8720 35232 8726 35244
rect 11882 35232 11888 35244
rect 11940 35232 11946 35284
rect 11974 35232 11980 35284
rect 12032 35232 12038 35284
rect 12066 35232 12072 35284
rect 12124 35272 12130 35284
rect 12124 35244 21404 35272
rect 12124 35232 12130 35244
rect 11900 35204 11928 35232
rect 14093 35207 14151 35213
rect 14093 35204 14105 35207
rect 11900 35176 14105 35204
rect 14093 35173 14105 35176
rect 14139 35204 14151 35207
rect 17494 35204 17500 35216
rect 14139 35176 17500 35204
rect 14139 35173 14151 35176
rect 14093 35167 14151 35173
rect 17494 35164 17500 35176
rect 17552 35164 17558 35216
rect 20714 35204 20720 35216
rect 18984 35176 20720 35204
rect 6546 35096 6552 35148
rect 6604 35096 6610 35148
rect 10505 35139 10563 35145
rect 10505 35105 10517 35139
rect 10551 35136 10563 35139
rect 10594 35136 10600 35148
rect 10551 35108 10600 35136
rect 10551 35105 10563 35108
rect 10505 35099 10563 35105
rect 10594 35096 10600 35108
rect 10652 35096 10658 35148
rect 17402 35096 17408 35148
rect 17460 35136 17466 35148
rect 18984 35136 19012 35176
rect 20714 35164 20720 35176
rect 20772 35164 20778 35216
rect 20898 35164 20904 35216
rect 20956 35164 20962 35216
rect 20916 35136 20944 35164
rect 17460 35108 19012 35136
rect 19352 35108 19656 35136
rect 20916 35108 21129 35136
rect 17460 35096 17466 35108
rect 19352 35080 19380 35108
rect 4433 35071 4491 35077
rect 4433 35037 4445 35071
rect 4479 35068 4491 35071
rect 5442 35068 5448 35080
rect 4479 35040 5448 35068
rect 4479 35037 4491 35040
rect 4433 35031 4491 35037
rect 5442 35028 5448 35040
rect 5500 35068 5506 35080
rect 7929 35071 7987 35077
rect 7929 35068 7941 35071
rect 5500 35040 7941 35068
rect 5500 35028 5506 35040
rect 7929 35037 7941 35040
rect 7975 35068 7987 35071
rect 9950 35068 9956 35080
rect 7975 35040 9956 35068
rect 7975 35037 7987 35040
rect 7929 35031 7987 35037
rect 9950 35028 9956 35040
rect 10008 35028 10014 35080
rect 10045 35071 10103 35077
rect 10045 35037 10057 35071
rect 10091 35068 10103 35071
rect 10229 35071 10287 35077
rect 10229 35068 10241 35071
rect 10091 35040 10241 35068
rect 10091 35037 10103 35040
rect 10045 35031 10103 35037
rect 10229 35037 10241 35040
rect 10275 35037 10287 35071
rect 10229 35031 10287 35037
rect 14277 35071 14335 35077
rect 14277 35037 14289 35071
rect 14323 35068 14335 35071
rect 14366 35068 14372 35080
rect 14323 35040 14372 35068
rect 14323 35037 14335 35040
rect 14277 35031 14335 35037
rect 14366 35028 14372 35040
rect 14424 35028 14430 35080
rect 14461 35071 14519 35077
rect 14461 35037 14473 35071
rect 14507 35068 14519 35071
rect 14826 35068 14832 35080
rect 14507 35040 14832 35068
rect 14507 35037 14519 35040
rect 14461 35031 14519 35037
rect 14826 35028 14832 35040
rect 14884 35068 14890 35080
rect 14884 35040 15424 35068
rect 14884 35028 14890 35040
rect 6365 35003 6423 35009
rect 6365 34969 6377 35003
rect 6411 35000 6423 35003
rect 6730 35000 6736 35012
rect 6411 34972 6736 35000
rect 6411 34969 6423 34972
rect 6365 34963 6423 34969
rect 6730 34960 6736 34972
rect 6788 35000 6794 35012
rect 9968 35000 9996 35028
rect 6788 34972 9444 35000
rect 9968 34972 10272 35000
rect 6788 34960 6794 34972
rect 9416 34944 9444 34972
rect 10244 34944 10272 34972
rect 10704 34972 10994 35000
rect 10704 34944 10732 34972
rect 15396 34944 15424 35040
rect 19334 35028 19340 35080
rect 19392 35028 19398 35080
rect 19426 35028 19432 35080
rect 19484 35028 19490 35080
rect 19628 35077 19656 35108
rect 19613 35071 19671 35077
rect 19613 35037 19625 35071
rect 19659 35037 19671 35071
rect 19613 35031 19671 35037
rect 19889 35071 19947 35077
rect 19889 35037 19901 35071
rect 19935 35068 19947 35071
rect 19978 35068 19984 35080
rect 19935 35040 19984 35068
rect 19935 35037 19947 35040
rect 19889 35031 19947 35037
rect 19978 35028 19984 35040
rect 20036 35068 20042 35080
rect 20898 35068 20904 35080
rect 20036 35040 20904 35068
rect 20036 35028 20042 35040
rect 20898 35028 20904 35040
rect 20956 35028 20962 35080
rect 20990 35028 20996 35080
rect 21048 35028 21054 35080
rect 21101 35077 21129 35108
rect 21376 35077 21404 35244
rect 22186 35232 22192 35284
rect 22244 35232 22250 35284
rect 22646 35232 22652 35284
rect 22704 35232 22710 35284
rect 27246 35232 27252 35284
rect 27304 35272 27310 35284
rect 27801 35275 27859 35281
rect 27801 35272 27813 35275
rect 27304 35244 27813 35272
rect 27304 35232 27310 35244
rect 27801 35241 27813 35244
rect 27847 35241 27859 35275
rect 27801 35235 27859 35241
rect 28258 35232 28264 35284
rect 28316 35272 28322 35284
rect 30466 35272 30472 35284
rect 28316 35244 30472 35272
rect 28316 35232 28322 35244
rect 30466 35232 30472 35244
rect 30524 35232 30530 35284
rect 30653 35275 30711 35281
rect 30653 35241 30665 35275
rect 30699 35272 30711 35275
rect 30926 35272 30932 35284
rect 30699 35244 30932 35272
rect 30699 35241 30711 35244
rect 30653 35235 30711 35241
rect 30926 35232 30932 35244
rect 30984 35232 30990 35284
rect 22204 35204 22232 35232
rect 22204 35176 22508 35204
rect 21086 35071 21144 35077
rect 21086 35037 21098 35071
rect 21132 35037 21144 35071
rect 21086 35031 21144 35037
rect 21361 35071 21419 35077
rect 21361 35037 21373 35071
rect 21407 35037 21419 35071
rect 21361 35031 21419 35037
rect 19521 35003 19579 35009
rect 19521 34969 19533 35003
rect 19567 34969 19579 35003
rect 19521 34963 19579 34969
rect 19751 35003 19809 35009
rect 19751 34969 19763 35003
rect 19797 35000 19809 35003
rect 21174 35000 21180 35012
rect 19797 34972 21180 35000
rect 19797 34969 19809 34972
rect 19751 34963 19809 34969
rect 4522 34892 4528 34944
rect 4580 34892 4586 34944
rect 6454 34892 6460 34944
rect 6512 34892 6518 34944
rect 8018 34892 8024 34944
rect 8076 34892 8082 34944
rect 9398 34892 9404 34944
rect 9456 34892 9462 34944
rect 10226 34892 10232 34944
rect 10284 34892 10290 34944
rect 10686 34892 10692 34944
rect 10744 34892 10750 34944
rect 10870 34892 10876 34944
rect 10928 34932 10934 34944
rect 11974 34932 11980 34944
rect 10928 34904 11980 34932
rect 10928 34892 10934 34904
rect 11974 34892 11980 34904
rect 12032 34892 12038 34944
rect 14369 34935 14427 34941
rect 14369 34901 14381 34935
rect 14415 34932 14427 34935
rect 14458 34932 14464 34944
rect 14415 34904 14464 34932
rect 14415 34901 14427 34904
rect 14369 34895 14427 34901
rect 14458 34892 14464 34904
rect 14516 34892 14522 34944
rect 14642 34892 14648 34944
rect 14700 34892 14706 34944
rect 15378 34892 15384 34944
rect 15436 34892 15442 34944
rect 18230 34892 18236 34944
rect 18288 34932 18294 34944
rect 19245 34935 19303 34941
rect 19245 34932 19257 34935
rect 18288 34904 19257 34932
rect 18288 34892 18294 34904
rect 19245 34901 19257 34904
rect 19291 34901 19303 34935
rect 19536 34932 19564 34963
rect 21174 34960 21180 34972
rect 21232 34960 21238 35012
rect 21266 34960 21272 35012
rect 21324 34960 21330 35012
rect 21376 35000 21404 35031
rect 21450 35028 21456 35080
rect 21508 35077 21514 35080
rect 21508 35068 21516 35077
rect 21508 35040 21553 35068
rect 21508 35031 21516 35040
rect 21508 35028 21514 35031
rect 21634 35028 21640 35080
rect 21692 35068 21698 35080
rect 22189 35071 22247 35077
rect 22189 35068 22201 35071
rect 21692 35040 22201 35068
rect 21692 35028 21698 35040
rect 22189 35037 22201 35040
rect 22235 35037 22247 35071
rect 22189 35031 22247 35037
rect 22278 35028 22284 35080
rect 22336 35068 22342 35080
rect 22480 35077 22508 35176
rect 22664 35136 22692 35232
rect 23382 35164 23388 35216
rect 23440 35204 23446 35216
rect 23440 35176 23520 35204
rect 23440 35164 23446 35176
rect 23492 35145 23520 35176
rect 25406 35164 25412 35216
rect 25464 35164 25470 35216
rect 25590 35164 25596 35216
rect 25648 35164 25654 35216
rect 23477 35139 23535 35145
rect 22664 35108 23336 35136
rect 22465 35071 22523 35077
rect 22336 35040 22381 35068
rect 22336 35028 22342 35040
rect 22465 35037 22477 35071
rect 22511 35037 22523 35071
rect 22465 35031 22523 35037
rect 22695 35071 22753 35077
rect 22695 35037 22707 35071
rect 22741 35068 22753 35071
rect 23106 35068 23112 35080
rect 22741 35040 23112 35068
rect 22741 35037 22753 35040
rect 22695 35031 22753 35037
rect 23106 35028 23112 35040
rect 23164 35028 23170 35080
rect 23308 35077 23336 35108
rect 23477 35105 23489 35139
rect 23523 35105 23535 35139
rect 23477 35099 23535 35105
rect 23569 35139 23627 35145
rect 23569 35105 23581 35139
rect 23615 35136 23627 35139
rect 24210 35136 24216 35148
rect 23615 35108 24216 35136
rect 23615 35105 23627 35108
rect 23569 35099 23627 35105
rect 24210 35096 24216 35108
rect 24268 35136 24274 35148
rect 25608 35136 25636 35164
rect 27157 35139 27215 35145
rect 24268 35108 25544 35136
rect 25608 35108 25912 35136
rect 24268 35096 24274 35108
rect 23293 35071 23351 35077
rect 23293 35037 23305 35071
rect 23339 35037 23351 35071
rect 23293 35031 23351 35037
rect 23382 35028 23388 35080
rect 23440 35028 23446 35080
rect 23753 35071 23811 35077
rect 23753 35037 23765 35071
rect 23799 35037 23811 35071
rect 23753 35031 23811 35037
rect 22557 35003 22615 35009
rect 22557 35000 22569 35003
rect 21376 34972 22569 35000
rect 22557 34969 22569 34972
rect 22603 35000 22615 35003
rect 22922 35000 22928 35012
rect 22603 34972 22928 35000
rect 22603 34969 22615 34972
rect 22557 34963 22615 34969
rect 22922 34960 22928 34972
rect 22980 34960 22986 35012
rect 19978 34932 19984 34944
rect 19536 34904 19984 34932
rect 19245 34895 19303 34901
rect 19978 34892 19984 34904
rect 20036 34892 20042 34944
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 21284 34932 21312 34960
rect 23768 34944 23796 35031
rect 24854 35028 24860 35080
rect 24912 35068 24918 35080
rect 24949 35071 25007 35077
rect 24949 35068 24961 35071
rect 24912 35040 24961 35068
rect 24912 35028 24918 35040
rect 24949 35037 24961 35040
rect 24995 35037 25007 35071
rect 24949 35031 25007 35037
rect 25041 35071 25099 35077
rect 25041 35037 25053 35071
rect 25087 35037 25099 35071
rect 25041 35031 25099 35037
rect 25056 35000 25084 35031
rect 25130 35028 25136 35080
rect 25188 35028 25194 35080
rect 25317 35071 25375 35077
rect 25317 35037 25329 35071
rect 25363 35037 25375 35071
rect 25516 35068 25544 35108
rect 25685 35071 25743 35077
rect 25685 35068 25697 35071
rect 25516 35040 25697 35068
rect 25317 35031 25375 35037
rect 25685 35037 25697 35040
rect 25731 35037 25743 35071
rect 25685 35031 25743 35037
rect 24964 34972 25084 35000
rect 25332 35000 25360 35031
rect 25774 35028 25780 35080
rect 25832 35028 25838 35080
rect 25884 35077 25912 35108
rect 27157 35105 27169 35139
rect 27203 35136 27215 35139
rect 28258 35136 28264 35148
rect 27203 35108 28264 35136
rect 27203 35105 27215 35108
rect 27157 35099 27215 35105
rect 28258 35096 28264 35108
rect 28316 35096 28322 35148
rect 31294 35096 31300 35148
rect 31352 35136 31358 35148
rect 33686 35136 33692 35148
rect 31352 35108 33692 35136
rect 31352 35096 31358 35108
rect 33686 35096 33692 35108
rect 33744 35096 33750 35148
rect 25869 35071 25927 35077
rect 25869 35037 25881 35071
rect 25915 35037 25927 35071
rect 25869 35031 25927 35037
rect 26053 35071 26111 35077
rect 26053 35037 26065 35071
rect 26099 35037 26111 35071
rect 26053 35031 26111 35037
rect 25590 35000 25596 35012
rect 25332 34972 25596 35000
rect 24964 34944 24992 34972
rect 25590 34960 25596 34972
rect 25648 35000 25654 35012
rect 26068 35000 26096 35031
rect 26970 35028 26976 35080
rect 27028 35068 27034 35080
rect 27341 35071 27399 35077
rect 27341 35068 27353 35071
rect 27028 35040 27353 35068
rect 27028 35028 27034 35040
rect 27341 35037 27353 35040
rect 27387 35037 27399 35071
rect 27341 35031 27399 35037
rect 27430 35028 27436 35080
rect 27488 35068 27494 35080
rect 27525 35071 27583 35077
rect 27525 35068 27537 35071
rect 27488 35040 27537 35068
rect 27488 35028 27494 35040
rect 27525 35037 27537 35040
rect 27571 35037 27583 35071
rect 27525 35031 27583 35037
rect 27614 35049 27672 35055
rect 27614 35015 27626 35049
rect 27660 35015 27672 35049
rect 27706 35028 27712 35080
rect 27764 35028 27770 35080
rect 29454 35028 29460 35080
rect 29512 35068 29518 35080
rect 31021 35071 31079 35077
rect 31021 35068 31033 35071
rect 29512 35040 31033 35068
rect 29512 35028 29518 35040
rect 31021 35037 31033 35040
rect 31067 35068 31079 35071
rect 31846 35068 31852 35080
rect 31067 35040 31852 35068
rect 31067 35037 31079 35040
rect 31021 35031 31079 35037
rect 31846 35028 31852 35040
rect 31904 35028 31910 35080
rect 27614 35009 27672 35015
rect 25648 34972 26096 35000
rect 25648 34960 25654 34972
rect 20772 34904 21312 34932
rect 21637 34935 21695 34941
rect 20772 34892 20778 34904
rect 21637 34901 21649 34935
rect 21683 34932 21695 34935
rect 22278 34932 22284 34944
rect 21683 34904 22284 34932
rect 21683 34901 21695 34904
rect 21637 34895 21695 34901
rect 22278 34892 22284 34904
rect 22336 34892 22342 34944
rect 22830 34892 22836 34944
rect 22888 34892 22894 34944
rect 23106 34892 23112 34944
rect 23164 34892 23170 34944
rect 23198 34892 23204 34944
rect 23256 34932 23262 34944
rect 23382 34932 23388 34944
rect 23256 34904 23388 34932
rect 23256 34892 23262 34904
rect 23382 34892 23388 34904
rect 23440 34892 23446 34944
rect 23750 34892 23756 34944
rect 23808 34892 23814 34944
rect 24673 34935 24731 34941
rect 24673 34901 24685 34935
rect 24719 34932 24731 34935
rect 24762 34932 24768 34944
rect 24719 34904 24768 34932
rect 24719 34901 24731 34904
rect 24673 34895 24731 34901
rect 24762 34892 24768 34904
rect 24820 34892 24826 34944
rect 24946 34892 24952 34944
rect 25004 34892 25010 34944
rect 25038 34892 25044 34944
rect 25096 34932 25102 34944
rect 27632 34932 27660 35009
rect 29546 35000 29552 35012
rect 29380 34972 29552 35000
rect 29380 34932 29408 34972
rect 29546 34960 29552 34972
rect 29604 34960 29610 35012
rect 25096 34904 29408 34932
rect 25096 34892 25102 34904
rect 31110 34892 31116 34944
rect 31168 34892 31174 34944
rect 1104 34842 38272 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38272 34842
rect 1104 34768 38272 34790
rect 4522 34688 4528 34740
rect 4580 34688 4586 34740
rect 6454 34688 6460 34740
rect 6512 34728 6518 34740
rect 6733 34731 6791 34737
rect 6733 34728 6745 34731
rect 6512 34700 6745 34728
rect 6512 34688 6518 34700
rect 6733 34697 6745 34700
rect 6779 34728 6791 34731
rect 8938 34728 8944 34740
rect 6779 34700 8944 34728
rect 6779 34697 6791 34700
rect 6733 34691 6791 34697
rect 8938 34688 8944 34700
rect 8996 34688 9002 34740
rect 9585 34731 9643 34737
rect 9585 34697 9597 34731
rect 9631 34728 9643 34731
rect 9674 34728 9680 34740
rect 9631 34700 9680 34728
rect 9631 34697 9643 34700
rect 9585 34691 9643 34697
rect 9674 34688 9680 34700
rect 9732 34728 9738 34740
rect 10870 34728 10876 34740
rect 9732 34700 10876 34728
rect 9732 34688 9738 34700
rect 10870 34688 10876 34700
rect 10928 34688 10934 34740
rect 16853 34731 16911 34737
rect 10980 34700 12572 34728
rect 4540 34660 4568 34688
rect 8018 34660 8024 34672
rect 4356 34632 4568 34660
rect 7852 34632 8024 34660
rect 4356 34601 4384 34632
rect 4341 34595 4399 34601
rect 4341 34561 4353 34595
rect 4387 34561 4399 34595
rect 6730 34592 6736 34604
rect 5750 34564 6736 34592
rect 4341 34555 4399 34561
rect 6730 34552 6736 34564
rect 6788 34552 6794 34604
rect 7852 34601 7880 34632
rect 8018 34620 8024 34632
rect 8076 34620 8082 34672
rect 9398 34620 9404 34672
rect 9456 34660 9462 34672
rect 10980 34660 11008 34700
rect 12544 34669 12572 34700
rect 16853 34697 16865 34731
rect 16899 34728 16911 34731
rect 19426 34728 19432 34740
rect 16899 34700 19432 34728
rect 16899 34697 16911 34700
rect 16853 34691 16911 34697
rect 19426 34688 19432 34700
rect 19484 34688 19490 34740
rect 20162 34688 20168 34740
rect 20220 34688 20226 34740
rect 20809 34731 20867 34737
rect 20809 34697 20821 34731
rect 20855 34728 20867 34731
rect 20990 34728 20996 34740
rect 20855 34700 20996 34728
rect 20855 34697 20867 34700
rect 20809 34691 20867 34697
rect 20990 34688 20996 34700
rect 21048 34688 21054 34740
rect 22830 34688 22836 34740
rect 22888 34688 22894 34740
rect 24029 34731 24087 34737
rect 24029 34728 24041 34731
rect 23584 34700 24041 34728
rect 12529 34663 12587 34669
rect 9456 34632 11008 34660
rect 11900 34632 12297 34660
rect 9456 34620 9462 34632
rect 11900 34604 11928 34632
rect 6825 34595 6883 34601
rect 6825 34561 6837 34595
rect 6871 34592 6883 34595
rect 7837 34595 7895 34601
rect 6871 34564 7788 34592
rect 6871 34561 6883 34564
rect 6825 34555 6883 34561
rect 4614 34484 4620 34536
rect 4672 34484 4678 34536
rect 6089 34527 6147 34533
rect 6089 34493 6101 34527
rect 6135 34524 6147 34527
rect 6840 34524 6868 34555
rect 7760 34536 7788 34564
rect 7837 34561 7849 34595
rect 7883 34561 7895 34595
rect 7837 34555 7895 34561
rect 9214 34552 9220 34604
rect 9272 34592 9278 34604
rect 10686 34592 10692 34604
rect 9272 34564 10692 34592
rect 9272 34552 9278 34564
rect 10686 34552 10692 34564
rect 10744 34592 10750 34604
rect 10870 34592 10876 34604
rect 10744 34564 10876 34592
rect 10744 34552 10750 34564
rect 10870 34552 10876 34564
rect 10928 34552 10934 34604
rect 11882 34552 11888 34604
rect 11940 34552 11946 34604
rect 12269 34601 12297 34632
rect 12529 34629 12541 34663
rect 12575 34660 12587 34663
rect 16114 34660 16120 34672
rect 12575 34632 16120 34660
rect 12575 34629 12587 34632
rect 12529 34623 12587 34629
rect 16114 34620 16120 34632
rect 16172 34620 16178 34672
rect 16758 34620 16764 34672
rect 16816 34660 16822 34672
rect 17218 34660 17224 34672
rect 16816 34632 17224 34660
rect 16816 34620 16822 34632
rect 17218 34620 17224 34632
rect 17276 34620 17282 34672
rect 17405 34663 17463 34669
rect 17405 34629 17417 34663
rect 17451 34660 17463 34663
rect 19794 34660 19800 34672
rect 17451 34632 19800 34660
rect 17451 34629 17463 34632
rect 17405 34623 17463 34629
rect 19794 34620 19800 34632
rect 19852 34620 19858 34672
rect 20073 34663 20131 34669
rect 20073 34629 20085 34663
rect 20119 34660 20131 34663
rect 20180 34660 20208 34688
rect 20119 34632 20208 34660
rect 20119 34629 20131 34632
rect 20073 34623 20131 34629
rect 20438 34620 20444 34672
rect 20496 34620 20502 34672
rect 20530 34620 20536 34672
rect 20588 34620 20594 34672
rect 20622 34620 20628 34672
rect 20680 34669 20686 34672
rect 20680 34663 20699 34669
rect 20687 34629 20699 34663
rect 20680 34623 20699 34629
rect 20680 34620 20686 34623
rect 21726 34620 21732 34672
rect 21784 34620 21790 34672
rect 22020 34632 22784 34660
rect 12161 34595 12219 34601
rect 12161 34561 12173 34595
rect 12207 34561 12219 34595
rect 12161 34555 12219 34561
rect 12254 34595 12312 34601
rect 12254 34561 12266 34595
rect 12300 34561 12312 34595
rect 12254 34555 12312 34561
rect 6135 34496 6868 34524
rect 6917 34527 6975 34533
rect 6135 34493 6147 34496
rect 6089 34487 6147 34493
rect 6917 34493 6929 34527
rect 6963 34493 6975 34527
rect 6917 34487 6975 34493
rect 6638 34416 6644 34468
rect 6696 34456 6702 34468
rect 6932 34456 6960 34487
rect 7742 34484 7748 34536
rect 7800 34484 7806 34536
rect 8110 34484 8116 34536
rect 8168 34484 8174 34536
rect 12176 34524 12204 34555
rect 12434 34552 12440 34604
rect 12492 34552 12498 34604
rect 12667 34595 12725 34601
rect 12667 34561 12679 34595
rect 12713 34592 12725 34595
rect 12894 34592 12900 34604
rect 12713 34564 12900 34592
rect 12713 34561 12725 34564
rect 12667 34555 12725 34561
rect 12894 34552 12900 34564
rect 12952 34592 12958 34604
rect 13170 34592 13176 34604
rect 12952 34564 13176 34592
rect 12952 34552 12958 34564
rect 13170 34552 13176 34564
rect 13228 34592 13234 34604
rect 15102 34592 15108 34604
rect 13228 34564 15108 34592
rect 13228 34552 13234 34564
rect 15102 34552 15108 34564
rect 15160 34552 15166 34604
rect 17129 34595 17187 34601
rect 17129 34592 17141 34595
rect 16776 34564 17141 34592
rect 16776 34524 16804 34564
rect 17129 34561 17141 34564
rect 17175 34561 17187 34595
rect 17129 34555 17187 34561
rect 17310 34552 17316 34604
rect 17368 34592 17374 34604
rect 17589 34595 17647 34601
rect 17589 34592 17601 34595
rect 17368 34564 17601 34592
rect 17368 34552 17374 34564
rect 17589 34561 17601 34564
rect 17635 34561 17647 34595
rect 17589 34555 17647 34561
rect 17678 34552 17684 34604
rect 17736 34552 17742 34604
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34592 17831 34595
rect 17862 34592 17868 34604
rect 17819 34564 17868 34592
rect 17819 34561 17831 34564
rect 17773 34555 17831 34561
rect 17862 34552 17868 34564
rect 17920 34552 17926 34604
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19889 34595 19947 34601
rect 19889 34592 19901 34595
rect 19484 34564 19901 34592
rect 19484 34552 19490 34564
rect 19889 34561 19901 34564
rect 19935 34561 19947 34595
rect 19889 34555 19947 34561
rect 20165 34595 20223 34601
rect 20165 34561 20177 34595
rect 20211 34561 20223 34595
rect 20165 34555 20223 34561
rect 12176 34496 12480 34524
rect 6696 34428 6960 34456
rect 12452 34456 12480 34496
rect 16408 34496 16804 34524
rect 12710 34456 12716 34468
rect 12452 34428 12716 34456
rect 6696 34416 6702 34428
rect 12710 34416 12716 34428
rect 12768 34416 12774 34468
rect 16408 34400 16436 34496
rect 16942 34484 16948 34536
rect 17000 34484 17006 34536
rect 17957 34527 18015 34533
rect 17957 34524 17969 34527
rect 17052 34496 17969 34524
rect 16666 34416 16672 34468
rect 16724 34456 16730 34468
rect 17052 34465 17080 34496
rect 17957 34493 17969 34496
rect 18003 34493 18015 34527
rect 17957 34487 18015 34493
rect 19978 34484 19984 34536
rect 20036 34484 20042 34536
rect 20180 34524 20208 34555
rect 20254 34552 20260 34604
rect 20312 34601 20318 34604
rect 20312 34595 20351 34601
rect 20339 34592 20351 34595
rect 20548 34592 20576 34620
rect 20339 34564 20576 34592
rect 20339 34561 20351 34564
rect 20312 34555 20351 34561
rect 20312 34552 20318 34555
rect 20806 34552 20812 34604
rect 20864 34552 20870 34604
rect 21744 34592 21772 34620
rect 22020 34601 22048 34632
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21744 34564 22017 34592
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22097 34595 22155 34601
rect 22097 34561 22109 34595
rect 22143 34592 22155 34595
rect 22186 34592 22192 34604
rect 22143 34564 22192 34592
rect 22143 34561 22155 34564
rect 22097 34555 22155 34561
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 22278 34552 22284 34604
rect 22336 34552 22342 34604
rect 22373 34595 22431 34601
rect 22373 34561 22385 34595
rect 22419 34561 22431 34595
rect 22373 34555 22431 34561
rect 20824 34524 20852 34552
rect 20180 34496 20852 34524
rect 21634 34484 21640 34536
rect 21692 34524 21698 34536
rect 22388 34524 22416 34555
rect 21692 34496 22416 34524
rect 21692 34484 21698 34496
rect 17037 34459 17095 34465
rect 16724 34428 16988 34456
rect 16724 34416 16730 34428
rect 6362 34348 6368 34400
rect 6420 34348 6426 34400
rect 12526 34348 12532 34400
rect 12584 34388 12590 34400
rect 12805 34391 12863 34397
rect 12805 34388 12817 34391
rect 12584 34360 12817 34388
rect 12584 34348 12590 34360
rect 12805 34357 12817 34360
rect 12851 34357 12863 34391
rect 12805 34351 12863 34357
rect 16390 34348 16396 34400
rect 16448 34348 16454 34400
rect 16850 34348 16856 34400
rect 16908 34348 16914 34400
rect 16960 34388 16988 34428
rect 17037 34425 17049 34459
rect 17083 34425 17095 34459
rect 22462 34456 22468 34468
rect 17037 34419 17095 34425
rect 19306 34428 22468 34456
rect 19306 34388 19334 34428
rect 22462 34416 22468 34428
rect 22520 34416 22526 34468
rect 22756 34456 22784 34632
rect 22848 34592 22876 34688
rect 23584 34660 23612 34700
rect 24029 34697 24041 34700
rect 24075 34697 24087 34731
rect 24029 34691 24087 34697
rect 24946 34688 24952 34740
rect 25004 34728 25010 34740
rect 25774 34728 25780 34740
rect 25004 34700 25780 34728
rect 25004 34688 25010 34700
rect 25774 34688 25780 34700
rect 25832 34688 25838 34740
rect 30929 34731 30987 34737
rect 25884 34700 29316 34728
rect 23124 34632 23612 34660
rect 23661 34663 23719 34669
rect 23124 34601 23152 34632
rect 23661 34629 23673 34663
rect 23707 34660 23719 34663
rect 24578 34660 24584 34672
rect 23707 34632 24584 34660
rect 23707 34629 23719 34632
rect 23661 34623 23719 34629
rect 24578 34620 24584 34632
rect 24636 34620 24642 34672
rect 25884 34660 25912 34700
rect 27246 34660 27252 34672
rect 25148 34632 25912 34660
rect 26988 34632 27252 34660
rect 23017 34595 23075 34601
rect 23017 34592 23029 34595
rect 22848 34564 23029 34592
rect 23017 34561 23029 34564
rect 23063 34561 23075 34595
rect 23017 34555 23075 34561
rect 23109 34595 23167 34601
rect 23109 34561 23121 34595
rect 23155 34561 23167 34595
rect 23109 34555 23167 34561
rect 23474 34552 23480 34604
rect 23532 34552 23538 34604
rect 23566 34552 23572 34604
rect 23624 34592 23630 34604
rect 23753 34595 23811 34601
rect 23753 34592 23765 34595
rect 23624 34564 23765 34592
rect 23624 34552 23630 34564
rect 23753 34561 23765 34564
rect 23799 34561 23811 34595
rect 23753 34555 23811 34561
rect 23845 34595 23903 34601
rect 23845 34561 23857 34595
rect 23891 34592 23903 34595
rect 25038 34592 25044 34604
rect 23891 34564 25044 34592
rect 23891 34561 23903 34564
rect 23845 34555 23903 34561
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25148 34601 25176 34632
rect 25133 34595 25191 34601
rect 25133 34561 25145 34595
rect 25179 34561 25191 34595
rect 25133 34555 25191 34561
rect 22833 34527 22891 34533
rect 22833 34493 22845 34527
rect 22879 34524 22891 34527
rect 22922 34524 22928 34536
rect 22879 34496 22928 34524
rect 22879 34493 22891 34496
rect 22833 34487 22891 34493
rect 22922 34484 22928 34496
rect 22980 34484 22986 34536
rect 23198 34484 23204 34536
rect 23256 34524 23262 34536
rect 23293 34527 23351 34533
rect 23293 34524 23305 34527
rect 23256 34496 23305 34524
rect 23256 34484 23262 34496
rect 23293 34493 23305 34496
rect 23339 34493 23351 34527
rect 23293 34487 23351 34493
rect 23382 34484 23388 34536
rect 23440 34484 23446 34536
rect 24486 34484 24492 34536
rect 24544 34524 24550 34536
rect 25148 34524 25176 34555
rect 25222 34552 25228 34604
rect 25280 34592 25286 34604
rect 25317 34595 25375 34601
rect 25317 34592 25329 34595
rect 25280 34564 25329 34592
rect 25280 34552 25286 34564
rect 25317 34561 25329 34564
rect 25363 34561 25375 34595
rect 25317 34555 25375 34561
rect 25409 34595 25467 34601
rect 25409 34561 25421 34595
rect 25455 34561 25467 34595
rect 25409 34555 25467 34561
rect 25501 34595 25559 34601
rect 25501 34561 25513 34595
rect 25547 34592 25559 34595
rect 25774 34592 25780 34604
rect 25547 34564 25780 34592
rect 25547 34561 25559 34564
rect 25501 34555 25559 34561
rect 24544 34496 25176 34524
rect 24544 34484 24550 34496
rect 25240 34456 25268 34552
rect 25424 34524 25452 34555
rect 25774 34552 25780 34564
rect 25832 34592 25838 34604
rect 25958 34592 25964 34604
rect 25832 34564 25964 34592
rect 25832 34552 25838 34564
rect 25958 34552 25964 34564
rect 26016 34552 26022 34604
rect 26510 34552 26516 34604
rect 26568 34552 26574 34604
rect 26988 34601 27016 34632
rect 27246 34620 27252 34632
rect 27304 34620 27310 34672
rect 27890 34620 27896 34672
rect 27948 34620 27954 34672
rect 26973 34595 27031 34601
rect 26973 34561 26985 34595
rect 27019 34561 27031 34595
rect 26973 34555 27031 34561
rect 29086 34552 29092 34604
rect 29144 34552 29150 34604
rect 29182 34595 29240 34601
rect 29182 34561 29194 34595
rect 29228 34561 29240 34595
rect 29288 34592 29316 34700
rect 30929 34697 30941 34731
rect 30975 34697 30987 34731
rect 30929 34691 30987 34697
rect 29362 34620 29368 34672
rect 29420 34660 29426 34672
rect 29914 34660 29920 34672
rect 29420 34632 29920 34660
rect 29420 34620 29426 34632
rect 29914 34620 29920 34632
rect 29972 34620 29978 34672
rect 29454 34592 29460 34604
rect 29288 34564 29460 34592
rect 29182 34555 29240 34561
rect 27249 34527 27307 34533
rect 27249 34524 27261 34527
rect 25424 34496 25544 34524
rect 25516 34468 25544 34496
rect 26344 34496 27261 34524
rect 22756 34428 25268 34456
rect 25498 34416 25504 34468
rect 25556 34416 25562 34468
rect 26344 34465 26372 34496
rect 27249 34493 27261 34496
rect 27295 34493 27307 34527
rect 27249 34487 27307 34493
rect 27890 34484 27896 34536
rect 27948 34524 27954 34536
rect 28534 34524 28540 34536
rect 27948 34496 28540 34524
rect 27948 34484 27954 34496
rect 28534 34484 28540 34496
rect 28592 34484 28598 34536
rect 29196 34524 29224 34555
rect 29454 34552 29460 34564
rect 29512 34552 29518 34604
rect 29595 34595 29653 34601
rect 29595 34561 29607 34595
rect 29641 34592 29653 34595
rect 30006 34592 30012 34604
rect 29641 34564 30012 34592
rect 29641 34561 29653 34564
rect 29595 34555 29653 34561
rect 30006 34552 30012 34564
rect 30064 34552 30070 34604
rect 30374 34552 30380 34604
rect 30432 34552 30438 34604
rect 30837 34595 30895 34601
rect 30837 34561 30849 34595
rect 30883 34592 30895 34595
rect 30944 34592 30972 34691
rect 30883 34564 30972 34592
rect 31297 34595 31355 34601
rect 30883 34561 30895 34564
rect 30837 34555 30895 34561
rect 31297 34561 31309 34595
rect 31343 34561 31355 34595
rect 31297 34555 31355 34561
rect 28966 34496 29224 34524
rect 30392 34524 30420 34552
rect 31110 34524 31116 34536
rect 30392 34496 31116 34524
rect 26329 34459 26387 34465
rect 26329 34425 26341 34459
rect 26375 34425 26387 34459
rect 26329 34419 26387 34425
rect 16960 34360 19334 34388
rect 20346 34348 20352 34400
rect 20404 34388 20410 34400
rect 20625 34391 20683 34397
rect 20625 34388 20637 34391
rect 20404 34360 20637 34388
rect 20404 34348 20410 34360
rect 20625 34357 20637 34360
rect 20671 34357 20683 34391
rect 20625 34351 20683 34357
rect 21818 34348 21824 34400
rect 21876 34348 21882 34400
rect 22738 34348 22744 34400
rect 22796 34388 22802 34400
rect 23198 34388 23204 34400
rect 22796 34360 23204 34388
rect 22796 34348 22802 34360
rect 23198 34348 23204 34360
rect 23256 34348 23262 34400
rect 25038 34348 25044 34400
rect 25096 34388 25102 34400
rect 25590 34388 25596 34400
rect 25096 34360 25596 34388
rect 25096 34348 25102 34360
rect 25590 34348 25596 34360
rect 25648 34348 25654 34400
rect 25682 34348 25688 34400
rect 25740 34348 25746 34400
rect 27246 34348 27252 34400
rect 27304 34388 27310 34400
rect 28721 34391 28779 34397
rect 28721 34388 28733 34391
rect 27304 34360 28733 34388
rect 27304 34348 27310 34360
rect 28721 34357 28733 34360
rect 28767 34388 28779 34391
rect 28966 34388 28994 34496
rect 31110 34484 31116 34496
rect 31168 34524 31174 34536
rect 31312 34524 31340 34555
rect 37550 34552 37556 34604
rect 37608 34552 37614 34604
rect 31168 34496 31340 34524
rect 31168 34484 31174 34496
rect 31386 34484 31392 34536
rect 31444 34484 31450 34536
rect 31481 34527 31539 34533
rect 31481 34493 31493 34527
rect 31527 34524 31539 34527
rect 33318 34524 33324 34536
rect 31527 34496 33324 34524
rect 31527 34493 31539 34496
rect 31481 34487 31539 34493
rect 29178 34416 29184 34468
rect 29236 34456 29242 34468
rect 31496 34456 31524 34487
rect 33318 34484 33324 34496
rect 33376 34484 33382 34536
rect 37829 34527 37887 34533
rect 37829 34493 37841 34527
rect 37875 34524 37887 34527
rect 37918 34524 37924 34536
rect 37875 34496 37924 34524
rect 37875 34493 37887 34496
rect 37829 34487 37887 34493
rect 37918 34484 37924 34496
rect 37976 34484 37982 34536
rect 29236 34428 31524 34456
rect 29236 34416 29242 34428
rect 28767 34360 28994 34388
rect 28767 34357 28779 34360
rect 28721 34351 28779 34357
rect 29730 34348 29736 34400
rect 29788 34348 29794 34400
rect 30650 34348 30656 34400
rect 30708 34348 30714 34400
rect 1104 34298 38272 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38272 34298
rect 1104 34224 38272 34246
rect 4614 34144 4620 34196
rect 4672 34184 4678 34196
rect 5353 34187 5411 34193
rect 5353 34184 5365 34187
rect 4672 34156 5365 34184
rect 4672 34144 4678 34156
rect 5353 34153 5365 34156
rect 5399 34153 5411 34187
rect 5353 34147 5411 34153
rect 8110 34144 8116 34196
rect 8168 34184 8174 34196
rect 8389 34187 8447 34193
rect 8389 34184 8401 34187
rect 8168 34156 8401 34184
rect 8168 34144 8174 34156
rect 8389 34153 8401 34156
rect 8435 34153 8447 34187
rect 8389 34147 8447 34153
rect 11974 34144 11980 34196
rect 12032 34184 12038 34196
rect 12802 34184 12808 34196
rect 12032 34156 12808 34184
rect 12032 34144 12038 34156
rect 12802 34144 12808 34156
rect 12860 34144 12866 34196
rect 14642 34144 14648 34196
rect 14700 34184 14706 34196
rect 14829 34187 14887 34193
rect 14829 34184 14841 34187
rect 14700 34156 14841 34184
rect 14700 34144 14706 34156
rect 14829 34153 14841 34156
rect 14875 34153 14887 34187
rect 14829 34147 14887 34153
rect 16117 34187 16175 34193
rect 16117 34153 16129 34187
rect 16163 34184 16175 34187
rect 16850 34184 16856 34196
rect 16163 34156 16856 34184
rect 16163 34153 16175 34156
rect 16117 34147 16175 34153
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 16942 34144 16948 34196
rect 17000 34184 17006 34196
rect 17405 34187 17463 34193
rect 17405 34184 17417 34187
rect 17000 34156 17417 34184
rect 17000 34144 17006 34156
rect 17405 34153 17417 34156
rect 17451 34153 17463 34187
rect 17405 34147 17463 34153
rect 20162 34144 20168 34196
rect 20220 34184 20226 34196
rect 22462 34184 22468 34196
rect 20220 34156 22468 34184
rect 20220 34144 20226 34156
rect 22462 34144 22468 34156
rect 22520 34144 22526 34196
rect 24949 34187 25007 34193
rect 24949 34153 24961 34187
rect 24995 34184 25007 34187
rect 25225 34187 25283 34193
rect 25225 34184 25237 34187
rect 24995 34156 25237 34184
rect 24995 34153 25007 34156
rect 24949 34147 25007 34153
rect 25225 34153 25237 34156
rect 25271 34153 25283 34187
rect 25225 34147 25283 34153
rect 26510 34144 26516 34196
rect 26568 34184 26574 34196
rect 26973 34187 27031 34193
rect 26973 34184 26985 34187
rect 26568 34156 26985 34184
rect 26568 34144 26574 34156
rect 26973 34153 26985 34156
rect 27019 34153 27031 34187
rect 26973 34147 27031 34153
rect 27430 34144 27436 34196
rect 27488 34184 27494 34196
rect 30374 34184 30380 34196
rect 27488 34156 30380 34184
rect 27488 34144 27494 34156
rect 30374 34144 30380 34156
rect 30432 34144 30438 34196
rect 30650 34144 30656 34196
rect 30708 34184 30714 34196
rect 30708 34156 31064 34184
rect 30708 34144 30714 34156
rect 12342 34076 12348 34128
rect 12400 34076 12406 34128
rect 14274 34076 14280 34128
rect 14332 34116 14338 34128
rect 14332 34088 30788 34116
rect 14332 34076 14338 34088
rect 7742 34008 7748 34060
rect 7800 34048 7806 34060
rect 7800 34020 9444 34048
rect 7800 34008 7806 34020
rect 4433 33983 4491 33989
rect 4433 33949 4445 33983
rect 4479 33980 4491 33983
rect 5442 33980 5448 33992
rect 4479 33952 5448 33980
rect 4479 33949 4491 33952
rect 4433 33943 4491 33949
rect 5442 33940 5448 33952
rect 5500 33940 5506 33992
rect 5537 33983 5595 33989
rect 5537 33949 5549 33983
rect 5583 33980 5595 33983
rect 6362 33980 6368 33992
rect 5583 33952 6368 33980
rect 5583 33949 5595 33952
rect 5537 33943 5595 33949
rect 6362 33940 6368 33952
rect 6420 33940 6426 33992
rect 7098 33940 7104 33992
rect 7156 33980 7162 33992
rect 8573 33983 8631 33989
rect 7156 33952 8248 33980
rect 7156 33940 7162 33952
rect 8220 33924 8248 33952
rect 8573 33949 8585 33983
rect 8619 33980 8631 33983
rect 8619 33952 9352 33980
rect 8619 33949 8631 33952
rect 8573 33943 8631 33949
rect 8202 33872 8208 33924
rect 8260 33872 8266 33924
rect 4522 33804 4528 33856
rect 4580 33804 4586 33856
rect 7190 33804 7196 33856
rect 7248 33804 7254 33856
rect 9324 33853 9352 33952
rect 9416 33912 9444 34020
rect 9950 34008 9956 34060
rect 10008 34008 10014 34060
rect 14461 34051 14519 34057
rect 14461 34017 14473 34051
rect 14507 34048 14519 34051
rect 18785 34051 18843 34057
rect 18785 34048 18797 34051
rect 14507 34020 18797 34048
rect 14507 34017 14519 34020
rect 14461 34011 14519 34017
rect 18785 34017 18797 34020
rect 18831 34017 18843 34051
rect 18785 34011 18843 34017
rect 19812 34020 20668 34048
rect 19812 33992 19840 34020
rect 9674 33940 9680 33992
rect 9732 33940 9738 33992
rect 10137 33983 10195 33989
rect 10137 33949 10149 33983
rect 10183 33980 10195 33983
rect 10226 33980 10232 33992
rect 10183 33952 10232 33980
rect 10183 33949 10195 33952
rect 10137 33943 10195 33949
rect 10226 33940 10232 33952
rect 10284 33940 10290 33992
rect 12335 33983 12393 33989
rect 12335 33949 12347 33983
rect 12381 33980 12393 33983
rect 12526 33980 12532 33992
rect 12381 33952 12532 33980
rect 12381 33949 12393 33952
rect 12335 33943 12393 33949
rect 12526 33940 12532 33952
rect 12584 33940 12590 33992
rect 12618 33940 12624 33992
rect 12676 33980 12682 33992
rect 12676 33952 13124 33980
rect 12676 33940 12682 33952
rect 9416 33884 12572 33912
rect 12544 33856 12572 33884
rect 13096 33856 13124 33952
rect 14734 33940 14740 33992
rect 14792 33940 14798 33992
rect 14918 33940 14924 33992
rect 14976 33940 14982 33992
rect 15197 33983 15255 33989
rect 15197 33949 15209 33983
rect 15243 33980 15255 33983
rect 15746 33980 15752 33992
rect 15243 33952 15752 33980
rect 15243 33949 15255 33952
rect 15197 33943 15255 33949
rect 15746 33940 15752 33952
rect 15804 33980 15810 33992
rect 16022 33980 16028 33992
rect 15804 33952 16028 33980
rect 15804 33940 15810 33952
rect 16022 33940 16028 33952
rect 16080 33940 16086 33992
rect 16114 33940 16120 33992
rect 16172 33980 16178 33992
rect 16393 33983 16451 33989
rect 16393 33980 16405 33983
rect 16172 33952 16405 33980
rect 16172 33940 16178 33952
rect 16393 33949 16405 33952
rect 16439 33949 16451 33983
rect 16393 33943 16451 33949
rect 16482 33940 16488 33992
rect 16540 33940 16546 33992
rect 16577 33983 16635 33989
rect 16577 33949 16589 33983
rect 16623 33949 16635 33983
rect 16577 33943 16635 33949
rect 15930 33872 15936 33924
rect 15988 33912 15994 33924
rect 16592 33912 16620 33943
rect 16666 33940 16672 33992
rect 16724 33940 16730 33992
rect 16761 33983 16819 33989
rect 16761 33949 16773 33983
rect 16807 33977 16819 33983
rect 16942 33980 16948 33992
rect 16868 33977 16948 33980
rect 16807 33952 16948 33977
rect 16807 33949 16896 33952
rect 16761 33943 16819 33949
rect 16942 33940 16948 33952
rect 17000 33980 17006 33992
rect 17221 33983 17279 33989
rect 17221 33980 17233 33983
rect 17000 33952 17233 33980
rect 17000 33940 17006 33952
rect 17221 33949 17233 33952
rect 17267 33949 17279 33983
rect 17221 33943 17279 33949
rect 17681 33983 17739 33989
rect 17681 33949 17693 33983
rect 17727 33949 17739 33983
rect 17681 33943 17739 33949
rect 15988 33884 16620 33912
rect 16684 33912 16712 33940
rect 16853 33915 16911 33921
rect 16853 33912 16865 33915
rect 16684 33884 16865 33912
rect 15988 33872 15994 33884
rect 9309 33847 9367 33853
rect 9309 33813 9321 33847
rect 9355 33813 9367 33847
rect 9309 33807 9367 33813
rect 9766 33804 9772 33856
rect 9824 33804 9830 33856
rect 9858 33804 9864 33856
rect 9916 33844 9922 33856
rect 10229 33847 10287 33853
rect 10229 33844 10241 33847
rect 9916 33816 10241 33844
rect 9916 33804 9922 33816
rect 10229 33813 10241 33816
rect 10275 33813 10287 33847
rect 10229 33807 10287 33813
rect 12526 33804 12532 33856
rect 12584 33804 12590 33856
rect 13078 33804 13084 33856
rect 13136 33804 13142 33856
rect 15105 33847 15163 33853
rect 15105 33813 15117 33847
rect 15151 33844 15163 33847
rect 16684 33844 16712 33884
rect 16853 33881 16865 33884
rect 16899 33881 16911 33915
rect 16853 33875 16911 33881
rect 17037 33915 17095 33921
rect 17037 33881 17049 33915
rect 17083 33912 17095 33915
rect 17083 33884 17264 33912
rect 17083 33881 17095 33884
rect 17037 33875 17095 33881
rect 17236 33856 17264 33884
rect 15151 33816 16712 33844
rect 15151 33813 15163 33816
rect 15105 33807 15163 33813
rect 17126 33804 17132 33856
rect 17184 33804 17190 33856
rect 17218 33804 17224 33856
rect 17276 33804 17282 33856
rect 17310 33804 17316 33856
rect 17368 33844 17374 33856
rect 17696 33844 17724 33943
rect 18046 33940 18052 33992
rect 18104 33940 18110 33992
rect 18509 33983 18567 33989
rect 18509 33980 18521 33983
rect 18248 33952 18521 33980
rect 17862 33872 17868 33924
rect 17920 33872 17926 33924
rect 17954 33872 17960 33924
rect 18012 33872 18018 33924
rect 18248 33853 18276 33952
rect 18509 33949 18521 33952
rect 18555 33949 18567 33983
rect 18509 33943 18567 33949
rect 18601 33983 18659 33989
rect 18601 33949 18613 33983
rect 18647 33949 18659 33983
rect 18601 33943 18659 33949
rect 17368 33816 17724 33844
rect 18233 33847 18291 33853
rect 17368 33804 17374 33816
rect 18233 33813 18245 33847
rect 18279 33813 18291 33847
rect 18233 33807 18291 33813
rect 18506 33804 18512 33856
rect 18564 33804 18570 33856
rect 18616 33844 18644 33943
rect 19794 33940 19800 33992
rect 19852 33940 19858 33992
rect 20349 33983 20407 33989
rect 20349 33949 20361 33983
rect 20395 33980 20407 33983
rect 20438 33980 20444 33992
rect 20395 33952 20444 33980
rect 20395 33949 20407 33952
rect 20349 33943 20407 33949
rect 20438 33940 20444 33952
rect 20496 33940 20502 33992
rect 20640 33989 20668 34020
rect 21174 34008 21180 34060
rect 21232 34048 21238 34060
rect 24302 34048 24308 34060
rect 21232 34020 24308 34048
rect 21232 34008 21238 34020
rect 24302 34008 24308 34020
rect 24360 34008 24366 34060
rect 24578 34008 24584 34060
rect 24636 34008 24642 34060
rect 27246 34048 27252 34060
rect 25332 34020 27252 34048
rect 20625 33983 20683 33989
rect 20625 33949 20637 33983
rect 20671 33949 20683 33983
rect 20625 33943 20683 33949
rect 20717 33983 20775 33989
rect 20717 33949 20729 33983
rect 20763 33980 20775 33983
rect 21726 33980 21732 33992
rect 20763 33952 21732 33980
rect 20763 33949 20775 33952
rect 20717 33943 20775 33949
rect 19334 33872 19340 33924
rect 19392 33912 19398 33924
rect 20530 33912 20536 33924
rect 19392 33884 20536 33912
rect 19392 33872 19398 33884
rect 20530 33872 20536 33884
rect 20588 33872 20594 33924
rect 20640 33912 20668 33943
rect 21726 33940 21732 33952
rect 21784 33980 21790 33992
rect 22370 33980 22376 33992
rect 21784 33952 22376 33980
rect 21784 33940 21790 33952
rect 22370 33940 22376 33952
rect 22428 33940 22434 33992
rect 25332 33980 25360 34020
rect 24504 33952 25360 33980
rect 24504 33912 24532 33952
rect 25406 33940 25412 33992
rect 25464 33940 25470 33992
rect 25516 33989 25544 34020
rect 27246 34008 27252 34020
rect 27304 34048 27310 34060
rect 27433 34051 27491 34057
rect 27433 34048 27445 34051
rect 27304 34020 27445 34048
rect 27304 34008 27310 34020
rect 27433 34017 27445 34020
rect 27479 34017 27491 34051
rect 27433 34011 27491 34017
rect 27522 34008 27528 34060
rect 27580 34048 27586 34060
rect 28626 34048 28632 34060
rect 27580 34020 28632 34048
rect 27580 34008 27586 34020
rect 28626 34008 28632 34020
rect 28684 34008 28690 34060
rect 29546 34008 29552 34060
rect 29604 34048 29610 34060
rect 29604 34020 30328 34048
rect 29604 34008 29610 34020
rect 25501 33983 25559 33989
rect 25501 33949 25513 33983
rect 25547 33949 25559 33983
rect 25501 33943 25559 33949
rect 25682 33940 25688 33992
rect 25740 33940 25746 33992
rect 25777 33983 25835 33989
rect 25777 33949 25789 33983
rect 25823 33980 25835 33983
rect 26050 33980 26056 33992
rect 25823 33952 26056 33980
rect 25823 33949 25835 33952
rect 25777 33943 25835 33949
rect 26050 33940 26056 33952
rect 26108 33940 26114 33992
rect 28261 33983 28319 33989
rect 28261 33949 28273 33983
rect 28307 33949 28319 33983
rect 28261 33943 28319 33949
rect 20640 33884 24532 33912
rect 24670 33872 24676 33924
rect 24728 33912 24734 33924
rect 27706 33912 27712 33924
rect 24728 33884 27712 33912
rect 24728 33872 24734 33884
rect 27706 33872 27712 33884
rect 27764 33912 27770 33924
rect 28276 33912 28304 33943
rect 29730 33940 29736 33992
rect 29788 33980 29794 33992
rect 30300 33989 30328 34020
rect 30009 33983 30067 33989
rect 30009 33980 30021 33983
rect 29788 33952 30021 33980
rect 29788 33940 29794 33952
rect 30009 33949 30021 33952
rect 30055 33949 30067 33983
rect 30009 33943 30067 33949
rect 30285 33983 30343 33989
rect 30285 33949 30297 33983
rect 30331 33980 30343 33983
rect 30374 33980 30380 33992
rect 30331 33952 30380 33980
rect 30331 33949 30343 33952
rect 30285 33943 30343 33949
rect 30374 33940 30380 33952
rect 30432 33940 30438 33992
rect 30760 33989 30788 34088
rect 31036 34048 31064 34156
rect 31386 34144 31392 34196
rect 31444 34184 31450 34196
rect 32769 34187 32827 34193
rect 32769 34184 32781 34187
rect 31444 34156 32781 34184
rect 31444 34144 31450 34156
rect 32769 34153 32781 34156
rect 32815 34153 32827 34187
rect 32769 34147 32827 34153
rect 32858 34144 32864 34196
rect 32916 34184 32922 34196
rect 33873 34187 33931 34193
rect 33873 34184 33885 34187
rect 32916 34156 33885 34184
rect 32916 34144 32922 34156
rect 33873 34153 33885 34156
rect 33919 34153 33931 34187
rect 33873 34147 33931 34153
rect 32953 34119 33011 34125
rect 32953 34085 32965 34119
rect 32999 34116 33011 34119
rect 32999 34088 34284 34116
rect 32999 34085 33011 34088
rect 32953 34079 33011 34085
rect 31297 34051 31355 34057
rect 31297 34048 31309 34051
rect 31036 34020 31309 34048
rect 31297 34017 31309 34020
rect 31343 34017 31355 34051
rect 31297 34011 31355 34017
rect 33597 34051 33655 34057
rect 33597 34017 33609 34051
rect 33643 34048 33655 34051
rect 33686 34048 33692 34060
rect 33643 34020 33692 34048
rect 33643 34017 33655 34020
rect 33597 34011 33655 34017
rect 33686 34008 33692 34020
rect 33744 34008 33750 34060
rect 30745 33983 30803 33989
rect 30745 33949 30757 33983
rect 30791 33949 30803 33983
rect 30745 33943 30803 33949
rect 30837 33983 30895 33989
rect 30837 33949 30849 33983
rect 30883 33980 30895 33983
rect 31021 33983 31079 33989
rect 31021 33980 31033 33983
rect 30883 33952 31033 33980
rect 30883 33949 30895 33952
rect 30837 33943 30895 33949
rect 31021 33949 31033 33952
rect 31067 33949 31079 33983
rect 32674 33980 32680 33992
rect 32430 33952 32680 33980
rect 31021 33943 31079 33949
rect 32674 33940 32680 33952
rect 32732 33940 32738 33992
rect 32766 33940 32772 33992
rect 32824 33980 32830 33992
rect 34256 33989 34284 34088
rect 33781 33983 33839 33989
rect 33781 33980 33793 33983
rect 32824 33952 33793 33980
rect 32824 33940 32830 33952
rect 33781 33949 33793 33952
rect 33827 33949 33839 33983
rect 33781 33943 33839 33949
rect 34241 33983 34299 33989
rect 34241 33949 34253 33983
rect 34287 33949 34299 33983
rect 34241 33943 34299 33949
rect 27764 33884 28304 33912
rect 29825 33915 29883 33921
rect 27764 33872 27770 33884
rect 29825 33881 29837 33915
rect 29871 33912 29883 33915
rect 30466 33912 30472 33924
rect 29871 33884 30472 33912
rect 29871 33881 29883 33884
rect 29825 33875 29883 33881
rect 30466 33872 30472 33884
rect 30524 33872 30530 33924
rect 32692 33912 32720 33940
rect 33134 33912 33140 33924
rect 32692 33884 33140 33912
rect 33134 33872 33140 33884
rect 33192 33872 33198 33924
rect 33413 33915 33471 33921
rect 33413 33912 33425 33915
rect 33244 33884 33425 33912
rect 33244 33856 33272 33884
rect 33413 33881 33425 33884
rect 33459 33881 33471 33915
rect 33796 33912 33824 33943
rect 34606 33912 34612 33924
rect 33796 33884 34612 33912
rect 33413 33875 33471 33881
rect 34606 33872 34612 33884
rect 34664 33872 34670 33924
rect 20901 33847 20959 33853
rect 20901 33844 20913 33847
rect 18616 33816 20913 33844
rect 20901 33813 20913 33816
rect 20947 33813 20959 33847
rect 20901 33807 20959 33813
rect 21542 33804 21548 33856
rect 21600 33844 21606 33856
rect 21910 33844 21916 33856
rect 21600 33816 21916 33844
rect 21600 33804 21606 33816
rect 21910 33804 21916 33816
rect 21968 33844 21974 33856
rect 22646 33844 22652 33856
rect 21968 33816 22652 33844
rect 21968 33804 21974 33816
rect 22646 33804 22652 33816
rect 22704 33804 22710 33856
rect 24949 33847 25007 33853
rect 24949 33813 24961 33847
rect 24995 33844 25007 33847
rect 25038 33844 25044 33856
rect 24995 33816 25044 33844
rect 24995 33813 25007 33816
rect 24949 33807 25007 33813
rect 25038 33804 25044 33816
rect 25096 33804 25102 33856
rect 25130 33804 25136 33856
rect 25188 33804 25194 33856
rect 26510 33804 26516 33856
rect 26568 33844 26574 33856
rect 27341 33847 27399 33853
rect 27341 33844 27353 33847
rect 26568 33816 27353 33844
rect 26568 33804 26574 33816
rect 27341 33813 27353 33816
rect 27387 33844 27399 33847
rect 27430 33844 27436 33856
rect 27387 33816 27436 33844
rect 27387 33813 27399 33816
rect 27341 33807 27399 33813
rect 27430 33804 27436 33816
rect 27488 33804 27494 33856
rect 28350 33804 28356 33856
rect 28408 33804 28414 33856
rect 28442 33804 28448 33856
rect 28500 33844 28506 33856
rect 30193 33847 30251 33853
rect 30193 33844 30205 33847
rect 28500 33816 30205 33844
rect 28500 33804 28506 33816
rect 30193 33813 30205 33816
rect 30239 33844 30251 33847
rect 31386 33844 31392 33856
rect 30239 33816 31392 33844
rect 30239 33813 30251 33816
rect 30193 33807 30251 33813
rect 31386 33804 31392 33816
rect 31444 33804 31450 33856
rect 33226 33804 33232 33856
rect 33284 33804 33290 33856
rect 33318 33804 33324 33856
rect 33376 33804 33382 33856
rect 34057 33847 34115 33853
rect 34057 33813 34069 33847
rect 34103 33844 34115 33847
rect 34146 33844 34152 33856
rect 34103 33816 34152 33844
rect 34103 33813 34115 33816
rect 34057 33807 34115 33813
rect 34146 33804 34152 33816
rect 34204 33804 34210 33856
rect 1104 33754 38272 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38272 33754
rect 1104 33680 38272 33702
rect 4522 33600 4528 33652
rect 4580 33600 4586 33652
rect 7190 33600 7196 33652
rect 7248 33600 7254 33652
rect 9858 33600 9864 33652
rect 9916 33600 9922 33652
rect 14737 33643 14795 33649
rect 14737 33609 14749 33643
rect 14783 33640 14795 33643
rect 14918 33640 14924 33652
rect 14783 33612 14924 33640
rect 14783 33609 14795 33612
rect 14737 33603 14795 33609
rect 14918 33600 14924 33612
rect 14976 33600 14982 33652
rect 17037 33643 17095 33649
rect 17037 33609 17049 33643
rect 17083 33609 17095 33643
rect 17037 33603 17095 33609
rect 4540 33572 4568 33600
rect 6822 33572 6828 33584
rect 4356 33544 4568 33572
rect 5842 33544 6828 33572
rect 4356 33513 4384 33544
rect 6822 33532 6828 33544
rect 6880 33532 6886 33584
rect 7208 33572 7236 33600
rect 9214 33572 9220 33584
rect 7024 33544 7236 33572
rect 8510 33544 9220 33572
rect 7024 33513 7052 33544
rect 9214 33532 9220 33544
rect 9272 33532 9278 33584
rect 9876 33572 9904 33600
rect 9508 33544 9904 33572
rect 9508 33513 9536 33544
rect 10318 33532 10324 33584
rect 10376 33532 10382 33584
rect 12526 33532 12532 33584
rect 12584 33572 12590 33584
rect 14090 33572 14096 33584
rect 12584 33544 14096 33572
rect 12584 33532 12590 33544
rect 14090 33532 14096 33544
rect 14148 33572 14154 33584
rect 14185 33575 14243 33581
rect 14185 33572 14197 33575
rect 14148 33544 14197 33572
rect 14148 33532 14154 33544
rect 14185 33541 14197 33544
rect 14231 33541 14243 33575
rect 14185 33535 14243 33541
rect 14458 33532 14464 33584
rect 14516 33572 14522 33584
rect 14516 33544 14688 33572
rect 14516 33532 14522 33544
rect 14660 33516 14688 33544
rect 16114 33532 16120 33584
rect 16172 33572 16178 33584
rect 16669 33575 16727 33581
rect 16669 33572 16681 33575
rect 16172 33544 16681 33572
rect 16172 33532 16178 33544
rect 4341 33507 4399 33513
rect 4341 33473 4353 33507
rect 4387 33473 4399 33507
rect 4341 33467 4399 33473
rect 7009 33507 7067 33513
rect 7009 33473 7021 33507
rect 7055 33473 7067 33507
rect 7009 33467 7067 33473
rect 9493 33507 9551 33513
rect 9493 33473 9505 33507
rect 9539 33473 9551 33507
rect 9493 33467 9551 33473
rect 14366 33464 14372 33516
rect 14424 33464 14430 33516
rect 14550 33464 14556 33516
rect 14608 33464 14614 33516
rect 14642 33464 14648 33516
rect 14700 33464 14706 33516
rect 4614 33396 4620 33448
rect 4672 33396 4678 33448
rect 7282 33396 7288 33448
rect 7340 33396 7346 33448
rect 9766 33396 9772 33448
rect 9824 33396 9830 33448
rect 11241 33439 11299 33445
rect 11241 33405 11253 33439
rect 11287 33436 11299 33439
rect 11609 33439 11667 33445
rect 11609 33436 11621 33439
rect 11287 33408 11621 33436
rect 11287 33405 11299 33408
rect 11241 33399 11299 33405
rect 11609 33405 11621 33408
rect 11655 33436 11667 33439
rect 16592 33436 16620 33544
rect 16669 33541 16681 33544
rect 16715 33541 16727 33575
rect 16669 33535 16727 33541
rect 16899 33541 16957 33547
rect 16899 33538 16911 33541
rect 16884 33516 16911 33538
rect 16850 33464 16856 33516
rect 16908 33507 16911 33516
rect 16945 33507 16957 33541
rect 16908 33501 16957 33507
rect 17052 33504 17080 33603
rect 18506 33600 18512 33652
rect 18564 33600 18570 33652
rect 23937 33643 23995 33649
rect 23937 33640 23949 33643
rect 18708 33612 23949 33640
rect 17402 33532 17408 33584
rect 17460 33532 17466 33584
rect 17494 33532 17500 33584
rect 17552 33532 17558 33584
rect 18524 33572 18552 33600
rect 18340 33544 18552 33572
rect 17129 33507 17187 33513
rect 17129 33504 17141 33507
rect 16908 33464 16914 33501
rect 17052 33476 17141 33504
rect 17129 33473 17141 33476
rect 17175 33473 17187 33507
rect 17129 33467 17187 33473
rect 17222 33507 17280 33513
rect 17222 33473 17234 33507
rect 17268 33504 17280 33507
rect 17635 33507 17693 33513
rect 17268 33476 17448 33504
rect 17268 33473 17280 33476
rect 17222 33467 17280 33473
rect 17420 33448 17448 33476
rect 17635 33473 17647 33507
rect 17681 33504 17693 33507
rect 17770 33504 17776 33516
rect 17681 33476 17776 33504
rect 17681 33473 17693 33476
rect 17635 33467 17693 33473
rect 17770 33464 17776 33476
rect 17828 33464 17834 33516
rect 18340 33513 18368 33544
rect 18141 33507 18199 33513
rect 18141 33473 18153 33507
rect 18187 33473 18199 33507
rect 18141 33467 18199 33473
rect 18325 33507 18383 33513
rect 18325 33473 18337 33507
rect 18371 33473 18383 33507
rect 18325 33467 18383 33473
rect 18509 33507 18567 33513
rect 18509 33473 18521 33507
rect 18555 33504 18567 33507
rect 18708 33504 18736 33612
rect 23937 33609 23949 33612
rect 23983 33609 23995 33643
rect 23937 33603 23995 33609
rect 24302 33600 24308 33652
rect 24360 33640 24366 33652
rect 24489 33643 24547 33649
rect 24489 33640 24501 33643
rect 24360 33612 24501 33640
rect 24360 33600 24366 33612
rect 24489 33609 24501 33612
rect 24535 33609 24547 33643
rect 24489 33603 24547 33609
rect 28350 33600 28356 33652
rect 28408 33600 28414 33652
rect 28828 33612 31754 33640
rect 19981 33575 20039 33581
rect 19981 33572 19993 33575
rect 19444 33544 19993 33572
rect 18555 33476 18736 33504
rect 18555 33473 18567 33476
rect 18509 33467 18567 33473
rect 17310 33436 17316 33448
rect 11655 33408 14044 33436
rect 16592 33408 17316 33436
rect 11655 33405 11667 33408
rect 11609 33399 11667 33405
rect 9490 33328 9496 33380
rect 9548 33328 9554 33380
rect 12526 33368 12532 33380
rect 10980 33340 12532 33368
rect 6089 33303 6147 33309
rect 6089 33269 6101 33303
rect 6135 33300 6147 33303
rect 6178 33300 6184 33312
rect 6135 33272 6184 33300
rect 6135 33269 6147 33272
rect 6089 33263 6147 33269
rect 6178 33260 6184 33272
rect 6236 33260 6242 33312
rect 8754 33260 8760 33312
rect 8812 33260 8818 33312
rect 9508 33300 9536 33328
rect 10980 33300 11008 33340
rect 12526 33328 12532 33340
rect 12584 33328 12590 33380
rect 14016 33368 14044 33408
rect 17310 33396 17316 33408
rect 17368 33396 17374 33448
rect 17402 33396 17408 33448
rect 17460 33396 17466 33448
rect 17954 33368 17960 33380
rect 14016 33340 17960 33368
rect 17954 33328 17960 33340
rect 18012 33328 18018 33380
rect 18156 33368 18184 33467
rect 18782 33464 18788 33516
rect 18840 33464 18846 33516
rect 19038 33507 19096 33513
rect 19038 33473 19050 33507
rect 19084 33504 19096 33507
rect 19444 33504 19472 33544
rect 19981 33541 19993 33544
rect 20027 33541 20039 33575
rect 19981 33535 20039 33541
rect 21082 33532 21088 33584
rect 21140 33572 21146 33584
rect 22002 33572 22008 33584
rect 21140 33544 22008 33572
rect 21140 33532 21146 33544
rect 22002 33532 22008 33544
rect 22060 33532 22066 33584
rect 22094 33532 22100 33584
rect 22152 33532 22158 33584
rect 22189 33575 22247 33581
rect 22189 33541 22201 33575
rect 22235 33572 22247 33575
rect 22738 33572 22744 33584
rect 22235 33544 22744 33572
rect 22235 33541 22247 33544
rect 22189 33535 22247 33541
rect 22738 33532 22744 33544
rect 22796 33572 22802 33584
rect 23290 33572 23296 33584
rect 22796 33544 23296 33572
rect 22796 33532 22802 33544
rect 23290 33532 23296 33544
rect 23348 33532 23354 33584
rect 24946 33572 24952 33584
rect 24412 33544 24952 33572
rect 19705 33507 19763 33513
rect 19705 33504 19717 33507
rect 19084 33476 19472 33504
rect 19536 33476 19717 33504
rect 19084 33473 19096 33476
rect 19038 33467 19096 33473
rect 18874 33396 18880 33448
rect 18932 33436 18938 33448
rect 19426 33436 19432 33448
rect 18932 33408 19432 33436
rect 18932 33396 18938 33408
rect 19426 33396 19432 33408
rect 19484 33436 19490 33448
rect 19536 33436 19564 33476
rect 19705 33473 19717 33476
rect 19751 33473 19763 33507
rect 19705 33467 19763 33473
rect 19886 33464 19892 33516
rect 19944 33504 19950 33516
rect 20530 33504 20536 33516
rect 19944 33476 20536 33504
rect 19944 33464 19950 33476
rect 20530 33464 20536 33476
rect 20588 33504 20594 33516
rect 21450 33504 21456 33516
rect 20588 33476 21456 33504
rect 20588 33464 20594 33476
rect 21450 33464 21456 33476
rect 21508 33464 21514 33516
rect 23750 33464 23756 33516
rect 23808 33504 23814 33516
rect 24412 33513 24440 33544
rect 24946 33532 24952 33544
rect 25004 33572 25010 33584
rect 28368 33572 28396 33600
rect 25004 33544 25728 33572
rect 25004 33532 25010 33544
rect 25700 33516 25728 33544
rect 28184 33544 28396 33572
rect 23845 33507 23903 33513
rect 23845 33504 23857 33507
rect 23808 33476 23857 33504
rect 23808 33464 23814 33476
rect 23845 33473 23857 33476
rect 23891 33473 23903 33507
rect 23845 33467 23903 33473
rect 24029 33507 24087 33513
rect 24029 33473 24041 33507
rect 24075 33473 24087 33507
rect 24029 33467 24087 33473
rect 24397 33507 24455 33513
rect 24397 33473 24409 33507
rect 24443 33473 24455 33507
rect 24397 33467 24455 33473
rect 24581 33507 24639 33513
rect 24581 33473 24593 33507
rect 24627 33473 24639 33507
rect 24581 33467 24639 33473
rect 19484 33408 19564 33436
rect 19484 33396 19490 33408
rect 19610 33396 19616 33448
rect 19668 33396 19674 33448
rect 19981 33439 20039 33445
rect 19981 33405 19993 33439
rect 20027 33436 20039 33439
rect 20027 33408 21956 33436
rect 20027 33405 20039 33408
rect 19981 33399 20039 33405
rect 19996 33368 20024 33399
rect 18156 33340 20024 33368
rect 21726 33328 21732 33380
rect 21784 33368 21790 33380
rect 21821 33371 21879 33377
rect 21821 33368 21833 33371
rect 21784 33340 21833 33368
rect 21784 33328 21790 33340
rect 21821 33337 21833 33340
rect 21867 33337 21879 33371
rect 21928 33368 21956 33408
rect 23382 33396 23388 33448
rect 23440 33396 23446 33448
rect 24044 33436 24072 33467
rect 24596 33436 24624 33467
rect 25682 33464 25688 33516
rect 25740 33464 25746 33516
rect 28184 33513 28212 33544
rect 28534 33532 28540 33584
rect 28592 33572 28598 33584
rect 28828 33572 28856 33612
rect 31726 33584 31754 33612
rect 33318 33600 33324 33652
rect 33376 33640 33382 33652
rect 34609 33643 34667 33649
rect 34609 33640 34621 33643
rect 33376 33612 34621 33640
rect 33376 33600 33382 33612
rect 34609 33609 34621 33612
rect 34655 33609 34667 33643
rect 34609 33603 34667 33609
rect 37369 33643 37427 33649
rect 37369 33609 37381 33643
rect 37415 33640 37427 33643
rect 37550 33640 37556 33652
rect 37415 33612 37556 33640
rect 37415 33609 37427 33612
rect 37369 33603 37427 33609
rect 37550 33600 37556 33612
rect 37608 33600 37614 33652
rect 28592 33544 28934 33572
rect 28592 33532 28598 33544
rect 31662 33532 31668 33584
rect 31720 33572 31754 33584
rect 33594 33572 33600 33584
rect 31720 33544 33600 33572
rect 31720 33532 31726 33544
rect 33594 33532 33600 33544
rect 33652 33532 33658 33584
rect 28169 33507 28227 33513
rect 28169 33473 28181 33507
rect 28215 33473 28227 33507
rect 28169 33467 28227 33473
rect 32858 33464 32864 33516
rect 32916 33464 32922 33516
rect 34146 33464 34152 33516
rect 34204 33464 34210 33516
rect 37550 33464 37556 33516
rect 37608 33464 37614 33516
rect 26234 33436 26240 33448
rect 24044 33408 26240 33436
rect 26234 33396 26240 33408
rect 26292 33396 26298 33448
rect 28442 33396 28448 33448
rect 28500 33396 28506 33448
rect 33137 33439 33195 33445
rect 33137 33405 33149 33439
rect 33183 33436 33195 33439
rect 34164 33436 34192 33464
rect 33183 33408 34192 33436
rect 33183 33405 33195 33408
rect 33137 33399 33195 33405
rect 23400 33368 23428 33396
rect 21928 33340 23428 33368
rect 21821 33331 21879 33337
rect 9508 33272 11008 33300
rect 11054 33260 11060 33312
rect 11112 33300 11118 33312
rect 12161 33303 12219 33309
rect 12161 33300 12173 33303
rect 11112 33272 12173 33300
rect 11112 33260 11118 33272
rect 12161 33269 12173 33272
rect 12207 33269 12219 33303
rect 12161 33263 12219 33269
rect 15930 33260 15936 33312
rect 15988 33300 15994 33312
rect 16853 33303 16911 33309
rect 16853 33300 16865 33303
rect 15988 33272 16865 33300
rect 15988 33260 15994 33272
rect 16853 33269 16865 33272
rect 16899 33269 16911 33303
rect 16853 33263 16911 33269
rect 17773 33303 17831 33309
rect 17773 33269 17785 33303
rect 17819 33300 17831 33303
rect 18322 33300 18328 33312
rect 17819 33272 18328 33300
rect 17819 33269 17831 33272
rect 17773 33263 17831 33269
rect 18322 33260 18328 33272
rect 18380 33260 18386 33312
rect 19797 33303 19855 33309
rect 19797 33269 19809 33303
rect 19843 33300 19855 33303
rect 21358 33300 21364 33312
rect 19843 33272 21364 33300
rect 19843 33269 19855 33272
rect 19797 33263 19855 33269
rect 21358 33260 21364 33272
rect 21416 33260 21422 33312
rect 22373 33303 22431 33309
rect 22373 33269 22385 33303
rect 22419 33300 22431 33303
rect 22830 33300 22836 33312
rect 22419 33272 22836 33300
rect 22419 33269 22431 33272
rect 22373 33263 22431 33269
rect 22830 33260 22836 33272
rect 22888 33260 22894 33312
rect 29730 33260 29736 33312
rect 29788 33300 29794 33312
rect 29917 33303 29975 33309
rect 29917 33300 29929 33303
rect 29788 33272 29929 33300
rect 29788 33260 29794 33272
rect 29917 33269 29929 33272
rect 29963 33269 29975 33303
rect 29917 33263 29975 33269
rect 30190 33260 30196 33312
rect 30248 33300 30254 33312
rect 33318 33300 33324 33312
rect 30248 33272 33324 33300
rect 30248 33260 30254 33272
rect 33318 33260 33324 33272
rect 33376 33260 33382 33312
rect 1104 33210 38272 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38272 33210
rect 1104 33136 38272 33158
rect 4614 33056 4620 33108
rect 4672 33096 4678 33108
rect 5169 33099 5227 33105
rect 5169 33096 5181 33099
rect 4672 33068 5181 33096
rect 4672 33056 4678 33068
rect 5169 33065 5181 33068
rect 5215 33065 5227 33099
rect 5169 33059 5227 33065
rect 7282 33056 7288 33108
rect 7340 33096 7346 33108
rect 7561 33099 7619 33105
rect 7561 33096 7573 33099
rect 7340 33068 7573 33096
rect 7340 33056 7346 33068
rect 7561 33065 7573 33068
rect 7607 33065 7619 33099
rect 7561 33059 7619 33065
rect 8110 33056 8116 33108
rect 8168 33096 8174 33108
rect 8168 33068 8432 33096
rect 8168 33056 8174 33068
rect 5721 33031 5779 33037
rect 5721 32997 5733 33031
rect 5767 32997 5779 33031
rect 5721 32991 5779 32997
rect 5353 32895 5411 32901
rect 5353 32861 5365 32895
rect 5399 32892 5411 32895
rect 5736 32892 5764 32991
rect 6365 32963 6423 32969
rect 6365 32929 6377 32963
rect 6411 32960 6423 32963
rect 6638 32960 6644 32972
rect 6411 32932 6644 32960
rect 6411 32929 6423 32932
rect 6365 32923 6423 32929
rect 6638 32920 6644 32932
rect 6696 32920 6702 32972
rect 8110 32960 8116 32972
rect 7484 32932 8116 32960
rect 5399 32864 5764 32892
rect 6089 32895 6147 32901
rect 5399 32861 5411 32864
rect 5353 32855 5411 32861
rect 6089 32861 6101 32895
rect 6135 32892 6147 32895
rect 7484 32892 7512 32932
rect 8110 32920 8116 32932
rect 8168 32960 8174 32972
rect 8297 32963 8355 32969
rect 8297 32960 8309 32963
rect 8168 32932 8309 32960
rect 8168 32920 8174 32932
rect 8297 32929 8309 32932
rect 8343 32929 8355 32963
rect 8404 32960 8432 33068
rect 9766 33056 9772 33108
rect 9824 33056 9830 33108
rect 10042 33096 10048 33108
rect 9876 33068 10048 33096
rect 9876 33028 9904 33068
rect 10042 33056 10048 33068
rect 10100 33096 10106 33108
rect 10502 33096 10508 33108
rect 10100 33068 10508 33096
rect 10100 33056 10106 33068
rect 10502 33056 10508 33068
rect 10560 33056 10566 33108
rect 16945 33099 17003 33105
rect 16945 33065 16957 33099
rect 16991 33096 17003 33099
rect 17126 33096 17132 33108
rect 16991 33068 17132 33096
rect 16991 33065 17003 33068
rect 16945 33059 17003 33065
rect 17126 33056 17132 33068
rect 17184 33096 17190 33108
rect 17402 33096 17408 33108
rect 17184 33068 17408 33096
rect 17184 33056 17190 33068
rect 17402 33056 17408 33068
rect 17460 33096 17466 33108
rect 17678 33096 17684 33108
rect 17460 33068 17684 33096
rect 17460 33056 17466 33068
rect 17678 33056 17684 33068
rect 17736 33056 17742 33108
rect 18322 33056 18328 33108
rect 18380 33056 18386 33108
rect 20162 33056 20168 33108
rect 20220 33096 20226 33108
rect 20220 33068 20760 33096
rect 20220 33056 20226 33068
rect 20438 33028 20444 33040
rect 9646 33000 9904 33028
rect 12361 33000 19012 33028
rect 8481 32963 8539 32969
rect 8481 32960 8493 32963
rect 8404 32932 8493 32960
rect 8297 32923 8355 32929
rect 8481 32929 8493 32932
rect 8527 32960 8539 32963
rect 9646 32960 9674 33000
rect 10229 32963 10287 32969
rect 8527 32932 9674 32960
rect 9784 32932 10180 32960
rect 8527 32929 8539 32932
rect 8481 32923 8539 32929
rect 6135 32864 7512 32892
rect 7745 32895 7803 32901
rect 6135 32861 6147 32864
rect 6089 32855 6147 32861
rect 7745 32861 7757 32895
rect 7791 32892 7803 32895
rect 8205 32895 8263 32901
rect 7791 32864 7880 32892
rect 7791 32861 7803 32864
rect 7745 32855 7803 32861
rect 6178 32716 6184 32768
rect 6236 32716 6242 32768
rect 7852 32765 7880 32864
rect 8205 32861 8217 32895
rect 8251 32892 8263 32895
rect 8754 32892 8760 32904
rect 8251 32864 8760 32892
rect 8251 32861 8263 32864
rect 8205 32855 8263 32861
rect 8754 32852 8760 32864
rect 8812 32852 8818 32904
rect 8938 32852 8944 32904
rect 8996 32892 9002 32904
rect 9490 32892 9496 32904
rect 8996 32864 9496 32892
rect 8996 32852 9002 32864
rect 9490 32852 9496 32864
rect 9548 32892 9554 32904
rect 9784 32892 9812 32932
rect 9548 32864 9812 32892
rect 9548 32852 9554 32864
rect 9950 32852 9956 32904
rect 10008 32852 10014 32904
rect 10042 32852 10048 32904
rect 10100 32852 10106 32904
rect 10152 32892 10180 32932
rect 10229 32929 10241 32963
rect 10275 32960 10287 32963
rect 10505 32963 10563 32969
rect 10505 32960 10517 32963
rect 10275 32932 10517 32960
rect 10275 32929 10287 32932
rect 10229 32923 10287 32929
rect 10505 32929 10517 32932
rect 10551 32929 10563 32963
rect 10505 32923 10563 32929
rect 12361 32901 12389 33000
rect 18984 32972 19012 33000
rect 19306 33000 20444 33028
rect 12636 32932 14504 32960
rect 12636 32901 12664 32932
rect 10321 32895 10379 32901
rect 10321 32892 10333 32895
rect 10152 32864 10333 32892
rect 10321 32861 10333 32864
rect 10367 32861 10379 32895
rect 10321 32855 10379 32861
rect 10413 32895 10471 32901
rect 10413 32861 10425 32895
rect 10459 32861 10471 32895
rect 12361 32895 12423 32901
rect 12361 32892 12377 32895
rect 10413 32855 10471 32861
rect 10612 32864 12377 32892
rect 8846 32784 8852 32836
rect 8904 32824 8910 32836
rect 10428 32824 10456 32855
rect 8904 32796 10456 32824
rect 8904 32784 8910 32796
rect 7837 32759 7895 32765
rect 7837 32725 7849 32759
rect 7883 32725 7895 32759
rect 7837 32719 7895 32725
rect 9398 32716 9404 32768
rect 9456 32756 9462 32768
rect 10612 32756 10640 32864
rect 12365 32861 12377 32864
rect 12411 32861 12423 32895
rect 12621 32895 12679 32901
rect 12621 32892 12633 32895
rect 12365 32855 12423 32861
rect 12452 32864 12633 32892
rect 10686 32784 10692 32836
rect 10744 32824 10750 32836
rect 12452 32824 12480 32864
rect 12621 32861 12633 32864
rect 12667 32861 12679 32895
rect 12621 32855 12679 32861
rect 12713 32895 12771 32901
rect 12713 32861 12725 32895
rect 12759 32892 12771 32895
rect 13078 32892 13084 32904
rect 12759 32864 13084 32892
rect 12759 32861 12771 32864
rect 12713 32855 12771 32861
rect 13078 32852 13084 32864
rect 13136 32852 13142 32904
rect 14476 32836 14504 32932
rect 15654 32920 15660 32972
rect 15712 32960 15718 32972
rect 16298 32960 16304 32972
rect 15712 32932 16304 32960
rect 15712 32920 15718 32932
rect 16298 32920 16304 32932
rect 16356 32960 16362 32972
rect 17862 32960 17868 32972
rect 16356 32932 17868 32960
rect 16356 32920 16362 32932
rect 17862 32920 17868 32932
rect 17920 32920 17926 32972
rect 18874 32960 18880 32972
rect 18156 32932 18880 32960
rect 17954 32852 17960 32904
rect 18012 32892 18018 32904
rect 18156 32901 18184 32932
rect 18874 32920 18880 32932
rect 18932 32920 18938 32972
rect 18966 32920 18972 32972
rect 19024 32920 19030 32972
rect 18141 32895 18199 32901
rect 18141 32892 18153 32895
rect 18012 32864 18153 32892
rect 18012 32852 18018 32864
rect 18141 32861 18153 32864
rect 18187 32861 18199 32895
rect 18141 32855 18199 32861
rect 18230 32852 18236 32904
rect 18288 32892 18294 32904
rect 18417 32895 18475 32901
rect 18417 32892 18429 32895
rect 18288 32864 18429 32892
rect 18288 32852 18294 32864
rect 18417 32861 18429 32864
rect 18463 32892 18475 32895
rect 19306 32892 19334 33000
rect 20438 32988 20444 33000
rect 20496 32988 20502 33040
rect 20732 32960 20760 33068
rect 22278 33056 22284 33108
rect 22336 33096 22342 33108
rect 23842 33096 23848 33108
rect 22336 33068 23848 33096
rect 22336 33056 22342 33068
rect 23842 33056 23848 33068
rect 23900 33056 23906 33108
rect 27893 33099 27951 33105
rect 27893 33065 27905 33099
rect 27939 33096 27951 33099
rect 28442 33096 28448 33108
rect 27939 33068 28448 33096
rect 27939 33065 27951 33068
rect 27893 33059 27951 33065
rect 28442 33056 28448 33068
rect 28500 33056 28506 33108
rect 30285 33099 30343 33105
rect 30285 33065 30297 33099
rect 30331 33096 30343 33099
rect 37550 33096 37556 33108
rect 30331 33068 37556 33096
rect 30331 33065 30343 33068
rect 30285 33059 30343 33065
rect 37550 33056 37556 33068
rect 37608 33056 37614 33108
rect 21910 32988 21916 33040
rect 21968 33028 21974 33040
rect 22738 33028 22744 33040
rect 21968 33000 22744 33028
rect 21968 32988 21974 33000
rect 22738 32988 22744 33000
rect 22796 32988 22802 33040
rect 28169 33031 28227 33037
rect 28169 33028 28181 33031
rect 27816 33000 28181 33028
rect 21269 32963 21327 32969
rect 21269 32960 21281 32963
rect 20732 32932 21281 32960
rect 21269 32929 21281 32932
rect 21315 32960 21327 32963
rect 21315 32932 21772 32960
rect 21315 32929 21327 32932
rect 21269 32923 21327 32929
rect 18463 32864 19334 32892
rect 18463 32861 18475 32864
rect 18417 32855 18475 32861
rect 20622 32852 20628 32904
rect 20680 32892 20686 32904
rect 20990 32892 20996 32904
rect 20680 32864 20996 32892
rect 20680 32852 20686 32864
rect 20990 32852 20996 32864
rect 21048 32892 21054 32904
rect 21637 32895 21695 32901
rect 21637 32892 21649 32895
rect 21048 32864 21649 32892
rect 21048 32852 21054 32864
rect 21637 32861 21649 32864
rect 21683 32861 21695 32895
rect 21637 32855 21695 32861
rect 10744 32796 12480 32824
rect 12529 32827 12587 32833
rect 10744 32784 10750 32796
rect 12529 32793 12541 32827
rect 12575 32824 12587 32827
rect 13446 32824 13452 32836
rect 12575 32796 13452 32824
rect 12575 32793 12587 32796
rect 12529 32787 12587 32793
rect 12728 32768 12756 32796
rect 13446 32784 13452 32796
rect 13504 32784 13510 32836
rect 14458 32784 14464 32836
rect 14516 32784 14522 32836
rect 16298 32784 16304 32836
rect 16356 32824 16362 32836
rect 16761 32827 16819 32833
rect 16761 32824 16773 32827
rect 16356 32796 16773 32824
rect 16356 32784 16362 32796
rect 16761 32793 16773 32796
rect 16807 32824 16819 32827
rect 17218 32824 17224 32836
rect 16807 32796 17224 32824
rect 16807 32793 16819 32796
rect 16761 32787 16819 32793
rect 17218 32784 17224 32796
rect 17276 32784 17282 32836
rect 18049 32827 18107 32833
rect 18049 32793 18061 32827
rect 18095 32793 18107 32827
rect 18049 32787 18107 32793
rect 18509 32827 18567 32833
rect 18509 32793 18521 32827
rect 18555 32824 18567 32827
rect 18690 32824 18696 32836
rect 18555 32796 18696 32824
rect 18555 32793 18567 32796
rect 18509 32787 18567 32793
rect 9456 32728 10640 32756
rect 9456 32716 9462 32728
rect 12710 32716 12716 32768
rect 12768 32716 12774 32768
rect 12802 32716 12808 32768
rect 12860 32756 12866 32768
rect 12897 32759 12955 32765
rect 12897 32756 12909 32759
rect 12860 32728 12909 32756
rect 12860 32716 12866 32728
rect 12897 32725 12909 32728
rect 12943 32725 12955 32759
rect 12897 32719 12955 32725
rect 16942 32716 16948 32768
rect 17000 32716 17006 32768
rect 17129 32759 17187 32765
rect 17129 32725 17141 32759
rect 17175 32756 17187 32759
rect 17586 32756 17592 32768
rect 17175 32728 17592 32756
rect 17175 32725 17187 32728
rect 17129 32719 17187 32725
rect 17586 32716 17592 32728
rect 17644 32716 17650 32768
rect 17954 32716 17960 32768
rect 18012 32756 18018 32768
rect 18064 32756 18092 32787
rect 18690 32784 18696 32796
rect 18748 32784 18754 32836
rect 19426 32784 19432 32836
rect 19484 32784 19490 32836
rect 21545 32827 21603 32833
rect 21545 32824 21557 32827
rect 20088 32796 21220 32824
rect 20088 32768 20116 32796
rect 21192 32768 21220 32796
rect 21376 32796 21557 32824
rect 19886 32756 19892 32768
rect 18012 32728 19892 32756
rect 18012 32716 18018 32728
rect 19886 32716 19892 32728
rect 19944 32716 19950 32768
rect 20070 32716 20076 32768
rect 20128 32716 20134 32768
rect 20622 32716 20628 32768
rect 20680 32756 20686 32768
rect 20717 32759 20775 32765
rect 20717 32756 20729 32759
rect 20680 32728 20729 32756
rect 20680 32716 20686 32728
rect 20717 32725 20729 32728
rect 20763 32725 20775 32759
rect 20717 32719 20775 32725
rect 21174 32716 21180 32768
rect 21232 32756 21238 32768
rect 21376 32756 21404 32796
rect 21545 32793 21557 32796
rect 21591 32793 21603 32827
rect 21744 32824 21772 32932
rect 22020 32932 22325 32960
rect 22020 32904 22048 32932
rect 22002 32852 22008 32904
rect 22060 32852 22066 32904
rect 22186 32852 22192 32904
rect 22244 32852 22250 32904
rect 22297 32901 22325 32932
rect 22572 32932 26280 32960
rect 22282 32895 22340 32901
rect 22282 32861 22294 32895
rect 22328 32892 22340 32895
rect 22572 32892 22600 32932
rect 22328 32864 22600 32892
rect 22328 32861 22340 32864
rect 22282 32855 22340 32861
rect 22646 32852 22652 32904
rect 22704 32901 22710 32904
rect 22704 32892 22712 32901
rect 22704 32864 22749 32892
rect 22704 32855 22712 32864
rect 22704 32852 22710 32855
rect 22830 32852 22836 32904
rect 22888 32892 22894 32904
rect 22925 32895 22983 32901
rect 22925 32892 22937 32895
rect 22888 32864 22937 32892
rect 22888 32852 22894 32864
rect 22925 32861 22937 32864
rect 22971 32861 22983 32895
rect 22925 32855 22983 32861
rect 23014 32852 23020 32904
rect 23072 32892 23078 32904
rect 23390 32895 23448 32901
rect 23072 32864 23117 32892
rect 23072 32852 23078 32864
rect 23390 32861 23402 32895
rect 23436 32861 23448 32895
rect 23390 32855 23448 32861
rect 21744 32796 22324 32824
rect 21545 32787 21603 32793
rect 21232 32728 21404 32756
rect 21232 32716 21238 32728
rect 21450 32716 21456 32768
rect 21508 32716 21514 32768
rect 21818 32716 21824 32768
rect 21876 32716 21882 32768
rect 22296 32756 22324 32796
rect 22370 32784 22376 32836
rect 22428 32824 22434 32836
rect 22465 32827 22523 32833
rect 22465 32824 22477 32827
rect 22428 32796 22477 32824
rect 22428 32784 22434 32796
rect 22465 32793 22477 32796
rect 22511 32793 22523 32827
rect 22465 32787 22523 32793
rect 22557 32827 22615 32833
rect 22557 32793 22569 32827
rect 22603 32793 22615 32827
rect 22557 32787 22615 32793
rect 23201 32827 23259 32833
rect 23201 32793 23213 32827
rect 23247 32793 23259 32827
rect 23201 32787 23259 32793
rect 22572 32756 22600 32787
rect 22296 32728 22600 32756
rect 22738 32716 22744 32768
rect 22796 32756 22802 32768
rect 22833 32759 22891 32765
rect 22833 32756 22845 32759
rect 22796 32728 22845 32756
rect 22796 32716 22802 32728
rect 22833 32725 22845 32728
rect 22879 32725 22891 32759
rect 22833 32719 22891 32725
rect 23106 32716 23112 32768
rect 23164 32756 23170 32768
rect 23216 32756 23244 32787
rect 23290 32784 23296 32836
rect 23348 32784 23354 32836
rect 23405 32824 23433 32855
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 25406 32892 25412 32904
rect 23900 32864 25412 32892
rect 23900 32852 23906 32864
rect 25406 32852 25412 32864
rect 25464 32892 25470 32904
rect 25774 32892 25780 32904
rect 25464 32864 25780 32892
rect 25464 32852 25470 32864
rect 25774 32852 25780 32864
rect 25832 32852 25838 32904
rect 25884 32901 25912 32932
rect 25869 32895 25927 32901
rect 25869 32861 25881 32895
rect 25915 32861 25927 32895
rect 25869 32855 25927 32861
rect 26050 32852 26056 32904
rect 26108 32852 26114 32904
rect 26142 32852 26148 32904
rect 26200 32852 26206 32904
rect 24026 32824 24032 32836
rect 23405 32796 24032 32824
rect 24026 32784 24032 32796
rect 24084 32824 24090 32836
rect 24302 32824 24308 32836
rect 24084 32796 24308 32824
rect 24084 32784 24090 32796
rect 24302 32784 24308 32796
rect 24360 32784 24366 32836
rect 26252 32824 26280 32932
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 26605 32895 26663 32901
rect 26605 32892 26617 32895
rect 26384 32864 26617 32892
rect 26384 32852 26390 32864
rect 26605 32861 26617 32864
rect 26651 32861 26663 32895
rect 26605 32855 26663 32861
rect 27062 32852 27068 32904
rect 27120 32852 27126 32904
rect 27816 32892 27844 33000
rect 28169 32997 28181 33000
rect 28215 32997 28227 33031
rect 31478 33028 31484 33040
rect 28169 32991 28227 32997
rect 28552 33000 31484 33028
rect 28552 32901 28580 33000
rect 31478 32988 31484 33000
rect 31536 32988 31542 33040
rect 32861 33031 32919 33037
rect 32861 32997 32873 33031
rect 32907 33028 32919 33031
rect 32907 33000 33916 33028
rect 32907 32997 32919 33000
rect 32861 32991 32919 32997
rect 28626 32920 28632 32972
rect 28684 32960 28690 32972
rect 28721 32963 28779 32969
rect 28721 32960 28733 32963
rect 28684 32932 28733 32960
rect 28684 32920 28690 32932
rect 28721 32929 28733 32932
rect 28767 32960 28779 32963
rect 28902 32960 28908 32972
rect 28767 32932 28908 32960
rect 28767 32929 28779 32932
rect 28721 32923 28779 32929
rect 28902 32920 28908 32932
rect 28960 32920 28966 32972
rect 28077 32895 28135 32901
rect 28077 32892 28089 32895
rect 27816 32864 28089 32892
rect 28077 32861 28089 32864
rect 28123 32861 28135 32895
rect 28537 32895 28595 32901
rect 28537 32892 28549 32895
rect 28077 32855 28135 32861
rect 28368 32864 28549 32892
rect 26252 32796 27292 32824
rect 23164 32728 23244 32756
rect 23164 32716 23170 32728
rect 23474 32716 23480 32768
rect 23532 32756 23538 32768
rect 23569 32759 23627 32765
rect 23569 32756 23581 32759
rect 23532 32728 23581 32756
rect 23532 32716 23538 32728
rect 23569 32725 23581 32728
rect 23615 32725 23627 32759
rect 23569 32719 23627 32725
rect 25590 32716 25596 32768
rect 25648 32716 25654 32768
rect 26418 32716 26424 32768
rect 26476 32716 26482 32768
rect 27154 32716 27160 32768
rect 27212 32716 27218 32768
rect 27264 32756 27292 32796
rect 27890 32784 27896 32836
rect 27948 32824 27954 32836
rect 28368 32824 28396 32864
rect 28537 32861 28549 32864
rect 28583 32861 28595 32895
rect 28537 32855 28595 32861
rect 28994 32852 29000 32904
rect 29052 32892 29058 32904
rect 29917 32895 29975 32901
rect 29917 32892 29929 32895
rect 29052 32864 29929 32892
rect 29052 32852 29058 32864
rect 29917 32861 29929 32864
rect 29963 32861 29975 32895
rect 29917 32855 29975 32861
rect 30101 32895 30159 32901
rect 30101 32861 30113 32895
rect 30147 32861 30159 32895
rect 31496 32892 31524 32988
rect 33410 32920 33416 32972
rect 33468 32920 33474 32972
rect 33226 32892 33232 32904
rect 31496 32864 33232 32892
rect 30101 32855 30159 32861
rect 27948 32796 28396 32824
rect 27948 32784 27954 32796
rect 28442 32784 28448 32836
rect 28500 32824 28506 32836
rect 30116 32824 30144 32855
rect 33226 32852 33232 32864
rect 33284 32852 33290 32904
rect 33888 32901 33916 33000
rect 33873 32895 33931 32901
rect 33873 32861 33885 32895
rect 33919 32861 33931 32895
rect 33873 32855 33931 32861
rect 34701 32895 34759 32901
rect 34701 32861 34713 32895
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 28500 32796 30144 32824
rect 28500 32784 28506 32796
rect 30742 32784 30748 32836
rect 30800 32824 30806 32836
rect 33321 32827 33379 32833
rect 33321 32824 33333 32827
rect 30800 32796 33333 32824
rect 30800 32784 30806 32796
rect 33321 32793 33333 32796
rect 33367 32824 33379 32827
rect 33962 32824 33968 32836
rect 33367 32796 33968 32824
rect 33367 32793 33379 32796
rect 33321 32787 33379 32793
rect 33962 32784 33968 32796
rect 34020 32784 34026 32836
rect 34606 32784 34612 32836
rect 34664 32824 34670 32836
rect 34716 32824 34744 32855
rect 34790 32852 34796 32904
rect 34848 32892 34854 32904
rect 34977 32895 35035 32901
rect 34977 32892 34989 32895
rect 34848 32864 34989 32892
rect 34848 32852 34854 32864
rect 34977 32861 34989 32864
rect 35023 32861 35035 32895
rect 34977 32855 35035 32861
rect 34664 32796 34744 32824
rect 34664 32784 34670 32796
rect 28629 32759 28687 32765
rect 28629 32756 28641 32759
rect 27264 32728 28641 32756
rect 28629 32725 28641 32728
rect 28675 32756 28687 32759
rect 29730 32756 29736 32768
rect 28675 32728 29736 32756
rect 28675 32725 28687 32728
rect 28629 32719 28687 32725
rect 29730 32716 29736 32728
rect 29788 32716 29794 32768
rect 33686 32716 33692 32768
rect 33744 32716 33750 32768
rect 34790 32716 34796 32768
rect 34848 32716 34854 32768
rect 35066 32716 35072 32768
rect 35124 32716 35130 32768
rect 1104 32666 38272 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38272 32666
rect 1104 32592 38272 32614
rect 8754 32512 8760 32564
rect 8812 32552 8818 32564
rect 12342 32552 12348 32564
rect 8812 32524 12348 32552
rect 8812 32512 8818 32524
rect 12342 32512 12348 32524
rect 12400 32552 12406 32564
rect 12400 32524 20944 32552
rect 12400 32512 12406 32524
rect 6178 32444 6184 32496
rect 6236 32484 6242 32496
rect 6236 32456 7880 32484
rect 6236 32444 6242 32456
rect 5350 32376 5356 32428
rect 5408 32416 5414 32428
rect 7745 32419 7803 32425
rect 7745 32416 7757 32419
rect 5408 32388 7757 32416
rect 5408 32376 5414 32388
rect 7745 32385 7757 32388
rect 7791 32385 7803 32419
rect 7852 32416 7880 32456
rect 10042 32444 10048 32496
rect 10100 32484 10106 32496
rect 11054 32484 11060 32496
rect 10100 32456 11060 32484
rect 10100 32444 10106 32456
rect 11054 32444 11060 32456
rect 11112 32444 11118 32496
rect 11900 32456 12664 32484
rect 10686 32416 10692 32428
rect 7852 32388 10692 32416
rect 7745 32379 7803 32385
rect 10686 32376 10692 32388
rect 10744 32376 10750 32428
rect 10873 32419 10931 32425
rect 10873 32385 10885 32419
rect 10919 32416 10931 32419
rect 11514 32416 11520 32428
rect 10919 32388 11520 32416
rect 10919 32385 10931 32388
rect 10873 32379 10931 32385
rect 11514 32376 11520 32388
rect 11572 32376 11578 32428
rect 6730 32308 6736 32360
rect 6788 32348 6794 32360
rect 11900 32348 11928 32456
rect 11974 32376 11980 32428
rect 12032 32416 12038 32428
rect 12253 32419 12311 32425
rect 12253 32416 12265 32419
rect 12032 32388 12265 32416
rect 12032 32376 12038 32388
rect 12253 32385 12265 32388
rect 12299 32385 12311 32419
rect 12253 32379 12311 32385
rect 12342 32376 12348 32428
rect 12400 32416 12406 32428
rect 12636 32425 12664 32456
rect 18248 32456 18553 32484
rect 18248 32428 18276 32456
rect 12529 32419 12587 32425
rect 12400 32388 12445 32416
rect 12400 32376 12406 32388
rect 12529 32385 12541 32419
rect 12575 32385 12587 32419
rect 12529 32379 12587 32385
rect 12621 32419 12679 32425
rect 12621 32385 12633 32419
rect 12667 32385 12679 32419
rect 12621 32379 12679 32385
rect 12759 32419 12817 32425
rect 12759 32385 12771 32419
rect 12805 32416 12817 32419
rect 12894 32416 12900 32428
rect 12805 32388 12900 32416
rect 12805 32385 12817 32388
rect 12759 32379 12817 32385
rect 6788 32320 11928 32348
rect 6788 32308 6794 32320
rect 12434 32308 12440 32360
rect 12492 32348 12498 32360
rect 12544 32348 12572 32379
rect 12492 32320 12572 32348
rect 12636 32348 12664 32379
rect 12894 32376 12900 32388
rect 12952 32376 12958 32428
rect 12989 32419 13047 32425
rect 12989 32385 13001 32419
rect 13035 32416 13047 32419
rect 15194 32416 15200 32428
rect 13035 32388 15200 32416
rect 13035 32385 13047 32388
rect 12989 32379 13047 32385
rect 15194 32376 15200 32388
rect 15252 32376 15258 32428
rect 18230 32376 18236 32428
rect 18288 32376 18294 32428
rect 18322 32376 18328 32428
rect 18380 32416 18386 32428
rect 18525 32425 18553 32456
rect 20714 32444 20720 32496
rect 20772 32444 20778 32496
rect 20916 32493 20944 32524
rect 21818 32512 21824 32564
rect 21876 32512 21882 32564
rect 22186 32512 22192 32564
rect 22244 32552 22250 32564
rect 22370 32552 22376 32564
rect 22244 32524 22376 32552
rect 22244 32512 22250 32524
rect 22370 32512 22376 32524
rect 22428 32512 22434 32564
rect 22646 32512 22652 32564
rect 22704 32552 22710 32564
rect 22925 32555 22983 32561
rect 22925 32552 22937 32555
rect 22704 32524 22937 32552
rect 22704 32512 22710 32524
rect 22925 32521 22937 32524
rect 22971 32521 22983 32555
rect 22925 32515 22983 32521
rect 23014 32512 23020 32564
rect 23072 32552 23078 32564
rect 23072 32524 23704 32552
rect 23072 32512 23078 32524
rect 20901 32487 20959 32493
rect 20901 32453 20913 32487
rect 20947 32484 20959 32487
rect 20947 32456 21128 32484
rect 20947 32453 20959 32456
rect 20901 32447 20959 32453
rect 18417 32419 18475 32425
rect 18417 32416 18429 32419
rect 18380 32388 18429 32416
rect 18380 32376 18386 32388
rect 18417 32385 18429 32388
rect 18463 32385 18475 32419
rect 18417 32379 18475 32385
rect 18509 32419 18567 32425
rect 18509 32385 18521 32419
rect 18555 32385 18567 32419
rect 18509 32379 18567 32385
rect 18690 32376 18696 32428
rect 18748 32376 18754 32428
rect 18785 32419 18843 32425
rect 18785 32385 18797 32419
rect 18831 32416 18843 32419
rect 18874 32416 18880 32428
rect 18831 32388 18880 32416
rect 18831 32385 18843 32388
rect 18785 32379 18843 32385
rect 18874 32376 18880 32388
rect 18932 32376 18938 32428
rect 19150 32376 19156 32428
rect 19208 32416 19214 32428
rect 19245 32419 19303 32425
rect 19245 32416 19257 32419
rect 19208 32388 19257 32416
rect 19208 32376 19214 32388
rect 19245 32385 19257 32388
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 19518 32376 19524 32428
rect 19576 32416 19582 32428
rect 20070 32416 20076 32428
rect 19576 32388 20076 32416
rect 19576 32376 19582 32388
rect 20070 32376 20076 32388
rect 20128 32376 20134 32428
rect 20625 32419 20683 32425
rect 20625 32385 20637 32419
rect 20671 32385 20683 32419
rect 20732 32416 20760 32444
rect 20809 32419 20867 32425
rect 20809 32416 20821 32419
rect 20732 32388 20821 32416
rect 20625 32379 20683 32385
rect 20809 32385 20821 32388
rect 20855 32385 20867 32419
rect 20809 32379 20867 32385
rect 20993 32419 21051 32425
rect 20993 32385 21005 32419
rect 21039 32385 21051 32419
rect 20993 32379 21051 32385
rect 12636 32320 14412 32348
rect 12492 32308 12498 32320
rect 12544 32280 12572 32320
rect 12618 32280 12624 32292
rect 12544 32252 12624 32280
rect 12618 32240 12624 32252
rect 12676 32240 12682 32292
rect 14384 32280 14412 32320
rect 14458 32308 14464 32360
rect 14516 32348 14522 32360
rect 20162 32348 20168 32360
rect 14516 32320 20168 32348
rect 14516 32308 14522 32320
rect 20162 32308 20168 32320
rect 20220 32348 20226 32360
rect 20640 32348 20668 32379
rect 21008 32348 21036 32379
rect 20220 32320 20668 32348
rect 20916 32320 21036 32348
rect 21100 32348 21128 32456
rect 21836 32425 21864 32512
rect 22301 32456 22968 32484
rect 22002 32425 22008 32428
rect 21821 32419 21879 32425
rect 21821 32385 21833 32419
rect 21867 32385 21879 32419
rect 21821 32379 21879 32385
rect 21969 32419 22008 32425
rect 21969 32385 21981 32419
rect 21969 32379 22008 32385
rect 22002 32376 22008 32379
rect 22060 32376 22066 32428
rect 22094 32376 22100 32428
rect 22152 32376 22158 32428
rect 22301 32425 22329 32456
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32385 22247 32419
rect 22189 32379 22247 32385
rect 22286 32419 22344 32425
rect 22286 32385 22298 32419
rect 22332 32385 22344 32419
rect 22286 32379 22344 32385
rect 21726 32348 21732 32360
rect 21100 32320 21732 32348
rect 20220 32308 20226 32320
rect 20714 32280 20720 32292
rect 14384 32252 20720 32280
rect 20714 32240 20720 32252
rect 20772 32240 20778 32292
rect 20916 32280 20944 32320
rect 21726 32308 21732 32320
rect 21784 32348 21790 32360
rect 22204 32348 22232 32379
rect 22664 32360 22692 32456
rect 22940 32428 22968 32456
rect 23106 32444 23112 32496
rect 23164 32484 23170 32496
rect 23382 32484 23388 32496
rect 23164 32456 23388 32484
rect 23164 32444 23170 32456
rect 23382 32444 23388 32456
rect 23440 32444 23446 32496
rect 23474 32444 23480 32496
rect 23532 32444 23538 32496
rect 23676 32484 23704 32524
rect 25590 32512 25596 32564
rect 25648 32512 25654 32564
rect 26053 32555 26111 32561
rect 26053 32521 26065 32555
rect 26099 32552 26111 32555
rect 26326 32552 26332 32564
rect 26099 32524 26332 32552
rect 26099 32521 26111 32524
rect 26053 32515 26111 32521
rect 26326 32512 26332 32524
rect 26384 32512 26390 32564
rect 26418 32512 26424 32564
rect 26476 32552 26482 32564
rect 26476 32524 26924 32552
rect 26476 32512 26482 32524
rect 25608 32484 25636 32512
rect 23676 32456 24624 32484
rect 25608 32456 25820 32484
rect 22738 32376 22744 32428
rect 22796 32376 22802 32428
rect 22922 32376 22928 32428
rect 22980 32376 22986 32428
rect 23201 32419 23259 32425
rect 23201 32385 23213 32419
rect 23247 32416 23336 32419
rect 23492 32416 23520 32444
rect 23676 32425 23704 32456
rect 24596 32428 24624 32456
rect 23247 32391 23520 32416
rect 23247 32385 23259 32391
rect 23308 32388 23520 32391
rect 23569 32419 23627 32425
rect 23201 32379 23259 32385
rect 23569 32385 23581 32419
rect 23615 32385 23627 32419
rect 23569 32379 23627 32385
rect 23661 32419 23719 32425
rect 23661 32385 23673 32419
rect 23707 32385 23719 32419
rect 23661 32379 23719 32385
rect 21784 32320 22232 32348
rect 21784 32308 21790 32320
rect 22646 32308 22652 32360
rect 22704 32308 22710 32360
rect 22278 32280 22284 32292
rect 20916 32252 22284 32280
rect 7466 32172 7472 32224
rect 7524 32212 7530 32224
rect 7837 32215 7895 32221
rect 7837 32212 7849 32215
rect 7524 32184 7849 32212
rect 7524 32172 7530 32184
rect 7837 32181 7849 32184
rect 7883 32181 7895 32215
rect 7837 32175 7895 32181
rect 10686 32172 10692 32224
rect 10744 32172 10750 32224
rect 12894 32172 12900 32224
rect 12952 32172 12958 32224
rect 13170 32172 13176 32224
rect 13228 32212 13234 32224
rect 14277 32215 14335 32221
rect 14277 32212 14289 32215
rect 13228 32184 14289 32212
rect 13228 32172 13234 32184
rect 14277 32181 14289 32184
rect 14323 32181 14335 32215
rect 14277 32175 14335 32181
rect 18230 32172 18236 32224
rect 18288 32172 18294 32224
rect 19886 32172 19892 32224
rect 19944 32212 19950 32224
rect 20073 32215 20131 32221
rect 20073 32212 20085 32215
rect 19944 32184 20085 32212
rect 19944 32172 19950 32184
rect 20073 32181 20085 32184
rect 20119 32181 20131 32215
rect 20073 32175 20131 32181
rect 20162 32172 20168 32224
rect 20220 32212 20226 32224
rect 20916 32212 20944 32252
rect 22278 32240 22284 32252
rect 22336 32240 22342 32292
rect 22756 32280 22784 32376
rect 23014 32308 23020 32360
rect 23072 32348 23078 32360
rect 23109 32351 23167 32357
rect 23109 32348 23121 32351
rect 23072 32320 23121 32348
rect 23072 32308 23078 32320
rect 23109 32317 23121 32320
rect 23155 32317 23167 32351
rect 23109 32311 23167 32317
rect 23293 32351 23351 32357
rect 23293 32317 23305 32351
rect 23339 32317 23351 32351
rect 23293 32311 23351 32317
rect 23308 32280 23336 32311
rect 23382 32308 23388 32360
rect 23440 32308 23446 32360
rect 23584 32348 23612 32379
rect 23842 32376 23848 32428
rect 23900 32376 23906 32428
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32385 23995 32419
rect 23937 32379 23995 32385
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32416 24087 32419
rect 24118 32416 24124 32428
rect 24075 32388 24124 32416
rect 24075 32385 24087 32388
rect 24029 32379 24087 32385
rect 23750 32348 23756 32360
rect 23584 32320 23756 32348
rect 22756 32252 23336 32280
rect 23584 32224 23612 32320
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 23952 32348 23980 32379
rect 24118 32376 24124 32388
rect 24176 32376 24182 32428
rect 24578 32376 24584 32428
rect 24636 32376 24642 32428
rect 24946 32376 24952 32428
rect 25004 32376 25010 32428
rect 25314 32376 25320 32428
rect 25372 32416 25378 32428
rect 25593 32419 25651 32425
rect 25593 32416 25605 32419
rect 25372 32388 25605 32416
rect 25372 32376 25378 32388
rect 25593 32385 25605 32388
rect 25639 32385 25651 32419
rect 25593 32379 25651 32385
rect 25682 32376 25688 32428
rect 25740 32376 25746 32428
rect 25792 32425 25820 32456
rect 26234 32444 26240 32496
rect 26292 32444 26298 32496
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32385 25835 32419
rect 25777 32379 25835 32385
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32385 26019 32419
rect 26252 32416 26280 32444
rect 26421 32419 26479 32425
rect 26421 32416 26433 32419
rect 26252 32388 26433 32416
rect 25961 32379 26019 32385
rect 26421 32385 26433 32388
rect 26467 32385 26479 32419
rect 26421 32379 26479 32385
rect 24964 32348 24992 32376
rect 23952 32320 24992 32348
rect 23952 32292 23980 32320
rect 25038 32308 25044 32360
rect 25096 32348 25102 32360
rect 25498 32348 25504 32360
rect 25096 32320 25504 32348
rect 25096 32308 25102 32320
rect 25498 32308 25504 32320
rect 25556 32348 25562 32360
rect 25976 32348 26004 32379
rect 25556 32320 26004 32348
rect 25556 32308 25562 32320
rect 23934 32240 23940 32292
rect 23992 32240 23998 32292
rect 24854 32240 24860 32292
rect 24912 32280 24918 32292
rect 26142 32280 26148 32292
rect 24912 32252 26148 32280
rect 24912 32240 24918 32252
rect 26142 32240 26148 32252
rect 26200 32240 26206 32292
rect 20220 32184 20944 32212
rect 21177 32215 21235 32221
rect 20220 32172 20226 32184
rect 21177 32181 21189 32215
rect 21223 32212 21235 32215
rect 21726 32212 21732 32224
rect 21223 32184 21732 32212
rect 21223 32181 21235 32184
rect 21177 32175 21235 32181
rect 21726 32172 21732 32184
rect 21784 32172 21790 32224
rect 22465 32215 22523 32221
rect 22465 32181 22477 32215
rect 22511 32212 22523 32215
rect 23474 32212 23480 32224
rect 22511 32184 23480 32212
rect 22511 32181 22523 32184
rect 22465 32175 22523 32181
rect 23474 32172 23480 32184
rect 23532 32172 23538 32224
rect 23566 32172 23572 32224
rect 23624 32172 23630 32224
rect 23842 32172 23848 32224
rect 23900 32212 23906 32224
rect 24213 32215 24271 32221
rect 24213 32212 24225 32215
rect 23900 32184 24225 32212
rect 23900 32172 23906 32184
rect 24213 32181 24225 32184
rect 24259 32181 24271 32215
rect 24213 32175 24271 32181
rect 25317 32215 25375 32221
rect 25317 32181 25329 32215
rect 25363 32212 25375 32215
rect 26234 32212 26240 32224
rect 25363 32184 26240 32212
rect 25363 32181 25375 32184
rect 25317 32175 25375 32181
rect 26234 32172 26240 32184
rect 26292 32172 26298 32224
rect 26436 32212 26464 32379
rect 26510 32308 26516 32360
rect 26568 32308 26574 32360
rect 26602 32308 26608 32360
rect 26660 32308 26666 32360
rect 26896 32348 26924 32524
rect 27154 32512 27160 32564
rect 27212 32512 27218 32564
rect 29086 32512 29092 32564
rect 29144 32552 29150 32564
rect 29638 32552 29644 32564
rect 29144 32524 29644 32552
rect 29144 32512 29150 32524
rect 29638 32512 29644 32524
rect 29696 32512 29702 32564
rect 30285 32555 30343 32561
rect 30285 32521 30297 32555
rect 30331 32521 30343 32555
rect 30285 32515 30343 32521
rect 27172 32484 27200 32512
rect 28534 32484 28540 32496
rect 26988 32456 27200 32484
rect 28474 32456 28540 32484
rect 26988 32425 27016 32456
rect 28534 32444 28540 32456
rect 28592 32444 28598 32496
rect 28626 32444 28632 32496
rect 28684 32484 28690 32496
rect 30009 32487 30067 32493
rect 30009 32484 30021 32487
rect 28684 32456 30021 32484
rect 28684 32444 28690 32456
rect 30009 32453 30021 32456
rect 30055 32484 30067 32487
rect 30190 32484 30196 32496
rect 30055 32456 30196 32484
rect 30055 32453 30067 32456
rect 30009 32447 30067 32453
rect 30190 32444 30196 32456
rect 30248 32444 30254 32496
rect 26973 32419 27031 32425
rect 26973 32385 26985 32419
rect 27019 32385 27031 32419
rect 26973 32379 27031 32385
rect 29638 32376 29644 32428
rect 29696 32376 29702 32428
rect 29730 32376 29736 32428
rect 29788 32416 29794 32428
rect 29917 32419 29975 32425
rect 29788 32388 29833 32416
rect 29788 32376 29794 32388
rect 29917 32385 29929 32419
rect 29963 32385 29975 32419
rect 29917 32379 29975 32385
rect 27249 32351 27307 32357
rect 27249 32348 27261 32351
rect 26896 32320 27261 32348
rect 27249 32317 27261 32320
rect 27295 32317 27307 32351
rect 27249 32311 27307 32317
rect 28994 32308 29000 32360
rect 29052 32308 29058 32360
rect 29932 32348 29960 32379
rect 30098 32376 30104 32428
rect 30156 32425 30162 32428
rect 30156 32416 30164 32425
rect 30300 32416 30328 32515
rect 30374 32512 30380 32564
rect 30432 32512 30438 32564
rect 30742 32512 30748 32564
rect 30800 32512 30806 32564
rect 31573 32555 31631 32561
rect 31573 32552 31585 32555
rect 30944 32524 31585 32552
rect 30392 32484 30420 32512
rect 30392 32456 30880 32484
rect 30852 32428 30880 32456
rect 30561 32419 30619 32425
rect 30561 32416 30573 32419
rect 30156 32388 30201 32416
rect 30300 32388 30573 32416
rect 30156 32379 30164 32388
rect 30561 32385 30573 32388
rect 30607 32385 30619 32419
rect 30561 32379 30619 32385
rect 30156 32376 30162 32379
rect 30834 32376 30840 32428
rect 30892 32376 30898 32428
rect 30006 32348 30012 32360
rect 29932 32320 30012 32348
rect 30006 32308 30012 32320
rect 30064 32308 30070 32360
rect 30944 32348 30972 32524
rect 31573 32521 31585 32524
rect 31619 32552 31631 32555
rect 32490 32552 32496 32564
rect 31619 32524 32496 32552
rect 31619 32521 31631 32524
rect 31573 32515 31631 32521
rect 32490 32512 32496 32524
rect 32548 32512 32554 32564
rect 34790 32552 34796 32564
rect 32692 32524 34796 32552
rect 31478 32444 31484 32496
rect 31536 32484 31542 32496
rect 31665 32487 31723 32493
rect 31665 32484 31677 32487
rect 31536 32456 31677 32484
rect 31536 32444 31542 32456
rect 31665 32453 31677 32456
rect 31711 32453 31723 32487
rect 31665 32447 31723 32453
rect 32692 32425 32720 32524
rect 34790 32512 34796 32524
rect 34848 32512 34854 32564
rect 35066 32512 35072 32564
rect 35124 32512 35130 32564
rect 33226 32444 33232 32496
rect 33284 32484 33290 32496
rect 35084 32484 35112 32512
rect 33284 32456 33442 32484
rect 34624 32456 35112 32484
rect 33284 32444 33290 32456
rect 32309 32419 32367 32425
rect 32309 32416 32321 32419
rect 30576 32320 30972 32348
rect 31772 32388 32321 32416
rect 29012 32212 29040 32308
rect 30576 32292 30604 32320
rect 30558 32240 30564 32292
rect 30616 32240 30622 32292
rect 31205 32283 31263 32289
rect 31205 32249 31217 32283
rect 31251 32280 31263 32283
rect 31772 32280 31800 32388
rect 32309 32385 32321 32388
rect 32355 32385 32367 32419
rect 32309 32379 32367 32385
rect 32677 32419 32735 32425
rect 32677 32385 32689 32419
rect 32723 32385 32735 32419
rect 32677 32379 32735 32385
rect 33962 32376 33968 32428
rect 34020 32376 34026 32428
rect 34624 32425 34652 32456
rect 34609 32419 34667 32425
rect 34609 32385 34621 32419
rect 34655 32385 34667 32419
rect 34609 32379 34667 32385
rect 35912 32388 36018 32416
rect 31849 32351 31907 32357
rect 31849 32317 31861 32351
rect 31895 32348 31907 32351
rect 32953 32351 33011 32357
rect 31895 32320 32260 32348
rect 31895 32317 31907 32320
rect 31849 32311 31907 32317
rect 31251 32252 31800 32280
rect 31251 32249 31263 32252
rect 31205 32243 31263 32249
rect 26436 32184 29040 32212
rect 30377 32215 30435 32221
rect 30377 32181 30389 32215
rect 30423 32212 30435 32215
rect 31478 32212 31484 32224
rect 30423 32184 31484 32212
rect 30423 32181 30435 32184
rect 30377 32175 30435 32181
rect 31478 32172 31484 32184
rect 31536 32172 31542 32224
rect 32122 32172 32128 32224
rect 32180 32172 32186 32224
rect 32232 32212 32260 32320
rect 32953 32317 32965 32351
rect 32999 32348 33011 32351
rect 33686 32348 33692 32360
rect 32999 32320 33692 32348
rect 32999 32317 33011 32320
rect 32953 32311 33011 32317
rect 33686 32308 33692 32320
rect 33744 32308 33750 32360
rect 33980 32280 34008 32376
rect 34238 32308 34244 32360
rect 34296 32348 34302 32360
rect 34885 32351 34943 32357
rect 34885 32348 34897 32351
rect 34296 32320 34897 32348
rect 34296 32308 34302 32320
rect 34885 32317 34897 32320
rect 34931 32317 34943 32351
rect 34885 32311 34943 32317
rect 34425 32283 34483 32289
rect 34425 32280 34437 32283
rect 33980 32252 34437 32280
rect 34425 32249 34437 32252
rect 34471 32249 34483 32283
rect 34425 32243 34483 32249
rect 35912 32224 35940 32388
rect 36630 32308 36636 32360
rect 36688 32308 36694 32360
rect 33962 32212 33968 32224
rect 32232 32184 33968 32212
rect 33962 32172 33968 32184
rect 34020 32172 34026 32224
rect 34146 32172 34152 32224
rect 34204 32212 34210 32224
rect 35894 32212 35900 32224
rect 34204 32184 35900 32212
rect 34204 32172 34210 32184
rect 35894 32172 35900 32184
rect 35952 32172 35958 32224
rect 1104 32122 38272 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38272 32122
rect 1104 32048 38272 32070
rect 6822 32008 6828 32020
rect 5736 31980 6828 32008
rect 3878 31764 3884 31816
rect 3936 31764 3942 31816
rect 5736 31804 5764 31980
rect 6822 31968 6828 31980
rect 6880 32008 6886 32020
rect 7834 32008 7840 32020
rect 6880 31980 7840 32008
rect 6880 31968 6886 31980
rect 7834 31968 7840 31980
rect 7892 31968 7898 32020
rect 8202 31968 8208 32020
rect 8260 32008 8266 32020
rect 11146 32008 11152 32020
rect 8260 31980 11152 32008
rect 8260 31968 8266 31980
rect 8018 31940 8024 31952
rect 7484 31912 8024 31940
rect 6089 31875 6147 31881
rect 6089 31841 6101 31875
rect 6135 31872 6147 31875
rect 7484 31872 7512 31912
rect 8018 31900 8024 31912
rect 8076 31900 8082 31952
rect 9398 31900 9404 31952
rect 9456 31900 9462 31952
rect 6135 31844 7512 31872
rect 7561 31875 7619 31881
rect 6135 31841 6147 31844
rect 6089 31835 6147 31841
rect 7561 31841 7573 31875
rect 7607 31872 7619 31875
rect 8938 31872 8944 31884
rect 7607 31844 7880 31872
rect 7607 31841 7619 31844
rect 7561 31835 7619 31841
rect 5290 31776 5764 31804
rect 4154 31696 4160 31748
rect 4212 31696 4218 31748
rect 5736 31736 5764 31776
rect 5810 31764 5816 31816
rect 5868 31764 5874 31816
rect 7852 31736 7880 31844
rect 7944 31844 8944 31872
rect 7944 31813 7972 31844
rect 8938 31832 8944 31844
rect 8996 31832 9002 31884
rect 7929 31807 7987 31813
rect 7929 31773 7941 31807
rect 7975 31773 7987 31807
rect 8113 31807 8171 31813
rect 8113 31804 8125 31807
rect 7929 31767 7987 31773
rect 8036 31776 8125 31804
rect 8036 31736 8064 31776
rect 8113 31773 8125 31776
rect 8159 31804 8171 31807
rect 9416 31804 9444 31900
rect 9508 31813 9536 31980
rect 11146 31968 11152 31980
rect 11204 32008 11210 32020
rect 11698 32008 11704 32020
rect 11204 31980 11704 32008
rect 11204 31968 11210 31980
rect 11698 31968 11704 31980
rect 11756 31968 11762 32020
rect 12710 31968 12716 32020
rect 12768 32008 12774 32020
rect 13449 32011 13507 32017
rect 13449 32008 13461 32011
rect 12768 31980 13461 32008
rect 12768 31968 12774 31980
rect 13449 31977 13461 31980
rect 13495 31977 13507 32011
rect 13449 31971 13507 31977
rect 18598 31968 18604 32020
rect 18656 32008 18662 32020
rect 20346 32008 20352 32020
rect 18656 31980 20352 32008
rect 18656 31968 18662 31980
rect 20346 31968 20352 31980
rect 20404 31968 20410 32020
rect 20732 31980 21864 32008
rect 20732 31952 20760 31980
rect 20622 31940 20628 31952
rect 19996 31912 20628 31940
rect 10226 31872 10232 31884
rect 10060 31844 10232 31872
rect 10060 31813 10088 31844
rect 10226 31832 10232 31844
rect 10284 31872 10290 31884
rect 10284 31844 11836 31872
rect 10284 31832 10290 31844
rect 8159 31776 9444 31804
rect 9493 31807 9551 31813
rect 8159 31773 8171 31776
rect 8113 31767 8171 31773
rect 9493 31773 9505 31807
rect 9539 31773 9551 31807
rect 9493 31767 9551 31773
rect 10045 31807 10103 31813
rect 10045 31773 10057 31807
rect 10091 31773 10103 31807
rect 10045 31767 10103 31773
rect 10137 31807 10195 31813
rect 10137 31773 10149 31807
rect 10183 31804 10195 31807
rect 10321 31807 10379 31813
rect 10321 31804 10333 31807
rect 10183 31776 10333 31804
rect 10183 31773 10195 31776
rect 10137 31767 10195 31773
rect 10321 31773 10333 31776
rect 10367 31773 10379 31807
rect 11808 31804 11836 31844
rect 12406 31844 14320 31872
rect 12406 31804 12434 31844
rect 11808 31776 12434 31804
rect 10321 31767 10379 31773
rect 12802 31764 12808 31816
rect 12860 31764 12866 31816
rect 12894 31764 12900 31816
rect 12952 31804 12958 31816
rect 13357 31807 13415 31813
rect 13357 31804 13369 31807
rect 12952 31776 13369 31804
rect 12952 31764 12958 31776
rect 13357 31773 13369 31776
rect 13403 31773 13415 31807
rect 13357 31767 13415 31773
rect 5736 31708 6578 31736
rect 7852 31708 8064 31736
rect 10594 31696 10600 31748
rect 10652 31696 10658 31748
rect 10870 31696 10876 31748
rect 10928 31736 10934 31748
rect 12820 31736 12848 31764
rect 14292 31748 14320 31844
rect 14734 31832 14740 31884
rect 14792 31872 14798 31884
rect 19996 31872 20024 31912
rect 20622 31900 20628 31912
rect 20680 31900 20686 31952
rect 20714 31900 20720 31952
rect 20772 31900 20778 31952
rect 20898 31900 20904 31952
rect 20956 31940 20962 31952
rect 21450 31940 21456 31952
rect 20956 31912 21456 31940
rect 20956 31900 20962 31912
rect 21450 31900 21456 31912
rect 21508 31900 21514 31952
rect 20346 31872 20352 31884
rect 14792 31844 20024 31872
rect 20272 31844 20352 31872
rect 14792 31832 14798 31844
rect 14369 31807 14427 31813
rect 14369 31773 14381 31807
rect 14415 31804 14427 31807
rect 14415 31776 15516 31804
rect 14415 31773 14427 31776
rect 14369 31767 14427 31773
rect 15488 31748 15516 31776
rect 16850 31764 16856 31816
rect 16908 31804 16914 31816
rect 17126 31804 17132 31816
rect 16908 31776 17132 31804
rect 16908 31764 16914 31776
rect 17126 31764 17132 31776
rect 17184 31804 17190 31816
rect 18877 31807 18935 31813
rect 17184 31776 18644 31804
rect 17184 31764 17190 31776
rect 13173 31739 13231 31745
rect 13173 31736 13185 31739
rect 10928 31708 11086 31736
rect 12820 31708 13185 31736
rect 10928 31696 10934 31708
rect 13173 31705 13185 31708
rect 13219 31705 13231 31739
rect 13173 31699 13231 31705
rect 14274 31696 14280 31748
rect 14332 31696 14338 31748
rect 14458 31696 14464 31748
rect 14516 31736 14522 31748
rect 14737 31739 14795 31745
rect 14737 31736 14749 31739
rect 14516 31708 14749 31736
rect 14516 31696 14522 31708
rect 14737 31705 14749 31708
rect 14783 31736 14795 31739
rect 14783 31708 15424 31736
rect 14783 31705 14795 31708
rect 14737 31699 14795 31705
rect 5629 31671 5687 31677
rect 5629 31637 5641 31671
rect 5675 31668 5687 31671
rect 6730 31668 6736 31680
rect 5675 31640 6736 31668
rect 5675 31637 5687 31640
rect 5629 31631 5687 31637
rect 6730 31628 6736 31640
rect 6788 31628 6794 31680
rect 7742 31628 7748 31680
rect 7800 31628 7806 31680
rect 8662 31628 8668 31680
rect 8720 31628 8726 31680
rect 9398 31628 9404 31680
rect 9456 31668 9462 31680
rect 9585 31671 9643 31677
rect 9585 31668 9597 31671
rect 9456 31640 9597 31668
rect 9456 31628 9462 31640
rect 9585 31637 9597 31640
rect 9631 31637 9643 31671
rect 9585 31631 9643 31637
rect 12066 31628 12072 31680
rect 12124 31628 12130 31680
rect 14366 31628 14372 31680
rect 14424 31668 14430 31680
rect 14553 31671 14611 31677
rect 14553 31668 14565 31671
rect 14424 31640 14565 31668
rect 14424 31628 14430 31640
rect 14553 31637 14565 31640
rect 14599 31637 14611 31671
rect 14553 31631 14611 31637
rect 14642 31628 14648 31680
rect 14700 31628 14706 31680
rect 14918 31628 14924 31680
rect 14976 31628 14982 31680
rect 15396 31668 15424 31708
rect 15470 31696 15476 31748
rect 15528 31696 15534 31748
rect 16298 31696 16304 31748
rect 16356 31736 16362 31748
rect 18616 31745 18644 31776
rect 18877 31773 18889 31807
rect 18923 31804 18935 31807
rect 19058 31804 19064 31816
rect 18923 31776 19064 31804
rect 18923 31773 18935 31776
rect 18877 31767 18935 31773
rect 19058 31764 19064 31776
rect 19116 31804 19122 31816
rect 19978 31804 19984 31816
rect 19116 31776 19984 31804
rect 19116 31764 19122 31776
rect 19978 31764 19984 31776
rect 20036 31764 20042 31816
rect 20272 31813 20300 31844
rect 20346 31832 20352 31844
rect 20404 31832 20410 31884
rect 20530 31832 20536 31884
rect 20588 31872 20594 31884
rect 20806 31872 20812 31884
rect 20588 31844 20812 31872
rect 20588 31832 20594 31844
rect 20806 31832 20812 31844
rect 20864 31832 20870 31884
rect 21174 31832 21180 31884
rect 21232 31872 21238 31884
rect 21836 31881 21864 31980
rect 22554 31968 22560 32020
rect 22612 32008 22618 32020
rect 23293 32011 23351 32017
rect 22612 31980 22932 32008
rect 22612 31968 22618 31980
rect 22904 31940 22932 31980
rect 23293 31977 23305 32011
rect 23339 32008 23351 32011
rect 23750 32008 23756 32020
rect 23339 31980 23756 32008
rect 23339 31977 23351 31980
rect 23293 31971 23351 31977
rect 23750 31968 23756 31980
rect 23808 31968 23814 32020
rect 25961 32011 26019 32017
rect 25961 31977 25973 32011
rect 26007 32008 26019 32011
rect 26050 32008 26056 32020
rect 26007 31980 26056 32008
rect 26007 31977 26019 31980
rect 25961 31971 26019 31977
rect 26050 31968 26056 31980
rect 26108 31968 26114 32020
rect 26234 31968 26240 32020
rect 26292 32008 26298 32020
rect 27154 32008 27160 32020
rect 26292 31980 27160 32008
rect 26292 31968 26298 31980
rect 27154 31968 27160 31980
rect 27212 32008 27218 32020
rect 27982 32008 27988 32020
rect 27212 31980 27988 32008
rect 27212 31968 27218 31980
rect 27982 31968 27988 31980
rect 28040 31968 28046 32020
rect 28350 31968 28356 32020
rect 28408 32008 28414 32020
rect 28408 31980 28994 32008
rect 28408 31968 28414 31980
rect 28966 31940 28994 31980
rect 30742 31968 30748 32020
rect 30800 31968 30806 32020
rect 31468 32011 31526 32017
rect 31468 31977 31480 32011
rect 31514 32008 31526 32011
rect 32122 32008 32128 32020
rect 31514 31980 32128 32008
rect 31514 31977 31526 31980
rect 31468 31971 31526 31977
rect 32122 31968 32128 31980
rect 32180 31968 32186 32020
rect 32490 31968 32496 32020
rect 32548 31968 32554 32020
rect 33594 31968 33600 32020
rect 33652 32008 33658 32020
rect 34146 32008 34152 32020
rect 33652 31980 34152 32008
rect 33652 31968 33658 31980
rect 34146 31968 34152 31980
rect 34204 31968 34210 32020
rect 34238 31968 34244 32020
rect 34296 31968 34302 32020
rect 30558 31940 30564 31952
rect 22904 31912 23152 31940
rect 28966 31912 30564 31940
rect 21729 31875 21787 31881
rect 21729 31872 21741 31875
rect 21232 31844 21741 31872
rect 21232 31832 21238 31844
rect 21729 31841 21741 31844
rect 21775 31841 21787 31875
rect 21729 31835 21787 31841
rect 21821 31875 21879 31881
rect 21821 31841 21833 31875
rect 21867 31872 21879 31875
rect 22002 31872 22008 31884
rect 21867 31844 22008 31872
rect 21867 31841 21879 31844
rect 21821 31835 21879 31841
rect 22002 31832 22008 31844
rect 22060 31872 22066 31884
rect 22060 31844 23060 31872
rect 22060 31832 22066 31844
rect 20257 31807 20315 31813
rect 20257 31773 20269 31807
rect 20303 31773 20315 31807
rect 21085 31807 21143 31813
rect 21085 31804 21097 31807
rect 20257 31767 20315 31773
rect 21008 31776 21097 31804
rect 21008 31748 21036 31776
rect 21085 31773 21097 31776
rect 21131 31804 21143 31807
rect 21637 31807 21695 31813
rect 21637 31804 21649 31807
rect 21131 31776 21649 31804
rect 21131 31773 21143 31776
rect 21085 31767 21143 31773
rect 21637 31773 21649 31776
rect 21683 31773 21695 31807
rect 21637 31767 21695 31773
rect 21913 31807 21971 31813
rect 21913 31773 21925 31807
rect 21959 31773 21971 31807
rect 21913 31767 21971 31773
rect 18417 31739 18475 31745
rect 18417 31736 18429 31739
rect 16356 31708 18429 31736
rect 16356 31696 16362 31708
rect 18417 31705 18429 31708
rect 18463 31705 18475 31739
rect 18417 31699 18475 31705
rect 18601 31739 18659 31745
rect 18601 31705 18613 31739
rect 18647 31705 18659 31739
rect 18601 31699 18659 31705
rect 18966 31696 18972 31748
rect 19024 31736 19030 31748
rect 19024 31708 20484 31736
rect 19024 31696 19030 31708
rect 18782 31668 18788 31680
rect 15396 31640 18788 31668
rect 18782 31628 18788 31640
rect 18840 31628 18846 31680
rect 19794 31628 19800 31680
rect 19852 31668 19858 31680
rect 20346 31668 20352 31680
rect 19852 31640 20352 31668
rect 19852 31628 19858 31640
rect 20346 31628 20352 31640
rect 20404 31628 20410 31680
rect 20456 31668 20484 31708
rect 20990 31696 20996 31748
rect 21048 31696 21054 31748
rect 21174 31668 21180 31680
rect 20456 31640 21180 31668
rect 21174 31628 21180 31640
rect 21232 31628 21238 31680
rect 21266 31628 21272 31680
rect 21324 31668 21330 31680
rect 21453 31671 21511 31677
rect 21453 31668 21465 31671
rect 21324 31640 21465 31668
rect 21324 31628 21330 31640
rect 21453 31637 21465 31640
rect 21499 31637 21511 31671
rect 21453 31631 21511 31637
rect 21634 31628 21640 31680
rect 21692 31668 21698 31680
rect 21928 31668 21956 31767
rect 22186 31764 22192 31816
rect 22244 31804 22250 31816
rect 22554 31804 22560 31816
rect 22244 31776 22560 31804
rect 22244 31764 22250 31776
rect 22554 31764 22560 31776
rect 22612 31764 22618 31816
rect 22738 31764 22744 31816
rect 22796 31764 22802 31816
rect 23032 31813 23060 31844
rect 23124 31813 23152 31912
rect 30558 31900 30564 31912
rect 30616 31900 30622 31952
rect 24946 31832 24952 31884
rect 25004 31872 25010 31884
rect 25004 31844 26188 31872
rect 25004 31832 25010 31844
rect 23017 31807 23075 31813
rect 23017 31773 23029 31807
rect 23063 31773 23075 31807
rect 23017 31767 23075 31773
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31804 23167 31807
rect 23382 31804 23388 31816
rect 23155 31776 23388 31804
rect 23155 31773 23167 31776
rect 23109 31767 23167 31773
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 24578 31764 24584 31816
rect 24636 31804 24642 31816
rect 25700 31813 25728 31844
rect 25409 31807 25467 31813
rect 25409 31804 25421 31807
rect 24636 31776 25421 31804
rect 24636 31764 24642 31776
rect 22925 31739 22983 31745
rect 22925 31705 22937 31739
rect 22971 31736 22983 31739
rect 22971 31708 23152 31736
rect 22971 31705 22983 31708
rect 22925 31699 22983 31705
rect 23124 31680 23152 31708
rect 21692 31640 21956 31668
rect 21692 31628 21698 31640
rect 22462 31628 22468 31680
rect 22520 31668 22526 31680
rect 23014 31668 23020 31680
rect 22520 31640 23020 31668
rect 22520 31628 22526 31640
rect 23014 31628 23020 31640
rect 23072 31628 23078 31680
rect 23106 31628 23112 31680
rect 23164 31628 23170 31680
rect 25148 31668 25176 31776
rect 25409 31773 25421 31776
rect 25455 31773 25467 31807
rect 25409 31767 25467 31773
rect 25593 31807 25651 31813
rect 25593 31773 25605 31807
rect 25639 31773 25651 31807
rect 25593 31767 25651 31773
rect 25685 31807 25743 31813
rect 25685 31773 25697 31807
rect 25731 31773 25743 31807
rect 25685 31767 25743 31773
rect 25777 31807 25835 31813
rect 25777 31773 25789 31807
rect 25823 31804 25835 31807
rect 25866 31804 25872 31816
rect 25823 31776 25872 31804
rect 25823 31773 25835 31776
rect 25777 31767 25835 31773
rect 25222 31696 25228 31748
rect 25280 31736 25286 31748
rect 25498 31736 25504 31748
rect 25280 31708 25504 31736
rect 25280 31696 25286 31708
rect 25498 31696 25504 31708
rect 25556 31736 25562 31748
rect 25608 31736 25636 31767
rect 25866 31764 25872 31776
rect 25924 31804 25930 31816
rect 26050 31804 26056 31816
rect 25924 31776 26056 31804
rect 25924 31764 25930 31776
rect 26050 31764 26056 31776
rect 26108 31764 26114 31816
rect 26160 31804 26188 31844
rect 28994 31832 29000 31884
rect 29052 31872 29058 31884
rect 29825 31875 29883 31881
rect 29825 31872 29837 31875
rect 29052 31844 29837 31872
rect 29052 31832 29058 31844
rect 29825 31841 29837 31844
rect 29871 31841 29883 31875
rect 30760 31872 30788 31968
rect 29825 31835 29883 31841
rect 29932 31844 30788 31872
rect 29932 31804 29960 31844
rect 31110 31832 31116 31884
rect 31168 31832 31174 31884
rect 31205 31875 31263 31881
rect 31205 31841 31217 31875
rect 31251 31872 31263 31875
rect 31846 31872 31852 31884
rect 31251 31844 31852 31872
rect 31251 31841 31263 31844
rect 31205 31835 31263 31841
rect 31846 31832 31852 31844
rect 31904 31832 31910 31884
rect 32508 31872 32536 31968
rect 33413 31943 33471 31949
rect 33413 31909 33425 31943
rect 33459 31940 33471 31943
rect 33459 31912 34468 31940
rect 33459 31909 33471 31912
rect 33413 31903 33471 31909
rect 33229 31875 33287 31881
rect 33229 31872 33241 31875
rect 32508 31844 33241 31872
rect 33229 31841 33241 31844
rect 33275 31841 33287 31875
rect 33229 31835 33287 31841
rect 33594 31832 33600 31884
rect 33652 31832 33658 31884
rect 33962 31832 33968 31884
rect 34020 31832 34026 31884
rect 26160 31776 29960 31804
rect 30190 31764 30196 31816
rect 30248 31764 30254 31816
rect 30374 31764 30380 31816
rect 30432 31764 30438 31816
rect 30466 31764 30472 31816
rect 30524 31804 30530 31816
rect 30745 31807 30803 31813
rect 30745 31804 30757 31807
rect 30524 31776 30757 31804
rect 30524 31764 30530 31776
rect 30745 31773 30757 31776
rect 30791 31773 30803 31807
rect 33612 31804 33640 31832
rect 34440 31813 34468 31912
rect 33873 31807 33931 31813
rect 33873 31804 33885 31807
rect 33612 31776 33885 31804
rect 30745 31767 30803 31773
rect 33873 31773 33885 31776
rect 33919 31773 33931 31807
rect 33873 31767 33931 31773
rect 34425 31807 34483 31813
rect 34425 31773 34437 31807
rect 34471 31773 34483 31807
rect 34425 31767 34483 31773
rect 25556 31708 25636 31736
rect 25556 31696 25562 31708
rect 28626 31696 28632 31748
rect 28684 31696 28690 31748
rect 29012 31708 31248 31736
rect 28644 31668 28672 31696
rect 29012 31680 29040 31708
rect 25148 31640 28672 31668
rect 28994 31628 29000 31680
rect 29052 31628 29058 31680
rect 31220 31668 31248 31708
rect 31754 31696 31760 31748
rect 31812 31736 31818 31748
rect 31812 31708 31970 31736
rect 31812 31696 31818 31708
rect 33781 31671 33839 31677
rect 33781 31668 33793 31671
rect 31220 31640 33793 31668
rect 33781 31637 33793 31640
rect 33827 31668 33839 31671
rect 36630 31668 36636 31680
rect 33827 31640 36636 31668
rect 33827 31637 33839 31640
rect 33781 31631 33839 31637
rect 36630 31628 36636 31640
rect 36688 31628 36694 31680
rect 1104 31578 38272 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38272 31578
rect 1104 31504 38272 31526
rect 3878 31424 3884 31476
rect 3936 31464 3942 31476
rect 4065 31467 4123 31473
rect 4065 31464 4077 31467
rect 3936 31436 4077 31464
rect 3936 31424 3942 31436
rect 4065 31433 4077 31436
rect 4111 31433 4123 31467
rect 4065 31427 4123 31433
rect 4154 31424 4160 31476
rect 4212 31464 4218 31476
rect 4893 31467 4951 31473
rect 4893 31464 4905 31467
rect 4212 31436 4905 31464
rect 4212 31424 4218 31436
rect 4893 31433 4905 31436
rect 4939 31433 4951 31467
rect 4893 31427 4951 31433
rect 5810 31424 5816 31476
rect 5868 31464 5874 31476
rect 5997 31467 6055 31473
rect 5997 31464 6009 31467
rect 5868 31436 6009 31464
rect 5868 31424 5874 31436
rect 5997 31433 6009 31436
rect 6043 31433 6055 31467
rect 5997 31427 6055 31433
rect 6730 31424 6736 31476
rect 6788 31424 6794 31476
rect 6825 31467 6883 31473
rect 6825 31433 6837 31467
rect 6871 31464 6883 31467
rect 8110 31464 8116 31476
rect 6871 31436 8116 31464
rect 6871 31433 6883 31436
rect 6825 31427 6883 31433
rect 8110 31424 8116 31436
rect 8168 31424 8174 31476
rect 11514 31424 11520 31476
rect 11572 31424 11578 31476
rect 14274 31424 14280 31476
rect 14332 31424 14338 31476
rect 18693 31467 18751 31473
rect 18693 31433 18705 31467
rect 18739 31433 18751 31467
rect 18693 31427 18751 31433
rect 20717 31467 20775 31473
rect 20717 31433 20729 31467
rect 20763 31433 20775 31467
rect 20717 31427 20775 31433
rect 3988 31368 5396 31396
rect 3988 31337 4016 31368
rect 5368 31340 5396 31368
rect 7742 31356 7748 31408
rect 7800 31356 7806 31408
rect 7834 31356 7840 31408
rect 7892 31396 7898 31408
rect 7892 31368 8234 31396
rect 7892 31356 7898 31368
rect 16574 31356 16580 31408
rect 16632 31396 16638 31408
rect 16669 31399 16727 31405
rect 16669 31396 16681 31399
rect 16632 31368 16681 31396
rect 16632 31356 16638 31368
rect 16669 31365 16681 31368
rect 16715 31396 16727 31399
rect 16942 31396 16948 31408
rect 16715 31368 16948 31396
rect 16715 31365 16727 31368
rect 16669 31359 16727 31365
rect 16942 31356 16948 31368
rect 17000 31356 17006 31408
rect 17313 31399 17371 31405
rect 17052 31368 17264 31396
rect 3973 31331 4031 31337
rect 3973 31297 3985 31331
rect 4019 31297 4031 31331
rect 3973 31291 4031 31297
rect 5077 31331 5135 31337
rect 5077 31297 5089 31331
rect 5123 31297 5135 31331
rect 5077 31291 5135 31297
rect 5092 31260 5120 31291
rect 5350 31288 5356 31340
rect 5408 31288 5414 31340
rect 5534 31288 5540 31340
rect 5592 31328 5598 31340
rect 5905 31331 5963 31337
rect 5905 31328 5917 31331
rect 5592 31300 5917 31328
rect 5592 31288 5598 31300
rect 5905 31297 5917 31300
rect 5951 31328 5963 31331
rect 6638 31328 6644 31340
rect 5951 31300 6644 31328
rect 5951 31297 5963 31300
rect 5905 31291 5963 31297
rect 6638 31288 6644 31300
rect 6696 31288 6702 31340
rect 7466 31288 7472 31340
rect 7524 31288 7530 31340
rect 11885 31331 11943 31337
rect 11885 31328 11897 31331
rect 5092 31232 6408 31260
rect 6380 31201 6408 31232
rect 6454 31220 6460 31272
rect 6512 31260 6518 31272
rect 6822 31260 6828 31272
rect 6512 31232 6828 31260
rect 6512 31220 6518 31232
rect 6822 31220 6828 31232
rect 6880 31260 6886 31272
rect 6917 31263 6975 31269
rect 6917 31260 6929 31263
rect 6880 31232 6929 31260
rect 6880 31220 6886 31232
rect 6917 31229 6929 31232
rect 6963 31229 6975 31263
rect 6917 31223 6975 31229
rect 9398 31220 9404 31272
rect 9456 31220 9462 31272
rect 9674 31220 9680 31272
rect 9732 31220 9738 31272
rect 10796 31260 10824 31314
rect 11072 31300 11897 31328
rect 10870 31260 10876 31272
rect 10796 31232 10876 31260
rect 10870 31220 10876 31232
rect 10928 31220 10934 31272
rect 6365 31195 6423 31201
rect 6365 31161 6377 31195
rect 6411 31161 6423 31195
rect 6365 31155 6423 31161
rect 11072 31136 11100 31300
rect 11885 31297 11897 31300
rect 11931 31297 11943 31331
rect 11885 31291 11943 31297
rect 12989 31331 13047 31337
rect 12989 31297 13001 31331
rect 13035 31328 13047 31331
rect 13722 31328 13728 31340
rect 13035 31300 13728 31328
rect 13035 31297 13047 31300
rect 12989 31291 13047 31297
rect 13722 31288 13728 31300
rect 13780 31328 13786 31340
rect 15286 31328 15292 31340
rect 13780 31300 15292 31328
rect 13780 31288 13786 31300
rect 15286 31288 15292 31300
rect 15344 31288 15350 31340
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 11977 31263 12035 31269
rect 11977 31229 11989 31263
rect 12023 31260 12035 31263
rect 12066 31260 12072 31272
rect 12023 31232 12072 31260
rect 12023 31229 12035 31232
rect 11977 31223 12035 31229
rect 12066 31220 12072 31232
rect 12124 31220 12130 31272
rect 12158 31220 12164 31272
rect 12216 31220 12222 31272
rect 16574 31220 16580 31272
rect 16632 31260 16638 31272
rect 16868 31260 16896 31291
rect 16632 31232 16896 31260
rect 16632 31220 16638 31232
rect 16942 31220 16948 31272
rect 17000 31260 17006 31272
rect 17052 31260 17080 31368
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31297 17187 31331
rect 17236 31328 17264 31368
rect 17313 31365 17325 31399
rect 17359 31396 17371 31399
rect 17586 31396 17592 31408
rect 17359 31368 17592 31396
rect 17359 31365 17371 31368
rect 17313 31359 17371 31365
rect 17586 31356 17592 31368
rect 17644 31356 17650 31408
rect 18708 31340 18736 31427
rect 18874 31356 18880 31408
rect 18932 31396 18938 31408
rect 19429 31399 19487 31405
rect 18932 31368 19334 31396
rect 18932 31356 18938 31368
rect 17405 31331 17463 31337
rect 17405 31328 17417 31331
rect 17236 31300 17417 31328
rect 17129 31291 17187 31297
rect 17405 31297 17417 31300
rect 17451 31297 17463 31331
rect 17405 31291 17463 31297
rect 17000 31232 17080 31260
rect 17000 31220 17006 31232
rect 17144 31192 17172 31291
rect 17494 31288 17500 31340
rect 17552 31288 17558 31340
rect 18598 31328 18604 31340
rect 17650 31300 18604 31328
rect 17650 31260 17678 31300
rect 18598 31288 18604 31300
rect 18656 31288 18662 31340
rect 18690 31288 18696 31340
rect 18748 31288 18754 31340
rect 19150 31288 19156 31340
rect 19208 31288 19214 31340
rect 19306 31328 19334 31368
rect 19429 31365 19441 31399
rect 19475 31396 19487 31399
rect 20530 31396 20536 31408
rect 19475 31368 20536 31396
rect 19475 31365 19487 31368
rect 19429 31359 19487 31365
rect 20530 31356 20536 31368
rect 20588 31356 20594 31408
rect 20732 31340 20760 31427
rect 20806 31424 20812 31476
rect 20864 31464 20870 31476
rect 22002 31464 22008 31476
rect 20864 31436 22008 31464
rect 20864 31424 20870 31436
rect 22002 31424 22008 31436
rect 22060 31464 22066 31476
rect 22557 31467 22615 31473
rect 22060 31436 22508 31464
rect 22060 31424 22066 31436
rect 22094 31356 22100 31408
rect 22152 31396 22158 31408
rect 22373 31399 22431 31405
rect 22373 31396 22385 31399
rect 22152 31368 22385 31396
rect 22152 31356 22158 31368
rect 22373 31365 22385 31368
rect 22419 31365 22431 31399
rect 22373 31359 22431 31365
rect 19886 31328 19892 31340
rect 19306 31300 19892 31328
rect 19886 31288 19892 31300
rect 19944 31288 19950 31340
rect 20714 31288 20720 31340
rect 20772 31288 20778 31340
rect 20898 31288 20904 31340
rect 20956 31328 20962 31340
rect 21542 31328 21548 31340
rect 20956 31300 21548 31328
rect 20956 31288 20962 31300
rect 21542 31288 21548 31300
rect 21600 31328 21606 31340
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 21600 31300 22201 31328
rect 21600 31288 21606 31300
rect 22189 31297 22201 31300
rect 22235 31297 22247 31331
rect 22480 31328 22508 31436
rect 22557 31433 22569 31467
rect 22603 31464 22615 31467
rect 22603 31436 22876 31464
rect 22603 31433 22615 31436
rect 22557 31427 22615 31433
rect 22848 31337 22876 31436
rect 22922 31424 22928 31476
rect 22980 31464 22986 31476
rect 23290 31464 23296 31476
rect 22980 31436 23296 31464
rect 22980 31424 22986 31436
rect 23290 31424 23296 31436
rect 23348 31424 23354 31476
rect 24210 31424 24216 31476
rect 24268 31464 24274 31476
rect 28810 31464 28816 31476
rect 24268 31436 28816 31464
rect 24268 31424 24274 31436
rect 28810 31424 28816 31436
rect 28868 31464 28874 31476
rect 28994 31464 29000 31476
rect 28868 31436 29000 31464
rect 28868 31424 28874 31436
rect 28994 31424 29000 31436
rect 29052 31424 29058 31476
rect 29549 31467 29607 31473
rect 29549 31433 29561 31467
rect 29595 31433 29607 31467
rect 29549 31427 29607 31433
rect 25682 31396 25688 31408
rect 25240 31368 25688 31396
rect 22649 31331 22707 31337
rect 22649 31328 22661 31331
rect 22480 31300 22661 31328
rect 22189 31291 22247 31297
rect 22649 31297 22661 31300
rect 22695 31297 22707 31331
rect 22649 31291 22707 31297
rect 22833 31331 22891 31337
rect 22833 31297 22845 31331
rect 22879 31297 22891 31331
rect 22833 31291 22891 31297
rect 22922 31288 22928 31340
rect 22980 31288 22986 31340
rect 23014 31288 23020 31340
rect 23072 31328 23078 31340
rect 23290 31328 23296 31340
rect 23072 31300 23296 31328
rect 23072 31288 23078 31300
rect 23290 31288 23296 31300
rect 23348 31288 23354 31340
rect 25240 31337 25268 31368
rect 25682 31356 25688 31368
rect 25740 31356 25746 31408
rect 25866 31356 25872 31408
rect 25924 31396 25930 31408
rect 25924 31368 28028 31396
rect 25924 31356 25930 31368
rect 28000 31340 28028 31368
rect 28626 31356 28632 31408
rect 28684 31396 28690 31408
rect 29564 31396 29592 31427
rect 30190 31424 30196 31476
rect 30248 31464 30254 31476
rect 31294 31464 31300 31476
rect 30248 31436 31300 31464
rect 30248 31424 30254 31436
rect 31294 31424 31300 31436
rect 31352 31424 31358 31476
rect 31757 31467 31815 31473
rect 31757 31433 31769 31467
rect 31803 31464 31815 31467
rect 31846 31464 31852 31476
rect 31803 31436 31852 31464
rect 31803 31433 31815 31436
rect 31757 31427 31815 31433
rect 31846 31424 31852 31436
rect 31904 31424 31910 31476
rect 28684 31368 29592 31396
rect 30484 31368 31708 31396
rect 28684 31356 28690 31368
rect 23385 31331 23443 31337
rect 23385 31297 23397 31331
rect 23431 31297 23443 31331
rect 25225 31331 25283 31337
rect 25225 31328 25237 31331
rect 23385 31291 23443 31297
rect 23860 31300 25237 31328
rect 17420 31232 17678 31260
rect 17420 31204 17448 31232
rect 18138 31220 18144 31272
rect 18196 31260 18202 31272
rect 20254 31260 20260 31272
rect 18196 31232 20260 31260
rect 18196 31220 18202 31232
rect 20254 31220 20260 31232
rect 20312 31220 20318 31272
rect 20622 31220 20628 31272
rect 20680 31260 20686 31272
rect 23400 31260 23428 31291
rect 23860 31272 23888 31300
rect 25225 31297 25237 31300
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 26142 31288 26148 31340
rect 26200 31328 26206 31340
rect 27890 31328 27896 31340
rect 26200 31300 27896 31328
rect 26200 31288 26206 31300
rect 27890 31288 27896 31300
rect 27948 31288 27954 31340
rect 27982 31288 27988 31340
rect 28040 31288 28046 31340
rect 28074 31288 28080 31340
rect 28132 31288 28138 31340
rect 28258 31288 28264 31340
rect 28316 31288 28322 31340
rect 28810 31288 28816 31340
rect 28868 31326 28874 31340
rect 28905 31331 28963 31337
rect 28905 31326 28917 31331
rect 28868 31298 28917 31326
rect 28868 31288 28874 31298
rect 28905 31297 28917 31298
rect 28951 31297 28963 31331
rect 28905 31291 28963 31297
rect 28994 31288 29000 31340
rect 29052 31288 29058 31340
rect 29086 31288 29092 31340
rect 29144 31288 29150 31340
rect 29270 31288 29276 31340
rect 29328 31288 29334 31340
rect 29365 31331 29423 31337
rect 29365 31297 29377 31331
rect 29411 31328 29423 31331
rect 29914 31328 29920 31340
rect 29411 31300 29920 31328
rect 29411 31297 29423 31300
rect 29365 31291 29423 31297
rect 20680 31232 23428 31260
rect 20680 31220 20686 31232
rect 23842 31220 23848 31272
rect 23900 31220 23906 31272
rect 27062 31220 27068 31272
rect 27120 31260 27126 31272
rect 29380 31260 29408 31291
rect 29914 31288 29920 31300
rect 29972 31328 29978 31340
rect 30484 31337 30512 31368
rect 30469 31331 30527 31337
rect 30469 31328 30481 31331
rect 29972 31300 30481 31328
rect 29972 31288 29978 31300
rect 30469 31297 30481 31300
rect 30515 31297 30527 31331
rect 30469 31291 30527 31297
rect 30558 31288 30564 31340
rect 30616 31328 30622 31340
rect 31205 31331 31263 31337
rect 31205 31328 31217 31331
rect 30616 31300 31217 31328
rect 30616 31288 30622 31300
rect 31205 31297 31217 31300
rect 31251 31297 31263 31331
rect 31205 31291 31263 31297
rect 31294 31288 31300 31340
rect 31352 31288 31358 31340
rect 31389 31331 31447 31337
rect 31389 31297 31401 31331
rect 31435 31297 31447 31331
rect 31389 31291 31447 31297
rect 31404 31260 31432 31291
rect 31570 31288 31576 31340
rect 31628 31288 31634 31340
rect 31680 31337 31708 31368
rect 31665 31331 31723 31337
rect 31665 31297 31677 31331
rect 31711 31297 31723 31331
rect 31665 31291 31723 31297
rect 32306 31288 32312 31340
rect 32364 31288 32370 31340
rect 34606 31288 34612 31340
rect 34664 31328 34670 31340
rect 34793 31331 34851 31337
rect 34793 31328 34805 31331
rect 34664 31300 34805 31328
rect 34664 31288 34670 31300
rect 34793 31297 34805 31300
rect 34839 31297 34851 31331
rect 34793 31291 34851 31297
rect 27120 31232 29408 31260
rect 30852 31232 31432 31260
rect 27120 31220 27126 31232
rect 16224 31164 17172 31192
rect 16224 31136 16252 31164
rect 9214 31084 9220 31136
rect 9272 31084 9278 31136
rect 11054 31084 11060 31136
rect 11112 31084 11118 31136
rect 11149 31127 11207 31133
rect 11149 31093 11161 31127
rect 11195 31124 11207 31127
rect 11238 31124 11244 31136
rect 11195 31096 11244 31124
rect 11195 31093 11207 31096
rect 11149 31087 11207 31093
rect 11238 31084 11244 31096
rect 11296 31084 11302 31136
rect 11514 31084 11520 31136
rect 11572 31124 11578 31136
rect 13262 31124 13268 31136
rect 11572 31096 13268 31124
rect 11572 31084 11578 31096
rect 13262 31084 13268 31096
rect 13320 31084 13326 31136
rect 16206 31084 16212 31136
rect 16264 31084 16270 31136
rect 17034 31084 17040 31136
rect 17092 31084 17098 31136
rect 17144 31124 17172 31164
rect 17402 31152 17408 31204
rect 17460 31152 17466 31204
rect 17604 31164 17908 31192
rect 17604 31124 17632 31164
rect 17144 31096 17632 31124
rect 17678 31084 17684 31136
rect 17736 31084 17742 31136
rect 17880 31124 17908 31164
rect 17954 31152 17960 31204
rect 18012 31192 18018 31204
rect 30653 31195 30711 31201
rect 30653 31192 30665 31195
rect 18012 31164 30665 31192
rect 18012 31152 18018 31164
rect 30653 31161 30665 31164
rect 30699 31161 30711 31195
rect 30653 31155 30711 31161
rect 18230 31124 18236 31136
rect 17880 31096 18236 31124
rect 18230 31084 18236 31096
rect 18288 31084 18294 31136
rect 18414 31084 18420 31136
rect 18472 31124 18478 31136
rect 19334 31124 19340 31136
rect 18472 31096 19340 31124
rect 18472 31084 18478 31096
rect 19334 31084 19340 31096
rect 19392 31084 19398 31136
rect 20622 31084 20628 31136
rect 20680 31124 20686 31136
rect 20990 31124 20996 31136
rect 20680 31096 20996 31124
rect 20680 31084 20686 31096
rect 20990 31084 20996 31096
rect 21048 31084 21054 31136
rect 21450 31084 21456 31136
rect 21508 31124 21514 31136
rect 22922 31124 22928 31136
rect 21508 31096 22928 31124
rect 21508 31084 21514 31096
rect 22922 31084 22928 31096
rect 22980 31084 22986 31136
rect 23198 31084 23204 31136
rect 23256 31084 23262 31136
rect 24026 31084 24032 31136
rect 24084 31124 24090 31136
rect 24673 31127 24731 31133
rect 24673 31124 24685 31127
rect 24084 31096 24685 31124
rect 24084 31084 24090 31096
rect 24673 31093 24685 31096
rect 24719 31093 24731 31127
rect 24673 31087 24731 31093
rect 25222 31084 25228 31136
rect 25280 31084 25286 31136
rect 25590 31084 25596 31136
rect 25648 31084 25654 31136
rect 27617 31127 27675 31133
rect 27617 31093 27629 31127
rect 27663 31124 27675 31127
rect 27706 31124 27712 31136
rect 27663 31096 27712 31124
rect 27663 31093 27675 31096
rect 27617 31087 27675 31093
rect 27706 31084 27712 31096
rect 27764 31084 27770 31136
rect 28074 31084 28080 31136
rect 28132 31124 28138 31136
rect 28629 31127 28687 31133
rect 28629 31124 28641 31127
rect 28132 31096 28641 31124
rect 28132 31084 28138 31096
rect 28629 31093 28641 31096
rect 28675 31093 28687 31127
rect 28629 31087 28687 31093
rect 28810 31084 28816 31136
rect 28868 31124 28874 31136
rect 29270 31124 29276 31136
rect 28868 31096 29276 31124
rect 28868 31084 28874 31096
rect 29270 31084 29276 31096
rect 29328 31124 29334 31136
rect 30466 31124 30472 31136
rect 29328 31096 30472 31124
rect 29328 31084 29334 31096
rect 30466 31084 30472 31096
rect 30524 31124 30530 31136
rect 30852 31124 30880 31232
rect 30524 31096 30880 31124
rect 30929 31127 30987 31133
rect 30524 31084 30530 31096
rect 30929 31093 30941 31127
rect 30975 31124 30987 31127
rect 32030 31124 32036 31136
rect 30975 31096 32036 31124
rect 30975 31093 30987 31096
rect 30929 31087 30987 31093
rect 32030 31084 32036 31096
rect 32088 31084 32094 31136
rect 32125 31127 32183 31133
rect 32125 31093 32137 31127
rect 32171 31124 32183 31127
rect 32398 31124 32404 31136
rect 32171 31096 32404 31124
rect 32171 31093 32183 31096
rect 32125 31087 32183 31093
rect 32398 31084 32404 31096
rect 32456 31084 32462 31136
rect 34790 31084 34796 31136
rect 34848 31124 34854 31136
rect 34885 31127 34943 31133
rect 34885 31124 34897 31127
rect 34848 31096 34897 31124
rect 34848 31084 34854 31096
rect 34885 31093 34897 31096
rect 34931 31093 34943 31127
rect 34885 31087 34943 31093
rect 1104 31034 38272 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38272 31034
rect 1104 30960 38272 30982
rect 8018 30880 8024 30932
rect 8076 30880 8082 30932
rect 8938 30880 8944 30932
rect 8996 30880 9002 30932
rect 9674 30880 9680 30932
rect 9732 30920 9738 30932
rect 10045 30923 10103 30929
rect 10045 30920 10057 30923
rect 9732 30892 10057 30920
rect 9732 30880 9738 30892
rect 10045 30889 10057 30892
rect 10091 30889 10103 30923
rect 10045 30883 10103 30889
rect 12066 30880 12072 30932
rect 12124 30920 12130 30932
rect 15470 30920 15476 30932
rect 12124 30892 15476 30920
rect 12124 30880 12130 30892
rect 10597 30855 10655 30861
rect 6840 30824 9536 30852
rect 6840 30796 6868 30824
rect 6822 30744 6828 30796
rect 6880 30744 6886 30796
rect 9508 30793 9536 30824
rect 10597 30821 10609 30855
rect 10643 30821 10655 30855
rect 10597 30815 10655 30821
rect 9493 30787 9551 30793
rect 7484 30756 8708 30784
rect 7484 30725 7512 30756
rect 8680 30728 8708 30756
rect 9493 30753 9505 30787
rect 9539 30753 9551 30787
rect 9493 30747 9551 30753
rect 6457 30719 6515 30725
rect 6457 30685 6469 30719
rect 6503 30716 6515 30719
rect 7469 30719 7527 30725
rect 6503 30688 6684 30716
rect 6503 30685 6515 30688
rect 6457 30679 6515 30685
rect 6656 30592 6684 30688
rect 7469 30685 7481 30719
rect 7515 30685 7527 30719
rect 7469 30679 7527 30685
rect 7837 30719 7895 30725
rect 7837 30685 7849 30719
rect 7883 30716 7895 30719
rect 7883 30688 8156 30716
rect 7883 30685 7895 30688
rect 7837 30679 7895 30685
rect 7653 30651 7711 30657
rect 7653 30617 7665 30651
rect 7699 30617 7711 30651
rect 7653 30611 7711 30617
rect 7745 30651 7803 30657
rect 7745 30617 7757 30651
rect 7791 30648 7803 30651
rect 7926 30648 7932 30660
rect 7791 30620 7932 30648
rect 7791 30617 7803 30620
rect 7745 30611 7803 30617
rect 6362 30540 6368 30592
rect 6420 30580 6426 30592
rect 6549 30583 6607 30589
rect 6549 30580 6561 30583
rect 6420 30552 6561 30580
rect 6420 30540 6426 30552
rect 6549 30549 6561 30552
rect 6595 30549 6607 30583
rect 6549 30543 6607 30549
rect 6638 30540 6644 30592
rect 6696 30540 6702 30592
rect 7668 30580 7696 30611
rect 7926 30608 7932 30620
rect 7984 30608 7990 30660
rect 8128 30648 8156 30688
rect 8202 30676 8208 30728
rect 8260 30676 8266 30728
rect 8312 30688 8616 30716
rect 8312 30648 8340 30688
rect 8128 30620 8340 30648
rect 8478 30608 8484 30660
rect 8536 30608 8542 30660
rect 8588 30648 8616 30688
rect 8662 30676 8668 30728
rect 8720 30676 8726 30728
rect 8938 30676 8944 30728
rect 8996 30676 9002 30728
rect 9214 30676 9220 30728
rect 9272 30716 9278 30728
rect 9309 30719 9367 30725
rect 9309 30716 9321 30719
rect 9272 30688 9321 30716
rect 9272 30676 9278 30688
rect 9309 30685 9321 30688
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 10229 30719 10287 30725
rect 10229 30685 10241 30719
rect 10275 30716 10287 30719
rect 10612 30716 10640 30815
rect 10686 30744 10692 30796
rect 10744 30784 10750 30796
rect 11149 30787 11207 30793
rect 11149 30784 11161 30787
rect 10744 30756 11161 30784
rect 10744 30744 10750 30756
rect 11149 30753 11161 30756
rect 11195 30753 11207 30787
rect 11149 30747 11207 30753
rect 10275 30688 10640 30716
rect 12437 30719 12495 30725
rect 10275 30685 10287 30688
rect 10229 30679 10287 30685
rect 12437 30685 12449 30719
rect 12483 30716 12495 30719
rect 12483 30688 12517 30716
rect 12483 30685 12495 30688
rect 12437 30679 12495 30685
rect 8956 30648 8984 30676
rect 8588 30620 8984 30648
rect 10965 30651 11023 30657
rect 10965 30617 10977 30651
rect 11011 30648 11023 30651
rect 11238 30648 11244 30660
rect 11011 30620 11244 30648
rect 11011 30617 11023 30620
rect 10965 30611 11023 30617
rect 11238 30608 11244 30620
rect 11296 30648 11302 30660
rect 12452 30648 12480 30679
rect 12618 30676 12624 30728
rect 12676 30676 12682 30728
rect 12728 30725 12756 30892
rect 15470 30880 15476 30892
rect 15528 30880 15534 30932
rect 16485 30923 16543 30929
rect 16485 30889 16497 30923
rect 16531 30920 16543 30923
rect 16758 30920 16764 30932
rect 16531 30892 16764 30920
rect 16531 30889 16543 30892
rect 16485 30883 16543 30889
rect 16758 30880 16764 30892
rect 16816 30880 16822 30932
rect 16942 30880 16948 30932
rect 17000 30880 17006 30932
rect 18141 30923 18199 30929
rect 18141 30889 18153 30923
rect 18187 30920 18199 30923
rect 19245 30923 19303 30929
rect 19245 30920 19257 30923
rect 18187 30892 19257 30920
rect 18187 30889 18199 30892
rect 18141 30883 18199 30889
rect 19245 30889 19257 30892
rect 19291 30889 19303 30923
rect 19245 30883 19303 30889
rect 19886 30880 19892 30932
rect 19944 30920 19950 30932
rect 19944 30892 21864 30920
rect 19944 30880 19950 30892
rect 14826 30812 14832 30864
rect 14884 30852 14890 30864
rect 16960 30852 16988 30880
rect 14884 30824 16988 30852
rect 14884 30812 14890 30824
rect 14844 30784 14872 30812
rect 14752 30756 14872 30784
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30685 12771 30719
rect 12713 30679 12771 30685
rect 12805 30719 12863 30725
rect 12805 30685 12817 30719
rect 12851 30716 12863 30719
rect 13078 30716 13084 30728
rect 12851 30688 13084 30716
rect 12851 30685 12863 30688
rect 12805 30679 12863 30685
rect 13078 30676 13084 30688
rect 13136 30676 13142 30728
rect 14752 30648 14780 30756
rect 14918 30744 14924 30796
rect 14976 30744 14982 30796
rect 16574 30784 16580 30796
rect 15212 30756 16580 30784
rect 14829 30719 14887 30725
rect 14829 30685 14841 30719
rect 14875 30685 14887 30719
rect 14829 30679 14887 30685
rect 11296 30620 14780 30648
rect 14844 30648 14872 30679
rect 15010 30676 15016 30728
rect 15068 30676 15074 30728
rect 15102 30676 15108 30728
rect 15160 30676 15166 30728
rect 15120 30648 15148 30676
rect 14844 30620 15148 30648
rect 11296 30608 11302 30620
rect 8496 30580 8524 30608
rect 7668 30552 8524 30580
rect 8754 30540 8760 30592
rect 8812 30540 8818 30592
rect 9214 30540 9220 30592
rect 9272 30580 9278 30592
rect 9401 30583 9459 30589
rect 9401 30580 9413 30583
rect 9272 30552 9413 30580
rect 9272 30540 9278 30552
rect 9401 30549 9413 30552
rect 9447 30580 9459 30583
rect 11054 30580 11060 30592
rect 9447 30552 11060 30580
rect 9447 30549 9459 30552
rect 9401 30543 9459 30549
rect 11054 30540 11060 30552
rect 11112 30540 11118 30592
rect 12989 30583 13047 30589
rect 12989 30549 13001 30583
rect 13035 30580 13047 30583
rect 13630 30580 13636 30592
rect 13035 30552 13636 30580
rect 13035 30549 13047 30552
rect 12989 30543 13047 30549
rect 13630 30540 13636 30552
rect 13688 30540 13694 30592
rect 14550 30540 14556 30592
rect 14608 30540 14614 30592
rect 14918 30540 14924 30592
rect 14976 30580 14982 30592
rect 15212 30589 15240 30756
rect 16574 30744 16580 30756
rect 16632 30744 16638 30796
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30716 15347 30719
rect 15654 30716 15660 30728
rect 15335 30688 15660 30716
rect 15335 30685 15347 30688
rect 15289 30679 15347 30685
rect 15654 30676 15660 30688
rect 15712 30676 15718 30728
rect 16022 30676 16028 30728
rect 16080 30716 16086 30728
rect 16301 30719 16359 30725
rect 16301 30716 16313 30719
rect 16080 30688 16313 30716
rect 16080 30676 16086 30688
rect 16301 30685 16313 30688
rect 16347 30685 16359 30719
rect 16301 30679 16359 30685
rect 16669 30719 16727 30725
rect 16669 30685 16681 30719
rect 16715 30685 16727 30719
rect 16669 30679 16727 30685
rect 16762 30719 16820 30725
rect 16762 30685 16774 30719
rect 16808 30685 16820 30719
rect 16960 30716 16988 30824
rect 17034 30812 17040 30864
rect 17092 30812 17098 30864
rect 17218 30812 17224 30864
rect 17276 30852 17282 30864
rect 17586 30852 17592 30864
rect 17276 30824 17592 30852
rect 17276 30812 17282 30824
rect 17586 30812 17592 30824
rect 17644 30812 17650 30864
rect 17862 30812 17868 30864
rect 17920 30852 17926 30864
rect 18785 30855 18843 30861
rect 18785 30852 18797 30855
rect 17920 30824 18797 30852
rect 17920 30812 17926 30824
rect 18785 30821 18797 30824
rect 18831 30821 18843 30855
rect 18785 30815 18843 30821
rect 18966 30812 18972 30864
rect 19024 30812 19030 30864
rect 20806 30812 20812 30864
rect 20864 30812 20870 30864
rect 21174 30852 21180 30864
rect 21008 30824 21180 30852
rect 17052 30784 17080 30812
rect 17052 30756 17816 30784
rect 17218 30725 17224 30728
rect 17037 30719 17095 30725
rect 17037 30716 17049 30719
rect 16960 30688 17049 30716
rect 16762 30679 16820 30685
rect 17037 30685 17049 30688
rect 17083 30685 17095 30719
rect 17037 30679 17095 30685
rect 17175 30719 17224 30725
rect 17175 30685 17187 30719
rect 17221 30685 17224 30719
rect 17175 30679 17224 30685
rect 16117 30651 16175 30657
rect 16117 30617 16129 30651
rect 16163 30648 16175 30651
rect 16684 30648 16712 30679
rect 16163 30620 16712 30648
rect 16163 30617 16175 30620
rect 16117 30611 16175 30617
rect 15197 30583 15255 30589
rect 15197 30580 15209 30583
rect 14976 30552 15209 30580
rect 14976 30540 14982 30552
rect 15197 30549 15209 30552
rect 15243 30549 15255 30583
rect 15197 30543 15255 30549
rect 15470 30540 15476 30592
rect 15528 30580 15534 30592
rect 16574 30580 16580 30592
rect 15528 30552 16580 30580
rect 15528 30540 15534 30552
rect 16574 30540 16580 30552
rect 16632 30580 16638 30592
rect 16777 30580 16805 30679
rect 17218 30676 17224 30679
rect 17276 30676 17282 30728
rect 17589 30719 17647 30725
rect 17589 30685 17601 30719
rect 17635 30685 17647 30719
rect 17589 30679 17647 30685
rect 16942 30608 16948 30660
rect 17000 30608 17006 30660
rect 16632 30552 16805 30580
rect 16632 30540 16638 30552
rect 17310 30540 17316 30592
rect 17368 30540 17374 30592
rect 17604 30580 17632 30679
rect 17788 30657 17816 30756
rect 18248 30756 18920 30784
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30716 18015 30719
rect 18138 30716 18144 30728
rect 18003 30688 18144 30716
rect 18003 30685 18015 30688
rect 17957 30679 18015 30685
rect 18138 30676 18144 30688
rect 18196 30676 18202 30728
rect 18248 30725 18276 30756
rect 18233 30719 18291 30725
rect 18233 30685 18245 30719
rect 18279 30685 18291 30719
rect 18233 30679 18291 30685
rect 18601 30719 18659 30725
rect 18601 30685 18613 30719
rect 18647 30716 18659 30719
rect 18690 30716 18696 30728
rect 18647 30688 18696 30716
rect 18647 30685 18659 30688
rect 18601 30679 18659 30685
rect 17773 30651 17831 30657
rect 17773 30617 17785 30651
rect 17819 30617 17831 30651
rect 17773 30611 17831 30617
rect 17865 30651 17923 30657
rect 17865 30617 17877 30651
rect 17911 30648 17923 30651
rect 18248 30648 18276 30679
rect 18690 30676 18696 30688
rect 18748 30676 18754 30728
rect 17911 30620 18276 30648
rect 17911 30617 17923 30620
rect 17865 30611 17923 30617
rect 18322 30608 18328 30660
rect 18380 30648 18386 30660
rect 18417 30651 18475 30657
rect 18417 30648 18429 30651
rect 18380 30620 18429 30648
rect 18380 30608 18386 30620
rect 18417 30617 18429 30620
rect 18463 30617 18475 30651
rect 18417 30611 18475 30617
rect 18506 30608 18512 30660
rect 18564 30608 18570 30660
rect 18892 30648 18920 30756
rect 18984 30716 19012 30812
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 18984 30688 19257 30716
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19334 30676 19340 30728
rect 19392 30676 19398 30728
rect 20824 30716 20852 30812
rect 21008 30725 21036 30824
rect 21174 30812 21180 30824
rect 21232 30852 21238 30864
rect 21450 30852 21456 30864
rect 21232 30824 21456 30852
rect 21232 30812 21238 30824
rect 21450 30812 21456 30824
rect 21508 30812 21514 30864
rect 21726 30784 21732 30796
rect 21192 30756 21732 30784
rect 21192 30725 21220 30756
rect 21726 30744 21732 30756
rect 21784 30744 21790 30796
rect 21836 30784 21864 30892
rect 23198 30880 23204 30932
rect 23256 30880 23262 30932
rect 23474 30880 23480 30932
rect 23532 30920 23538 30932
rect 23934 30920 23940 30932
rect 23532 30892 23940 30920
rect 23532 30880 23538 30892
rect 23934 30880 23940 30892
rect 23992 30880 23998 30932
rect 27982 30880 27988 30932
rect 28040 30920 28046 30932
rect 28994 30920 29000 30932
rect 28040 30892 29000 30920
rect 28040 30880 28046 30892
rect 28994 30880 29000 30892
rect 29052 30920 29058 30932
rect 30190 30920 30196 30932
rect 29052 30892 30196 30920
rect 29052 30880 29058 30892
rect 30190 30880 30196 30892
rect 30248 30880 30254 30932
rect 34790 30880 34796 30932
rect 34848 30880 34854 30932
rect 23216 30852 23244 30880
rect 23845 30855 23903 30861
rect 23845 30852 23857 30855
rect 23216 30824 23857 30852
rect 23845 30821 23857 30824
rect 23891 30821 23903 30855
rect 23845 30815 23903 30821
rect 23952 30824 25268 30852
rect 23952 30784 23980 30824
rect 25240 30793 25268 30824
rect 25590 30812 25596 30864
rect 25648 30812 25654 30864
rect 28629 30855 28687 30861
rect 28629 30821 28641 30855
rect 28675 30852 28687 30855
rect 29270 30852 29276 30864
rect 28675 30824 29276 30852
rect 28675 30821 28687 30824
rect 28629 30815 28687 30821
rect 29270 30812 29276 30824
rect 29328 30812 29334 30864
rect 25225 30787 25283 30793
rect 21836 30756 22228 30784
rect 20901 30719 20959 30725
rect 20901 30716 20913 30719
rect 20824 30688 20913 30716
rect 20901 30685 20913 30688
rect 20947 30685 20959 30719
rect 20901 30679 20959 30685
rect 20993 30719 21051 30725
rect 20993 30685 21005 30719
rect 21039 30685 21051 30719
rect 20993 30679 21051 30685
rect 21177 30719 21235 30725
rect 21177 30685 21189 30719
rect 21223 30685 21235 30719
rect 21177 30679 21235 30685
rect 21266 30676 21272 30728
rect 21324 30676 21330 30728
rect 21358 30676 21364 30728
rect 21416 30676 21422 30728
rect 21450 30676 21456 30728
rect 21508 30676 21514 30728
rect 21545 30719 21603 30725
rect 21545 30685 21557 30719
rect 21591 30716 21603 30719
rect 21818 30716 21824 30728
rect 21591 30688 21824 30716
rect 21591 30685 21603 30688
rect 21545 30679 21603 30685
rect 21818 30676 21824 30688
rect 21876 30676 21882 30728
rect 21468 30648 21496 30676
rect 18892 30620 21496 30648
rect 21729 30651 21787 30657
rect 21729 30617 21741 30651
rect 21775 30648 21787 30651
rect 22200 30648 22228 30756
rect 22388 30756 23980 30784
rect 24044 30756 24900 30784
rect 22388 30728 22416 30756
rect 22370 30676 22376 30728
rect 22428 30676 22434 30728
rect 22830 30676 22836 30728
rect 22888 30716 22894 30728
rect 23109 30719 23167 30725
rect 23109 30716 23121 30719
rect 22888 30688 23121 30716
rect 22888 30676 22894 30688
rect 23109 30685 23121 30688
rect 23155 30685 23167 30719
rect 23109 30679 23167 30685
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30716 23443 30719
rect 23658 30716 23664 30728
rect 23431 30688 23664 30716
rect 23431 30685 23443 30688
rect 23385 30679 23443 30685
rect 23658 30676 23664 30688
rect 23716 30676 23722 30728
rect 23750 30676 23756 30728
rect 23808 30676 23814 30728
rect 23934 30676 23940 30728
rect 23992 30676 23998 30728
rect 24044 30725 24072 30756
rect 24029 30719 24087 30725
rect 24029 30685 24041 30719
rect 24075 30685 24087 30719
rect 24029 30679 24087 30685
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 23569 30651 23627 30657
rect 21775 30620 23428 30648
rect 21775 30617 21787 30620
rect 21729 30611 21787 30617
rect 18046 30580 18052 30592
rect 17604 30552 18052 30580
rect 18046 30540 18052 30552
rect 18104 30540 18110 30592
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 19613 30583 19671 30589
rect 19613 30580 19625 30583
rect 19392 30552 19625 30580
rect 19392 30540 19398 30552
rect 19613 30549 19625 30552
rect 19659 30549 19671 30583
rect 19613 30543 19671 30549
rect 20717 30583 20775 30589
rect 20717 30549 20729 30583
rect 20763 30580 20775 30583
rect 22370 30580 22376 30592
rect 20763 30552 22376 30580
rect 20763 30549 20775 30552
rect 20717 30543 20775 30549
rect 22370 30540 22376 30552
rect 22428 30540 22434 30592
rect 22922 30540 22928 30592
rect 22980 30540 22986 30592
rect 23290 30540 23296 30592
rect 23348 30540 23354 30592
rect 23400 30580 23428 30620
rect 23569 30617 23581 30651
rect 23615 30648 23627 30651
rect 24780 30648 24808 30679
rect 23615 30620 24808 30648
rect 24872 30648 24900 30756
rect 25225 30753 25237 30787
rect 25271 30753 25283 30787
rect 25608 30784 25636 30812
rect 25225 30747 25283 30753
rect 25409 30756 25636 30784
rect 25041 30719 25099 30725
rect 25041 30685 25053 30719
rect 25087 30716 25099 30719
rect 25314 30716 25320 30728
rect 25087 30688 25320 30716
rect 25087 30685 25099 30688
rect 25041 30679 25099 30685
rect 25314 30676 25320 30688
rect 25372 30676 25378 30728
rect 25409 30648 25437 30756
rect 25866 30744 25872 30796
rect 25924 30744 25930 30796
rect 34701 30787 34759 30793
rect 34701 30753 34713 30787
rect 34747 30784 34759 30787
rect 34808 30784 34836 30880
rect 34747 30756 34836 30784
rect 34747 30753 34759 30756
rect 34701 30747 34759 30753
rect 25590 30676 25596 30728
rect 25648 30676 25654 30728
rect 27062 30676 27068 30728
rect 27120 30676 27126 30728
rect 28810 30676 28816 30728
rect 28868 30676 28874 30728
rect 29178 30676 29184 30728
rect 29236 30676 29242 30728
rect 32769 30719 32827 30725
rect 32769 30685 32781 30719
rect 32815 30716 32827 30719
rect 32815 30688 33088 30716
rect 32815 30685 32827 30688
rect 32769 30679 32827 30685
rect 24872 30620 25437 30648
rect 23615 30617 23627 30620
rect 23569 30611 23627 30617
rect 28994 30608 29000 30660
rect 29052 30648 29058 30660
rect 30929 30651 30987 30657
rect 30929 30648 30941 30651
rect 29052 30620 30941 30648
rect 29052 30608 29058 30620
rect 30929 30617 30941 30620
rect 30975 30617 30987 30651
rect 30929 30611 30987 30617
rect 33060 30592 33088 30688
rect 34330 30676 34336 30728
rect 34388 30676 34394 30728
rect 34977 30651 35035 30657
rect 34977 30648 34989 30651
rect 34164 30620 34989 30648
rect 23658 30580 23664 30592
rect 23400 30552 23664 30580
rect 23658 30540 23664 30552
rect 23716 30540 23722 30592
rect 26970 30540 26976 30592
rect 27028 30580 27034 30592
rect 27157 30583 27215 30589
rect 27157 30580 27169 30583
rect 27028 30552 27169 30580
rect 27028 30540 27034 30552
rect 27157 30549 27169 30552
rect 27203 30549 27215 30583
rect 27157 30543 27215 30549
rect 29086 30540 29092 30592
rect 29144 30580 29150 30592
rect 29273 30583 29331 30589
rect 29273 30580 29285 30583
rect 29144 30552 29285 30580
rect 29144 30540 29150 30552
rect 29273 30549 29285 30552
rect 29319 30549 29331 30583
rect 29273 30543 29331 30549
rect 32214 30540 32220 30592
rect 32272 30540 32278 30592
rect 32490 30540 32496 30592
rect 32548 30580 32554 30592
rect 32861 30583 32919 30589
rect 32861 30580 32873 30583
rect 32548 30552 32873 30580
rect 32548 30540 32554 30552
rect 32861 30549 32873 30552
rect 32907 30549 32919 30583
rect 32861 30543 32919 30549
rect 33042 30540 33048 30592
rect 33100 30540 33106 30592
rect 34164 30589 34192 30620
rect 34977 30617 34989 30620
rect 35023 30617 35035 30651
rect 34977 30611 35035 30617
rect 35986 30608 35992 30660
rect 36044 30608 36050 30660
rect 36725 30651 36783 30657
rect 36725 30617 36737 30651
rect 36771 30617 36783 30651
rect 36725 30611 36783 30617
rect 34149 30583 34207 30589
rect 34149 30549 34161 30583
rect 34195 30549 34207 30583
rect 34149 30543 34207 30549
rect 34514 30540 34520 30592
rect 34572 30580 34578 30592
rect 36740 30580 36768 30611
rect 34572 30552 36768 30580
rect 34572 30540 34578 30552
rect 1104 30490 38272 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38272 30490
rect 1104 30416 38272 30438
rect 8754 30376 8760 30388
rect 8312 30348 8760 30376
rect 8018 30240 8024 30252
rect 7774 30212 8024 30240
rect 8018 30200 8024 30212
rect 8076 30200 8082 30252
rect 8312 30249 8340 30348
rect 8754 30336 8760 30348
rect 8812 30336 8818 30388
rect 9306 30336 9312 30388
rect 9364 30376 9370 30388
rect 14918 30376 14924 30388
rect 9364 30348 14924 30376
rect 9364 30336 9370 30348
rect 8478 30268 8484 30320
rect 8536 30308 8542 30320
rect 8536 30280 10548 30308
rect 8536 30268 8542 30280
rect 10520 30252 10548 30280
rect 10962 30268 10968 30320
rect 11020 30268 11026 30320
rect 8297 30243 8355 30249
rect 8297 30209 8309 30243
rect 8343 30209 8355 30243
rect 8297 30203 8355 30209
rect 8569 30243 8627 30249
rect 8569 30209 8581 30243
rect 8615 30209 8627 30243
rect 8569 30203 8627 30209
rect 8665 30243 8723 30249
rect 8665 30209 8677 30243
rect 8711 30238 8723 30243
rect 8938 30240 8944 30252
rect 8772 30238 8944 30240
rect 8711 30212 8944 30238
rect 8711 30210 8800 30212
rect 8711 30209 8723 30210
rect 8665 30203 8723 30209
rect 6362 30132 6368 30184
rect 6420 30132 6426 30184
rect 6641 30175 6699 30181
rect 6641 30141 6653 30175
rect 6687 30172 6699 30175
rect 8588 30172 8616 30203
rect 8938 30200 8944 30212
rect 8996 30200 9002 30252
rect 9214 30200 9220 30252
rect 9272 30200 9278 30252
rect 9950 30200 9956 30252
rect 10008 30240 10014 30252
rect 10045 30243 10103 30249
rect 10045 30240 10057 30243
rect 10008 30212 10057 30240
rect 10008 30200 10014 30212
rect 10045 30209 10057 30212
rect 10091 30240 10103 30243
rect 10091 30212 10364 30240
rect 10091 30209 10103 30212
rect 10045 30203 10103 30209
rect 9232 30172 9260 30200
rect 9766 30172 9772 30184
rect 6687 30144 7696 30172
rect 8588 30144 9260 30172
rect 9508 30144 9772 30172
rect 6687 30141 6699 30144
rect 6641 30135 6699 30141
rect 7668 30104 7696 30144
rect 8849 30107 8907 30113
rect 8849 30104 8861 30107
rect 7668 30076 8861 30104
rect 8849 30073 8861 30076
rect 8895 30073 8907 30107
rect 8849 30067 8907 30073
rect 8113 30039 8171 30045
rect 8113 30005 8125 30039
rect 8159 30036 8171 30039
rect 8202 30036 8208 30048
rect 8159 30008 8208 30036
rect 8159 30005 8171 30008
rect 8113 29999 8171 30005
rect 8202 29996 8208 30008
rect 8260 30036 8266 30048
rect 9508 30036 9536 30144
rect 9766 30132 9772 30144
rect 9824 30132 9830 30184
rect 10336 30104 10364 30212
rect 10502 30200 10508 30252
rect 10560 30200 10566 30252
rect 10980 30172 11008 30268
rect 11974 30200 11980 30252
rect 12032 30240 12038 30252
rect 12360 30249 12388 30348
rect 14918 30336 14924 30348
rect 14976 30336 14982 30388
rect 15010 30336 15016 30388
rect 15068 30336 15074 30388
rect 17310 30336 17316 30388
rect 17368 30376 17374 30388
rect 18414 30376 18420 30388
rect 17368 30348 18420 30376
rect 17368 30336 17374 30348
rect 18414 30336 18420 30348
rect 18472 30336 18478 30388
rect 18966 30336 18972 30388
rect 19024 30376 19030 30388
rect 19245 30379 19303 30385
rect 19245 30376 19257 30379
rect 19024 30348 19257 30376
rect 19024 30336 19030 30348
rect 19245 30345 19257 30348
rect 19291 30345 19303 30379
rect 19245 30339 19303 30345
rect 19996 30348 21220 30376
rect 12434 30268 12440 30320
rect 12492 30308 12498 30320
rect 12529 30311 12587 30317
rect 12529 30308 12541 30311
rect 12492 30280 12541 30308
rect 12492 30268 12498 30280
rect 12529 30277 12541 30280
rect 12575 30308 12587 30311
rect 12894 30308 12900 30320
rect 12575 30280 12900 30308
rect 12575 30277 12587 30280
rect 12529 30271 12587 30277
rect 12894 30268 12900 30280
rect 12952 30268 12958 30320
rect 12989 30311 13047 30317
rect 12989 30277 13001 30311
rect 13035 30308 13047 30311
rect 14734 30308 14740 30320
rect 13035 30280 14740 30308
rect 13035 30277 13047 30280
rect 12989 30271 13047 30277
rect 14734 30268 14740 30280
rect 14792 30268 14798 30320
rect 14826 30268 14832 30320
rect 14884 30268 14890 30320
rect 15028 30308 15056 30336
rect 15381 30311 15439 30317
rect 15381 30308 15393 30311
rect 15028 30280 15393 30308
rect 15381 30277 15393 30280
rect 15427 30277 15439 30311
rect 15381 30271 15439 30277
rect 16666 30268 16672 30320
rect 16724 30308 16730 30320
rect 16724 30280 17908 30308
rect 16724 30268 16730 30280
rect 17236 30252 17264 30280
rect 12253 30243 12311 30249
rect 12253 30240 12265 30243
rect 12032 30212 12265 30240
rect 12032 30200 12038 30212
rect 12253 30209 12265 30212
rect 12299 30209 12311 30243
rect 12253 30203 12311 30209
rect 12346 30243 12404 30249
rect 12346 30209 12358 30243
rect 12392 30209 12404 30243
rect 12346 30203 12404 30209
rect 12621 30243 12679 30249
rect 12621 30209 12633 30243
rect 12667 30209 12679 30243
rect 12621 30203 12679 30209
rect 12759 30243 12817 30249
rect 12759 30209 12771 30243
rect 12805 30240 12817 30243
rect 13446 30240 13452 30252
rect 12805 30212 13452 30240
rect 12805 30209 12817 30212
rect 12759 30203 12817 30209
rect 12636 30172 12664 30203
rect 13446 30200 13452 30212
rect 13504 30200 13510 30252
rect 14366 30200 14372 30252
rect 14424 30240 14430 30252
rect 15010 30240 15016 30252
rect 14424 30212 15016 30240
rect 14424 30200 14430 30212
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 15105 30243 15163 30249
rect 15105 30209 15117 30243
rect 15151 30209 15163 30243
rect 15105 30203 15163 30209
rect 15197 30243 15255 30249
rect 15197 30209 15209 30243
rect 15243 30240 15255 30243
rect 15286 30240 15292 30252
rect 15243 30212 15292 30240
rect 15243 30209 15255 30212
rect 15197 30203 15255 30209
rect 10980 30144 14688 30172
rect 10962 30104 10968 30116
rect 10336 30076 10968 30104
rect 10962 30064 10968 30076
rect 11020 30064 11026 30116
rect 13998 30064 14004 30116
rect 14056 30104 14062 30116
rect 14277 30107 14335 30113
rect 14277 30104 14289 30107
rect 14056 30076 14289 30104
rect 14056 30064 14062 30076
rect 14277 30073 14289 30076
rect 14323 30073 14335 30107
rect 14277 30067 14335 30073
rect 8260 30008 9536 30036
rect 10137 30039 10195 30045
rect 8260 29996 8266 30008
rect 10137 30005 10149 30039
rect 10183 30036 10195 30039
rect 10502 30036 10508 30048
rect 10183 30008 10508 30036
rect 10183 30005 10195 30008
rect 10137 29999 10195 30005
rect 10502 29996 10508 30008
rect 10560 29996 10566 30048
rect 12894 29996 12900 30048
rect 12952 29996 12958 30048
rect 14660 30036 14688 30144
rect 14734 30064 14740 30116
rect 14792 30104 14798 30116
rect 15120 30104 15148 30203
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 16942 30200 16948 30252
rect 17000 30200 17006 30252
rect 17038 30243 17096 30249
rect 17038 30209 17050 30243
rect 17084 30209 17096 30243
rect 17038 30203 17096 30209
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 17052 30172 17080 30203
rect 17218 30200 17224 30252
rect 17276 30200 17282 30252
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 17451 30243 17509 30249
rect 17451 30209 17463 30243
rect 17497 30240 17509 30243
rect 17678 30240 17684 30252
rect 17497 30212 17684 30240
rect 17497 30209 17509 30212
rect 17451 30203 17509 30209
rect 16632 30144 17080 30172
rect 16632 30132 16638 30144
rect 14792 30076 15148 30104
rect 14792 30064 14798 30076
rect 17328 30036 17356 30203
rect 17678 30200 17684 30212
rect 17736 30200 17742 30252
rect 17880 30172 17908 30280
rect 17954 30268 17960 30320
rect 18012 30268 18018 30320
rect 18782 30268 18788 30320
rect 18840 30308 18846 30320
rect 19996 30308 20024 30348
rect 18840 30280 20024 30308
rect 18840 30268 18846 30280
rect 20070 30268 20076 30320
rect 20128 30308 20134 30320
rect 20441 30311 20499 30317
rect 20441 30308 20453 30311
rect 20128 30280 20453 30308
rect 20128 30268 20134 30280
rect 20441 30277 20453 30280
rect 20487 30308 20499 30311
rect 20530 30308 20536 30320
rect 20487 30280 20536 30308
rect 20487 30277 20499 30280
rect 20441 30271 20499 30277
rect 20530 30268 20536 30280
rect 20588 30268 20594 30320
rect 20622 30268 20628 30320
rect 20680 30268 20686 30320
rect 20806 30268 20812 30320
rect 20864 30308 20870 30320
rect 21082 30308 21088 30320
rect 20864 30280 21088 30308
rect 20864 30268 20870 30280
rect 21082 30268 21088 30280
rect 21140 30268 21146 30320
rect 21192 30308 21220 30348
rect 21818 30336 21824 30388
rect 21876 30376 21882 30388
rect 22738 30376 22744 30388
rect 21876 30348 22744 30376
rect 21876 30336 21882 30348
rect 22738 30336 22744 30348
rect 22796 30336 22802 30388
rect 25038 30336 25044 30388
rect 25096 30376 25102 30388
rect 25682 30376 25688 30388
rect 25096 30348 25688 30376
rect 25096 30336 25102 30348
rect 25682 30336 25688 30348
rect 25740 30336 25746 30388
rect 26142 30336 26148 30388
rect 26200 30376 26206 30388
rect 26421 30379 26479 30385
rect 26421 30376 26433 30379
rect 26200 30348 26433 30376
rect 26200 30336 26206 30348
rect 26421 30345 26433 30348
rect 26467 30345 26479 30379
rect 26421 30339 26479 30345
rect 29196 30348 29500 30376
rect 21266 30308 21272 30320
rect 21192 30280 21272 30308
rect 21266 30268 21272 30280
rect 21324 30268 21330 30320
rect 21450 30268 21456 30320
rect 21508 30308 21514 30320
rect 25593 30311 25651 30317
rect 25593 30308 25605 30311
rect 21508 30280 25605 30308
rect 21508 30268 21514 30280
rect 25593 30277 25605 30280
rect 25639 30308 25651 30311
rect 26513 30311 26571 30317
rect 25639 30280 26464 30308
rect 25639 30277 25651 30280
rect 25593 30271 25651 30277
rect 18230 30200 18236 30252
rect 18288 30240 18294 30252
rect 18288 30212 19380 30240
rect 18288 30200 18294 30212
rect 18782 30172 18788 30184
rect 17880 30144 18788 30172
rect 18782 30132 18788 30144
rect 18840 30132 18846 30184
rect 19352 30172 19380 30212
rect 19886 30200 19892 30252
rect 19944 30240 19950 30252
rect 19981 30243 20039 30249
rect 19981 30240 19993 30243
rect 19944 30212 19993 30240
rect 19944 30200 19950 30212
rect 19981 30209 19993 30212
rect 20027 30209 20039 30243
rect 19981 30203 20039 30209
rect 20162 30200 20168 30252
rect 20220 30200 20226 30252
rect 20254 30200 20260 30252
rect 20312 30200 20318 30252
rect 20714 30200 20720 30252
rect 20772 30240 20778 30252
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 20772 30212 23397 30240
rect 20772 30200 20778 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 25317 30243 25375 30249
rect 25317 30209 25329 30243
rect 25363 30209 25375 30243
rect 25317 30203 25375 30209
rect 25332 30172 25360 30203
rect 25498 30200 25504 30252
rect 25556 30200 25562 30252
rect 25682 30200 25688 30252
rect 25740 30240 25746 30252
rect 26050 30240 26056 30252
rect 25740 30212 26056 30240
rect 25740 30200 25746 30212
rect 26050 30200 26056 30212
rect 26108 30200 26114 30252
rect 26326 30172 26332 30184
rect 19352 30144 26332 30172
rect 26326 30132 26332 30144
rect 26384 30132 26390 30184
rect 17589 30107 17647 30113
rect 17589 30073 17601 30107
rect 17635 30104 17647 30107
rect 19150 30104 19156 30116
rect 17635 30076 19156 30104
rect 17635 30073 17647 30076
rect 17589 30067 17647 30073
rect 19150 30064 19156 30076
rect 19208 30064 19214 30116
rect 19702 30064 19708 30116
rect 19760 30104 19766 30116
rect 20809 30107 20867 30113
rect 20809 30104 20821 30107
rect 19760 30076 20821 30104
rect 19760 30064 19766 30076
rect 20809 30073 20821 30076
rect 20855 30104 20867 30107
rect 20855 30076 21772 30104
rect 20855 30073 20867 30076
rect 20809 30067 20867 30073
rect 17954 30036 17960 30048
rect 14660 30008 17960 30036
rect 17954 29996 17960 30008
rect 18012 30036 18018 30048
rect 18506 30036 18512 30048
rect 18012 30008 18512 30036
rect 18012 29996 18018 30008
rect 18506 29996 18512 30008
rect 18564 29996 18570 30048
rect 19794 29996 19800 30048
rect 19852 29996 19858 30048
rect 20346 29996 20352 30048
rect 20404 30036 20410 30048
rect 20625 30039 20683 30045
rect 20625 30036 20637 30039
rect 20404 30008 20637 30036
rect 20404 29996 20410 30008
rect 20625 30005 20637 30008
rect 20671 30005 20683 30039
rect 20625 29999 20683 30005
rect 21266 29996 21272 30048
rect 21324 29996 21330 30048
rect 21453 30039 21511 30045
rect 21453 30005 21465 30039
rect 21499 30036 21511 30039
rect 21634 30036 21640 30048
rect 21499 30008 21640 30036
rect 21499 30005 21511 30008
rect 21453 29999 21511 30005
rect 21634 29996 21640 30008
rect 21692 29996 21698 30048
rect 21744 30036 21772 30076
rect 22646 30064 22652 30116
rect 22704 30064 22710 30116
rect 23198 30064 23204 30116
rect 23256 30104 23262 30116
rect 24302 30104 24308 30116
rect 23256 30076 24308 30104
rect 23256 30064 23262 30076
rect 24302 30064 24308 30076
rect 24360 30064 24366 30116
rect 24670 30064 24676 30116
rect 24728 30064 24734 30116
rect 22664 30036 22692 30064
rect 21744 30008 22692 30036
rect 22922 29996 22928 30048
rect 22980 30036 22986 30048
rect 23106 30036 23112 30048
rect 22980 30008 23112 30036
rect 22980 29996 22986 30008
rect 23106 29996 23112 30008
rect 23164 29996 23170 30048
rect 25866 29996 25872 30048
rect 25924 29996 25930 30048
rect 26050 29996 26056 30048
rect 26108 29996 26114 30048
rect 26436 30036 26464 30280
rect 26513 30277 26525 30311
rect 26559 30308 26571 30311
rect 27154 30308 27160 30320
rect 26559 30280 27160 30308
rect 26559 30277 26571 30280
rect 26513 30271 26571 30277
rect 27154 30268 27160 30280
rect 27212 30268 27218 30320
rect 28534 30308 28540 30320
rect 28474 30280 28540 30308
rect 28534 30268 28540 30280
rect 28592 30308 28598 30320
rect 29196 30308 29224 30348
rect 28592 30280 29224 30308
rect 28592 30268 28598 30280
rect 29270 30268 29276 30320
rect 29328 30308 29334 30320
rect 29365 30311 29423 30317
rect 29365 30308 29377 30311
rect 29328 30280 29377 30308
rect 29328 30268 29334 30280
rect 29365 30277 29377 30280
rect 29411 30277 29423 30311
rect 29472 30308 29500 30348
rect 32490 30336 32496 30388
rect 32548 30336 32554 30388
rect 34057 30379 34115 30385
rect 34057 30345 34069 30379
rect 34103 30376 34115 30379
rect 34330 30376 34336 30388
rect 34103 30348 34336 30376
rect 34103 30345 34115 30348
rect 34057 30339 34115 30345
rect 34330 30336 34336 30348
rect 34388 30336 34394 30388
rect 29472 30280 29854 30308
rect 29365 30271 29423 30277
rect 30834 30268 30840 30320
rect 30892 30308 30898 30320
rect 32508 30308 32536 30336
rect 30892 30280 31524 30308
rect 30892 30268 30898 30280
rect 30742 30200 30748 30252
rect 30800 30240 30806 30252
rect 31496 30249 31524 30280
rect 32140 30280 32536 30308
rect 32140 30249 32168 30280
rect 33134 30268 33140 30320
rect 33192 30268 33198 30320
rect 34425 30311 34483 30317
rect 34425 30277 34437 30311
rect 34471 30308 34483 30311
rect 34514 30308 34520 30320
rect 34471 30280 34520 30308
rect 34471 30277 34483 30280
rect 34425 30271 34483 30277
rect 34514 30268 34520 30280
rect 34572 30268 34578 30320
rect 31205 30243 31263 30249
rect 31205 30240 31217 30243
rect 30800 30212 31217 30240
rect 30800 30200 30806 30212
rect 31205 30209 31217 30212
rect 31251 30209 31263 30243
rect 31205 30203 31263 30209
rect 31389 30243 31447 30249
rect 31389 30209 31401 30243
rect 31435 30209 31447 30243
rect 31389 30203 31447 30209
rect 31481 30243 31539 30249
rect 31481 30209 31493 30243
rect 31527 30209 31539 30243
rect 31481 30203 31539 30209
rect 32125 30243 32183 30249
rect 32125 30209 32137 30243
rect 32171 30209 32183 30243
rect 32125 30203 32183 30209
rect 26694 30132 26700 30184
rect 26752 30172 26758 30184
rect 26878 30172 26884 30184
rect 26752 30144 26884 30172
rect 26752 30132 26758 30144
rect 26878 30132 26884 30144
rect 26936 30132 26942 30184
rect 26970 30132 26976 30184
rect 27028 30132 27034 30184
rect 27246 30132 27252 30184
rect 27304 30132 27310 30184
rect 27890 30132 27896 30184
rect 27948 30172 27954 30184
rect 28997 30175 29055 30181
rect 28997 30172 29009 30175
rect 27948 30144 29009 30172
rect 27948 30132 27954 30144
rect 28997 30141 29009 30144
rect 29043 30141 29055 30175
rect 28997 30135 29055 30141
rect 29086 30132 29092 30184
rect 29144 30132 29150 30184
rect 31404 30172 31432 30203
rect 29196 30144 31432 30172
rect 29196 30036 29224 30144
rect 26436 30008 29224 30036
rect 29822 29996 29828 30048
rect 29880 30036 29886 30048
rect 30837 30039 30895 30045
rect 30837 30036 30849 30039
rect 29880 30008 30849 30036
rect 29880 29996 29886 30008
rect 30837 30005 30849 30008
rect 30883 30005 30895 30039
rect 30837 29999 30895 30005
rect 31018 29996 31024 30048
rect 31076 29996 31082 30048
rect 31404 30036 31432 30144
rect 32398 30132 32404 30184
rect 32456 30132 32462 30184
rect 33778 30132 33784 30184
rect 33836 30132 33842 30184
rect 34238 30132 34244 30184
rect 34296 30172 34302 30184
rect 34517 30175 34575 30181
rect 34517 30172 34529 30175
rect 34296 30144 34529 30172
rect 34296 30132 34302 30144
rect 34517 30141 34529 30144
rect 34563 30141 34575 30175
rect 34517 30135 34575 30141
rect 34609 30175 34667 30181
rect 34609 30141 34621 30175
rect 34655 30141 34667 30175
rect 34609 30135 34667 30141
rect 33796 30104 33824 30132
rect 34624 30104 34652 30135
rect 33796 30076 34652 30104
rect 31662 30036 31668 30048
rect 31404 30008 31668 30036
rect 31662 29996 31668 30008
rect 31720 30036 31726 30048
rect 33873 30039 33931 30045
rect 33873 30036 33885 30039
rect 31720 30008 33885 30036
rect 31720 29996 31726 30008
rect 33873 30005 33885 30008
rect 33919 30005 33931 30039
rect 33873 29999 33931 30005
rect 1104 29946 38272 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38272 29946
rect 1104 29872 38272 29894
rect 12526 29792 12532 29844
rect 12584 29792 12590 29844
rect 12894 29792 12900 29844
rect 12952 29792 12958 29844
rect 16853 29835 16911 29841
rect 16853 29801 16865 29835
rect 16899 29832 16911 29835
rect 16942 29832 16948 29844
rect 16899 29804 16948 29832
rect 16899 29801 16911 29804
rect 16853 29795 16911 29801
rect 16942 29792 16948 29804
rect 17000 29792 17006 29844
rect 17494 29792 17500 29844
rect 17552 29832 17558 29844
rect 19702 29832 19708 29844
rect 17552 29804 19708 29832
rect 17552 29792 17558 29804
rect 19702 29792 19708 29804
rect 19760 29792 19766 29844
rect 20070 29792 20076 29844
rect 20128 29792 20134 29844
rect 20162 29792 20168 29844
rect 20220 29832 20226 29844
rect 20257 29835 20315 29841
rect 20257 29832 20269 29835
rect 20220 29804 20269 29832
rect 20220 29792 20226 29804
rect 20257 29801 20269 29804
rect 20303 29801 20315 29835
rect 20257 29795 20315 29801
rect 20346 29792 20352 29844
rect 20404 29832 20410 29844
rect 20625 29835 20683 29841
rect 20625 29832 20637 29835
rect 20404 29804 20637 29832
rect 20404 29792 20410 29804
rect 20625 29801 20637 29804
rect 20671 29801 20683 29835
rect 20625 29795 20683 29801
rect 20714 29792 20720 29844
rect 20772 29832 20778 29844
rect 23937 29835 23995 29841
rect 23937 29832 23949 29835
rect 20772 29804 23949 29832
rect 20772 29792 20778 29804
rect 23937 29801 23949 29804
rect 23983 29832 23995 29835
rect 25222 29832 25228 29844
rect 23983 29804 25228 29832
rect 23983 29801 23995 29804
rect 23937 29795 23995 29801
rect 25222 29792 25228 29804
rect 25280 29792 25286 29844
rect 25774 29792 25780 29844
rect 25832 29792 25838 29844
rect 25866 29792 25872 29844
rect 25924 29792 25930 29844
rect 26050 29792 26056 29844
rect 26108 29792 26114 29844
rect 26326 29792 26332 29844
rect 26384 29792 26390 29844
rect 26421 29835 26479 29841
rect 26421 29801 26433 29835
rect 26467 29832 26479 29835
rect 27246 29832 27252 29844
rect 26467 29804 27252 29832
rect 26467 29801 26479 29804
rect 26421 29795 26479 29801
rect 27246 29792 27252 29804
rect 27304 29792 27310 29844
rect 28353 29835 28411 29841
rect 28353 29801 28365 29835
rect 28399 29832 28411 29835
rect 28810 29832 28816 29844
rect 28399 29804 28816 29832
rect 28399 29801 28411 29804
rect 28353 29795 28411 29801
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 30377 29835 30435 29841
rect 30377 29801 30389 29835
rect 30423 29832 30435 29835
rect 30742 29832 30748 29844
rect 30423 29804 30748 29832
rect 30423 29801 30435 29804
rect 30377 29795 30435 29801
rect 30742 29792 30748 29804
rect 30800 29792 30806 29844
rect 34514 29832 34520 29844
rect 31726 29804 34520 29832
rect 8018 29724 8024 29776
rect 8076 29764 8082 29776
rect 9122 29764 9128 29776
rect 8076 29736 9128 29764
rect 8076 29724 8082 29736
rect 9122 29724 9128 29736
rect 9180 29724 9186 29776
rect 4448 29668 6684 29696
rect 4448 29637 4476 29668
rect 6656 29640 6684 29668
rect 4433 29631 4491 29637
rect 4433 29597 4445 29631
rect 4479 29597 4491 29631
rect 4433 29591 4491 29597
rect 5718 29588 5724 29640
rect 5776 29588 5782 29640
rect 6638 29588 6644 29640
rect 6696 29628 6702 29640
rect 7561 29631 7619 29637
rect 7561 29628 7573 29631
rect 6696 29600 7573 29628
rect 6696 29588 6702 29600
rect 7561 29597 7573 29600
rect 7607 29597 7619 29631
rect 7561 29591 7619 29597
rect 6270 29520 6276 29572
rect 6328 29560 6334 29572
rect 8036 29560 8064 29724
rect 9585 29631 9643 29637
rect 9585 29628 9597 29631
rect 6328 29532 8064 29560
rect 8496 29600 9597 29628
rect 6328 29520 6334 29532
rect 8496 29504 8524 29600
rect 9585 29597 9597 29600
rect 9631 29597 9643 29631
rect 9585 29591 9643 29597
rect 12253 29631 12311 29637
rect 12253 29597 12265 29631
rect 12299 29597 12311 29631
rect 12253 29591 12311 29597
rect 9122 29520 9128 29572
rect 9180 29560 9186 29572
rect 10318 29560 10324 29572
rect 9180 29532 10324 29560
rect 9180 29520 9186 29532
rect 10318 29520 10324 29532
rect 10376 29520 10382 29572
rect 12268 29560 12296 29591
rect 12342 29588 12348 29640
rect 12400 29588 12406 29640
rect 12912 29628 12940 29792
rect 14921 29767 14979 29773
rect 14921 29733 14933 29767
rect 14967 29764 14979 29767
rect 16209 29767 16267 29773
rect 16209 29764 16221 29767
rect 14967 29736 16221 29764
rect 14967 29733 14979 29736
rect 14921 29727 14979 29733
rect 16209 29733 16221 29736
rect 16255 29733 16267 29767
rect 21818 29764 21824 29776
rect 16209 29727 16267 29733
rect 16500 29736 21824 29764
rect 13817 29699 13875 29705
rect 13817 29665 13829 29699
rect 13863 29696 13875 29699
rect 14645 29699 14703 29705
rect 14645 29696 14657 29699
rect 13863 29668 14657 29696
rect 13863 29665 13875 29668
rect 13817 29659 13875 29665
rect 14645 29665 14657 29668
rect 14691 29665 14703 29699
rect 14645 29659 14703 29665
rect 15013 29699 15071 29705
rect 15013 29665 15025 29699
rect 15059 29696 15071 29699
rect 15562 29696 15568 29708
rect 15059 29668 15568 29696
rect 15059 29665 15071 29668
rect 15013 29659 15071 29665
rect 15562 29656 15568 29668
rect 15620 29656 15626 29708
rect 15672 29668 16252 29696
rect 13541 29631 13599 29637
rect 13541 29628 13553 29631
rect 12912 29600 13553 29628
rect 13541 29597 13553 29600
rect 13587 29597 13599 29631
rect 13541 29591 13599 29597
rect 13630 29588 13636 29640
rect 13688 29588 13694 29640
rect 13906 29588 13912 29640
rect 13964 29588 13970 29640
rect 14550 29588 14556 29640
rect 14608 29628 14614 29640
rect 14829 29631 14887 29637
rect 14829 29628 14841 29631
rect 14608 29600 14841 29628
rect 14608 29588 14614 29600
rect 14829 29597 14841 29600
rect 14875 29597 14887 29631
rect 14829 29591 14887 29597
rect 15105 29631 15163 29637
rect 15105 29597 15117 29631
rect 15151 29597 15163 29631
rect 15105 29591 15163 29597
rect 15120 29560 15148 29591
rect 15286 29588 15292 29640
rect 15344 29588 15350 29640
rect 15672 29637 15700 29668
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29597 15715 29631
rect 15657 29591 15715 29597
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 15841 29631 15899 29637
rect 15841 29628 15853 29631
rect 15804 29600 15853 29628
rect 15804 29588 15810 29600
rect 15841 29597 15853 29600
rect 15887 29597 15899 29631
rect 15841 29591 15899 29597
rect 15933 29631 15991 29637
rect 15933 29597 15945 29631
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29628 16083 29631
rect 16114 29628 16120 29640
rect 16071 29600 16120 29628
rect 16071 29597 16083 29600
rect 16025 29591 16083 29597
rect 15562 29560 15568 29572
rect 12268 29532 15568 29560
rect 15562 29520 15568 29532
rect 15620 29520 15626 29572
rect 4522 29452 4528 29504
rect 4580 29452 4586 29504
rect 7650 29452 7656 29504
rect 7708 29452 7714 29504
rect 8478 29452 8484 29504
rect 8536 29452 8542 29504
rect 9674 29452 9680 29504
rect 9732 29452 9738 29504
rect 11974 29452 11980 29504
rect 12032 29492 12038 29504
rect 12894 29492 12900 29504
rect 12032 29464 12900 29492
rect 12032 29452 12038 29464
rect 12894 29452 12900 29464
rect 12952 29452 12958 29504
rect 13354 29452 13360 29504
rect 13412 29452 13418 29504
rect 15856 29492 15884 29591
rect 15948 29560 15976 29591
rect 16114 29588 16120 29600
rect 16172 29588 16178 29640
rect 16224 29628 16252 29668
rect 16301 29631 16359 29637
rect 16301 29628 16313 29631
rect 16224 29600 16313 29628
rect 16301 29597 16313 29600
rect 16347 29628 16359 29631
rect 16500 29628 16528 29736
rect 21818 29724 21824 29736
rect 21876 29724 21882 29776
rect 22002 29724 22008 29776
rect 22060 29724 22066 29776
rect 23290 29724 23296 29776
rect 23348 29764 23354 29776
rect 24121 29767 24179 29773
rect 24121 29764 24133 29767
rect 23348 29736 24133 29764
rect 23348 29724 23354 29736
rect 24121 29733 24133 29736
rect 24167 29733 24179 29767
rect 25792 29764 25820 29792
rect 24121 29727 24179 29733
rect 25516 29736 25820 29764
rect 18506 29656 18512 29708
rect 18564 29656 18570 29708
rect 18782 29656 18788 29708
rect 18840 29696 18846 29708
rect 19610 29696 19616 29708
rect 18840 29668 19616 29696
rect 18840 29656 18846 29668
rect 19610 29656 19616 29668
rect 19668 29656 19674 29708
rect 20162 29696 20168 29708
rect 20088 29668 20168 29696
rect 16347 29600 16528 29628
rect 16347 29597 16359 29600
rect 16301 29591 16359 29597
rect 16574 29588 16580 29640
rect 16632 29628 16638 29640
rect 16669 29631 16727 29637
rect 16669 29628 16681 29631
rect 16632 29600 16681 29628
rect 16632 29588 16638 29600
rect 16669 29597 16681 29600
rect 16715 29628 16727 29631
rect 17126 29628 17132 29640
rect 16715 29600 17132 29628
rect 16715 29597 16727 29600
rect 16669 29591 16727 29597
rect 17126 29588 17132 29600
rect 17184 29588 17190 29640
rect 17954 29588 17960 29640
rect 18012 29628 18018 29640
rect 18187 29631 18245 29637
rect 18187 29628 18199 29631
rect 18012 29600 18199 29628
rect 18012 29588 18018 29600
rect 18187 29597 18199 29600
rect 18233 29597 18245 29631
rect 18187 29591 18245 29597
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29597 18383 29631
rect 18325 29591 18383 29597
rect 18417 29631 18475 29637
rect 18417 29597 18429 29631
rect 18463 29628 18475 29631
rect 18524 29628 18552 29656
rect 18463 29600 18552 29628
rect 18601 29631 18659 29637
rect 18463 29597 18475 29600
rect 18417 29591 18475 29597
rect 18601 29597 18613 29631
rect 18647 29628 18659 29631
rect 19150 29628 19156 29640
rect 18647 29600 19156 29628
rect 18647 29597 18659 29600
rect 18601 29591 18659 29597
rect 16206 29560 16212 29572
rect 15948 29532 16212 29560
rect 16206 29520 16212 29532
rect 16264 29520 16270 29572
rect 18340 29560 18368 29591
rect 19150 29588 19156 29600
rect 19208 29588 19214 29640
rect 19889 29631 19947 29637
rect 19889 29597 19901 29631
rect 19935 29628 19947 29631
rect 19978 29628 19984 29640
rect 19935 29600 19984 29628
rect 19935 29597 19947 29600
rect 19889 29591 19947 29597
rect 19242 29560 19248 29572
rect 18248 29532 19248 29560
rect 18248 29504 18276 29532
rect 19242 29520 19248 29532
rect 19300 29560 19306 29572
rect 19904 29560 19932 29591
rect 19978 29588 19984 29600
rect 20036 29588 20042 29640
rect 20088 29637 20116 29668
rect 20162 29656 20168 29668
rect 20220 29656 20226 29708
rect 20806 29696 20812 29708
rect 20640 29668 20812 29696
rect 20073 29631 20131 29637
rect 20073 29597 20085 29631
rect 20119 29597 20131 29631
rect 20073 29591 20131 29597
rect 20254 29588 20260 29640
rect 20312 29628 20318 29640
rect 20640 29628 20668 29668
rect 20806 29656 20812 29668
rect 20864 29656 20870 29708
rect 20312 29600 20668 29628
rect 22020 29628 22048 29724
rect 24210 29656 24216 29708
rect 24268 29656 24274 29708
rect 22281 29631 22339 29637
rect 22281 29628 22293 29631
rect 22020 29600 22293 29628
rect 20312 29588 20318 29600
rect 19300 29532 19932 29560
rect 20441 29563 20499 29569
rect 19300 29520 19306 29532
rect 20441 29529 20453 29563
rect 20487 29560 20499 29563
rect 20530 29560 20536 29572
rect 20487 29532 20536 29560
rect 20487 29529 20499 29532
rect 20441 29523 20499 29529
rect 20530 29520 20536 29532
rect 20588 29520 20594 29572
rect 20640 29569 20668 29600
rect 22281 29597 22293 29600
rect 22327 29597 22339 29631
rect 22649 29631 22707 29637
rect 22281 29591 22339 29597
rect 22388 29600 22600 29628
rect 20625 29563 20683 29569
rect 20625 29529 20637 29563
rect 20671 29529 20683 29563
rect 20625 29523 20683 29529
rect 22002 29520 22008 29572
rect 22060 29560 22066 29572
rect 22388 29560 22416 29600
rect 22060 29532 22416 29560
rect 22060 29520 22066 29532
rect 22462 29520 22468 29572
rect 22520 29520 22526 29572
rect 22572 29569 22600 29600
rect 22649 29597 22661 29631
rect 22695 29628 22707 29631
rect 22922 29628 22928 29640
rect 22695 29600 22928 29628
rect 22695 29597 22707 29600
rect 22649 29591 22707 29597
rect 22922 29588 22928 29600
rect 22980 29588 22986 29640
rect 23106 29588 23112 29640
rect 23164 29628 23170 29640
rect 23753 29631 23811 29637
rect 23753 29628 23765 29631
rect 23164 29600 23765 29628
rect 23164 29588 23170 29600
rect 23753 29597 23765 29600
rect 23799 29628 23811 29631
rect 23842 29628 23848 29640
rect 23799 29600 23848 29628
rect 23799 29597 23811 29600
rect 23753 29591 23811 29597
rect 23842 29588 23848 29600
rect 23900 29588 23906 29640
rect 23937 29631 23995 29637
rect 23937 29597 23949 29631
rect 23983 29628 23995 29631
rect 24228 29628 24256 29656
rect 23983 29600 24256 29628
rect 23983 29597 23995 29600
rect 23937 29591 23995 29597
rect 25406 29588 25412 29640
rect 25464 29588 25470 29640
rect 25516 29637 25544 29736
rect 25884 29696 25912 29792
rect 25792 29668 25912 29696
rect 25792 29637 25820 29668
rect 25501 29631 25559 29637
rect 25501 29597 25513 29631
rect 25547 29597 25559 29631
rect 25501 29591 25559 29597
rect 25593 29631 25651 29637
rect 25593 29597 25605 29631
rect 25639 29597 25651 29631
rect 25593 29591 25651 29597
rect 25777 29631 25835 29637
rect 25777 29597 25789 29631
rect 25823 29597 25835 29631
rect 25777 29591 25835 29597
rect 25869 29631 25927 29637
rect 25869 29597 25881 29631
rect 25915 29597 25927 29631
rect 26068 29628 26096 29792
rect 26344 29764 26372 29792
rect 31726 29764 31754 29804
rect 34514 29792 34520 29804
rect 34572 29792 34578 29844
rect 26344 29736 31754 29764
rect 33781 29767 33839 29773
rect 26510 29656 26516 29708
rect 26568 29696 26574 29708
rect 28813 29699 28871 29705
rect 28813 29696 28825 29699
rect 26568 29668 28825 29696
rect 26568 29656 26574 29668
rect 28813 29665 28825 29668
rect 28859 29665 28871 29699
rect 28813 29659 28871 29665
rect 26605 29631 26663 29637
rect 26605 29628 26617 29631
rect 26068 29600 26617 29628
rect 25869 29591 25927 29597
rect 26605 29597 26617 29600
rect 26651 29597 26663 29631
rect 26605 29591 26663 29597
rect 22557 29563 22615 29569
rect 22557 29529 22569 29563
rect 22603 29529 22615 29563
rect 25424 29560 25452 29588
rect 25608 29560 25636 29591
rect 25884 29560 25912 29591
rect 26510 29560 26516 29572
rect 22557 29523 22615 29529
rect 22664 29532 23704 29560
rect 25424 29532 25636 29560
rect 25792 29532 26516 29560
rect 15930 29492 15936 29504
rect 15856 29464 15936 29492
rect 15930 29452 15936 29464
rect 15988 29452 15994 29504
rect 16390 29452 16396 29504
rect 16448 29492 16454 29504
rect 16485 29495 16543 29501
rect 16485 29492 16497 29495
rect 16448 29464 16497 29492
rect 16448 29452 16454 29464
rect 16485 29461 16497 29464
rect 16531 29461 16543 29495
rect 16485 29455 16543 29461
rect 16577 29495 16635 29501
rect 16577 29461 16589 29495
rect 16623 29492 16635 29495
rect 16666 29492 16672 29504
rect 16623 29464 16672 29492
rect 16623 29461 16635 29464
rect 16577 29455 16635 29461
rect 16666 29452 16672 29464
rect 16724 29492 16730 29504
rect 17402 29492 17408 29504
rect 16724 29464 17408 29492
rect 16724 29452 16730 29464
rect 17402 29452 17408 29464
rect 17460 29452 17466 29504
rect 17954 29452 17960 29504
rect 18012 29452 18018 29504
rect 18230 29452 18236 29504
rect 18288 29452 18294 29504
rect 18506 29452 18512 29504
rect 18564 29492 18570 29504
rect 19334 29492 19340 29504
rect 18564 29464 19340 29492
rect 18564 29452 18570 29464
rect 19334 29452 19340 29464
rect 19392 29452 19398 29504
rect 19610 29452 19616 29504
rect 19668 29492 19674 29504
rect 20809 29495 20867 29501
rect 20809 29492 20821 29495
rect 19668 29464 20821 29492
rect 19668 29452 19674 29464
rect 20809 29461 20821 29464
rect 20855 29492 20867 29495
rect 21174 29492 21180 29504
rect 20855 29464 21180 29492
rect 20855 29461 20867 29464
rect 20809 29455 20867 29461
rect 21174 29452 21180 29464
rect 21232 29492 21238 29504
rect 22664 29492 22692 29532
rect 23676 29504 23704 29532
rect 25792 29504 25820 29532
rect 26510 29520 26516 29532
rect 26568 29520 26574 29572
rect 28828 29560 28856 29659
rect 28902 29656 28908 29708
rect 28960 29656 28966 29708
rect 30098 29656 30104 29708
rect 30156 29656 30162 29708
rect 29454 29588 29460 29640
rect 29512 29628 29518 29640
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 29512 29600 29745 29628
rect 29512 29588 29518 29600
rect 29733 29597 29745 29600
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29822 29588 29828 29640
rect 29880 29588 29886 29640
rect 30116 29628 30144 29656
rect 30198 29631 30256 29637
rect 30198 29628 30210 29631
rect 30116 29600 30210 29628
rect 30198 29597 30210 29600
rect 30244 29597 30256 29631
rect 30198 29591 30256 29597
rect 29840 29560 29868 29588
rect 28828 29532 29868 29560
rect 30006 29520 30012 29572
rect 30064 29520 30070 29572
rect 30101 29563 30159 29569
rect 30101 29529 30113 29563
rect 30147 29560 30159 29563
rect 30300 29560 30328 29736
rect 33781 29733 33793 29767
rect 33827 29764 33839 29767
rect 33827 29736 35204 29764
rect 33827 29733 33839 29736
rect 33781 29727 33839 29733
rect 31018 29696 31024 29708
rect 30484 29668 31024 29696
rect 30484 29637 30512 29668
rect 31018 29656 31024 29668
rect 31076 29656 31082 29708
rect 31128 29668 33088 29696
rect 30469 29631 30527 29637
rect 30469 29597 30481 29631
rect 30515 29597 30527 29631
rect 30469 29591 30527 29597
rect 30650 29588 30656 29640
rect 30708 29588 30714 29640
rect 30745 29631 30803 29637
rect 30745 29597 30757 29631
rect 30791 29597 30803 29631
rect 30745 29591 30803 29597
rect 30871 29625 30929 29631
rect 31128 29628 31156 29668
rect 30871 29591 30883 29625
rect 30917 29622 30929 29625
rect 31036 29622 31156 29628
rect 30917 29600 31156 29622
rect 31205 29631 31263 29637
rect 30917 29594 31064 29600
rect 30917 29591 30929 29594
rect 30147 29532 30328 29560
rect 30147 29529 30159 29532
rect 30101 29523 30159 29529
rect 30374 29520 30380 29572
rect 30432 29560 30438 29572
rect 30760 29560 30788 29591
rect 30871 29585 30929 29591
rect 30432 29532 30788 29560
rect 30432 29520 30438 29532
rect 21232 29464 22692 29492
rect 21232 29452 21238 29464
rect 22830 29452 22836 29504
rect 22888 29452 22894 29504
rect 23658 29452 23664 29504
rect 23716 29452 23722 29504
rect 25317 29495 25375 29501
rect 25317 29461 25329 29495
rect 25363 29492 25375 29495
rect 25498 29492 25504 29504
rect 25363 29464 25504 29492
rect 25363 29461 25375 29464
rect 25317 29455 25375 29461
rect 25498 29452 25504 29464
rect 25556 29452 25562 29504
rect 25774 29452 25780 29504
rect 25832 29452 25838 29504
rect 27982 29452 27988 29504
rect 28040 29492 28046 29504
rect 28721 29495 28779 29501
rect 28721 29492 28733 29495
rect 28040 29464 28733 29492
rect 28040 29452 28046 29464
rect 28721 29461 28733 29464
rect 28767 29461 28779 29495
rect 28721 29455 28779 29461
rect 28902 29452 28908 29504
rect 28960 29492 28966 29504
rect 31036 29492 31064 29594
rect 31205 29597 31217 29631
rect 31251 29628 31263 29631
rect 31754 29628 31760 29640
rect 31251 29600 31760 29628
rect 31251 29597 31263 29600
rect 31205 29591 31263 29597
rect 31754 29588 31760 29600
rect 31812 29628 31818 29640
rect 32214 29628 32220 29640
rect 31812 29600 32220 29628
rect 31812 29588 31818 29600
rect 32214 29588 32220 29600
rect 32272 29588 32278 29640
rect 31113 29563 31171 29569
rect 31113 29529 31125 29563
rect 31159 29560 31171 29563
rect 32858 29560 32864 29572
rect 31159 29532 32864 29560
rect 31159 29529 31171 29532
rect 31113 29523 31171 29529
rect 32858 29520 32864 29532
rect 32916 29520 32922 29572
rect 32950 29520 32956 29572
rect 33008 29520 33014 29572
rect 33060 29560 33088 29668
rect 34330 29656 34336 29708
rect 34388 29656 34394 29708
rect 34698 29588 34704 29640
rect 34756 29588 34762 29640
rect 35176 29637 35204 29736
rect 35161 29631 35219 29637
rect 35161 29597 35173 29631
rect 35207 29597 35219 29631
rect 35161 29591 35219 29597
rect 34149 29563 34207 29569
rect 34149 29560 34161 29563
rect 33060 29532 34161 29560
rect 34149 29529 34161 29532
rect 34195 29560 34207 29563
rect 34195 29532 36400 29560
rect 34195 29529 34207 29532
rect 34149 29523 34207 29529
rect 36372 29504 36400 29532
rect 28960 29464 31064 29492
rect 28960 29452 28966 29464
rect 32490 29452 32496 29504
rect 32548 29492 32554 29504
rect 34238 29492 34244 29504
rect 32548 29464 34244 29492
rect 32548 29452 32554 29464
rect 34238 29452 34244 29464
rect 34296 29452 34302 29504
rect 34790 29452 34796 29504
rect 34848 29452 34854 29504
rect 34974 29452 34980 29504
rect 35032 29452 35038 29504
rect 36354 29452 36360 29504
rect 36412 29452 36418 29504
rect 1104 29402 38272 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38272 29402
rect 1104 29328 38272 29350
rect 4522 29248 4528 29300
rect 4580 29248 4586 29300
rect 6825 29291 6883 29297
rect 6825 29288 6837 29291
rect 6196 29260 6837 29288
rect 4540 29220 4568 29248
rect 6196 29229 6224 29260
rect 6825 29257 6837 29260
rect 6871 29288 6883 29291
rect 16298 29288 16304 29300
rect 6871 29260 16304 29288
rect 6871 29257 6883 29260
rect 6825 29251 6883 29257
rect 16298 29248 16304 29260
rect 16356 29248 16362 29300
rect 17954 29248 17960 29300
rect 18012 29288 18018 29300
rect 18782 29288 18788 29300
rect 18012 29260 18644 29288
rect 18012 29248 18018 29260
rect 4172 29192 4568 29220
rect 6181 29223 6239 29229
rect 4172 29161 4200 29192
rect 6181 29189 6193 29223
rect 6227 29189 6239 29223
rect 7650 29220 7656 29232
rect 6181 29183 6239 29189
rect 7484 29192 7656 29220
rect 4157 29155 4215 29161
rect 4157 29121 4169 29155
rect 4203 29121 4215 29155
rect 6270 29152 6276 29164
rect 5566 29124 6276 29152
rect 4157 29115 4215 29121
rect 6270 29112 6276 29124
rect 6328 29112 6334 29164
rect 6730 29112 6736 29164
rect 6788 29112 6794 29164
rect 7484 29161 7512 29192
rect 7650 29180 7656 29192
rect 7708 29180 7714 29232
rect 9122 29220 9128 29232
rect 8970 29192 9128 29220
rect 9122 29180 9128 29192
rect 9180 29180 9186 29232
rect 9674 29220 9680 29232
rect 9508 29192 9680 29220
rect 9508 29161 9536 29192
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 10318 29180 10324 29232
rect 10376 29180 10382 29232
rect 12250 29180 12256 29232
rect 12308 29220 12314 29232
rect 13998 29220 14004 29232
rect 12308 29192 14004 29220
rect 12308 29180 12314 29192
rect 13998 29180 14004 29192
rect 14056 29180 14062 29232
rect 16206 29220 16212 29232
rect 14108 29192 16212 29220
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29121 7527 29155
rect 7469 29115 7527 29121
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29121 9551 29155
rect 12342 29152 12348 29164
rect 9493 29115 9551 29121
rect 11900 29124 12348 29152
rect 11900 29096 11928 29124
rect 12342 29112 12348 29124
rect 12400 29152 12406 29164
rect 12437 29155 12495 29161
rect 12437 29152 12449 29155
rect 12400 29124 12449 29152
rect 12400 29112 12406 29124
rect 12437 29121 12449 29124
rect 12483 29152 12495 29155
rect 13173 29155 13231 29161
rect 13173 29152 13185 29155
rect 12483 29124 13185 29152
rect 12483 29121 12495 29124
rect 12437 29115 12495 29121
rect 13173 29121 13185 29124
rect 13219 29121 13231 29155
rect 13173 29115 13231 29121
rect 6638 29044 6644 29096
rect 6696 29084 6702 29096
rect 7009 29087 7067 29093
rect 7009 29084 7021 29087
rect 6696 29056 7021 29084
rect 6696 29044 6702 29056
rect 7009 29053 7021 29056
rect 7055 29084 7067 29087
rect 7374 29084 7380 29096
rect 7055 29056 7380 29084
rect 7055 29053 7067 29056
rect 7009 29047 7067 29053
rect 7374 29044 7380 29056
rect 7432 29044 7438 29096
rect 7742 29044 7748 29096
rect 7800 29044 7806 29096
rect 7834 29044 7840 29096
rect 7892 29084 7898 29096
rect 11241 29087 11299 29093
rect 7892 29056 10824 29084
rect 7892 29044 7898 29056
rect 10796 29016 10824 29056
rect 11241 29053 11253 29087
rect 11287 29084 11299 29087
rect 11514 29084 11520 29096
rect 11287 29056 11520 29084
rect 11287 29053 11299 29056
rect 11241 29047 11299 29053
rect 11514 29044 11520 29056
rect 11572 29044 11578 29096
rect 11882 29044 11888 29096
rect 11940 29044 11946 29096
rect 12066 29044 12072 29096
rect 12124 29084 12130 29096
rect 12253 29087 12311 29093
rect 12253 29084 12265 29087
rect 12124 29056 12265 29084
rect 12124 29044 12130 29056
rect 12253 29053 12265 29056
rect 12299 29053 12311 29087
rect 12253 29047 12311 29053
rect 12989 29087 13047 29093
rect 12989 29053 13001 29087
rect 13035 29084 13047 29087
rect 14108 29084 14136 29192
rect 16206 29180 16212 29192
rect 16264 29180 16270 29232
rect 18417 29223 18475 29229
rect 18417 29220 18429 29223
rect 18064 29192 18429 29220
rect 14182 29112 14188 29164
rect 14240 29152 14246 29164
rect 14918 29152 14924 29164
rect 14240 29124 14924 29152
rect 14240 29112 14246 29124
rect 14918 29112 14924 29124
rect 14976 29152 14982 29164
rect 14976 29124 17908 29152
rect 14976 29112 14982 29124
rect 13035 29056 14136 29084
rect 17880 29084 17908 29124
rect 18064 29084 18092 29192
rect 18417 29189 18429 29192
rect 18463 29189 18475 29223
rect 18417 29183 18475 29189
rect 18234 29155 18292 29161
rect 18234 29121 18246 29155
rect 18280 29121 18292 29155
rect 18234 29115 18292 29121
rect 18327 29155 18385 29161
rect 18506 29155 18512 29164
rect 18327 29121 18339 29155
rect 18373 29150 18385 29155
rect 18432 29150 18512 29155
rect 18373 29127 18512 29150
rect 18373 29122 18460 29127
rect 18373 29121 18385 29122
rect 18327 29115 18385 29121
rect 17880 29056 18092 29084
rect 13035 29053 13047 29056
rect 12989 29047 13047 29053
rect 12621 29019 12679 29025
rect 12621 29016 12633 29019
rect 10796 28988 12633 29016
rect 12621 28985 12633 28988
rect 12667 28985 12679 29019
rect 12621 28979 12679 28985
rect 13354 28976 13360 29028
rect 13412 28976 13418 29028
rect 16206 28976 16212 29028
rect 16264 29016 16270 29028
rect 16666 29016 16672 29028
rect 16264 28988 16672 29016
rect 16264 28976 16270 28988
rect 16666 28976 16672 28988
rect 16724 28976 16730 29028
rect 18046 28976 18052 29028
rect 18104 28976 18110 29028
rect 18248 29016 18276 29115
rect 18506 29112 18512 29127
rect 18564 29112 18570 29164
rect 18616 29161 18644 29260
rect 18708 29260 18788 29288
rect 18708 29161 18736 29260
rect 18782 29248 18788 29260
rect 18840 29248 18846 29300
rect 19058 29248 19064 29300
rect 19116 29288 19122 29300
rect 21910 29288 21916 29300
rect 19116 29260 21916 29288
rect 19116 29248 19122 29260
rect 21910 29248 21916 29260
rect 21968 29248 21974 29300
rect 22002 29248 22008 29300
rect 22060 29248 22066 29300
rect 22189 29291 22247 29297
rect 22189 29257 22201 29291
rect 22235 29288 22247 29291
rect 22462 29288 22468 29300
rect 22235 29260 22468 29288
rect 22235 29257 22247 29260
rect 22189 29251 22247 29257
rect 22462 29248 22468 29260
rect 22520 29248 22526 29300
rect 22554 29248 22560 29300
rect 22612 29248 22618 29300
rect 22830 29248 22836 29300
rect 22888 29248 22894 29300
rect 23842 29248 23848 29300
rect 23900 29288 23906 29300
rect 25406 29288 25412 29300
rect 23900 29260 25412 29288
rect 23900 29248 23906 29260
rect 25406 29248 25412 29260
rect 25464 29248 25470 29300
rect 28718 29288 28724 29300
rect 25516 29260 28724 29288
rect 19242 29220 19248 29232
rect 18897 29192 19248 29220
rect 18808 29161 18866 29167
rect 18601 29155 18659 29161
rect 18601 29121 18613 29155
rect 18647 29121 18659 29155
rect 18601 29115 18659 29121
rect 18693 29155 18751 29161
rect 18693 29121 18705 29155
rect 18739 29121 18751 29155
rect 18808 29127 18820 29161
rect 18854 29158 18866 29161
rect 18897 29158 18925 29192
rect 19242 29180 19248 29192
rect 19300 29180 19306 29232
rect 22020 29220 22048 29248
rect 22572 29220 22600 29248
rect 22020 29192 22416 29220
rect 22388 29164 22416 29192
rect 22480 29192 22600 29220
rect 22480 29164 22508 29192
rect 18854 29130 18925 29158
rect 18854 29127 18866 29130
rect 18808 29121 18866 29127
rect 18693 29115 18751 29121
rect 20714 29112 20720 29164
rect 20772 29152 20778 29164
rect 21542 29152 21548 29164
rect 20772 29124 21548 29152
rect 20772 29112 20778 29124
rect 21542 29112 21548 29124
rect 21600 29152 21606 29164
rect 21821 29155 21879 29161
rect 21821 29152 21833 29155
rect 21600 29124 21833 29152
rect 21600 29112 21606 29124
rect 21821 29121 21833 29124
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 22002 29112 22008 29164
rect 22060 29112 22066 29164
rect 22278 29112 22284 29164
rect 22336 29112 22342 29164
rect 22370 29112 22376 29164
rect 22428 29112 22434 29164
rect 22462 29112 22468 29164
rect 22520 29112 22526 29164
rect 22554 29112 22560 29164
rect 22612 29112 22618 29164
rect 22646 29112 22652 29164
rect 22704 29112 22710 29164
rect 22848 29152 22876 29248
rect 25516 29220 25544 29260
rect 24044 29192 25544 29220
rect 25608 29192 26004 29220
rect 24044 29164 24072 29192
rect 23201 29155 23259 29161
rect 23201 29152 23213 29155
rect 22848 29124 23213 29152
rect 23201 29121 23213 29124
rect 23247 29121 23259 29155
rect 23201 29115 23259 29121
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29152 23535 29155
rect 23566 29152 23572 29164
rect 23523 29124 23572 29152
rect 23523 29121 23535 29124
rect 23477 29115 23535 29121
rect 23566 29112 23572 29124
rect 23624 29112 23630 29164
rect 23658 29112 23664 29164
rect 23716 29112 23722 29164
rect 24026 29112 24032 29164
rect 24084 29112 24090 29164
rect 25317 29155 25375 29161
rect 25317 29121 25329 29155
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 18877 29087 18935 29093
rect 18877 29053 18889 29087
rect 18923 29084 18935 29087
rect 19058 29084 19064 29096
rect 18923 29056 19064 29084
rect 18923 29053 18935 29056
rect 18877 29047 18935 29053
rect 19058 29044 19064 29056
rect 19116 29084 19122 29096
rect 25332 29084 25360 29115
rect 25406 29112 25412 29164
rect 25464 29112 25470 29164
rect 25498 29112 25504 29164
rect 25556 29112 25562 29164
rect 25608 29084 25636 29192
rect 25685 29155 25743 29161
rect 25685 29121 25697 29155
rect 25731 29152 25743 29155
rect 25731 29124 25912 29152
rect 25731 29121 25743 29124
rect 25685 29115 25743 29121
rect 19116 29056 25636 29084
rect 19116 29044 19122 29056
rect 19153 29019 19211 29025
rect 19153 29016 19165 29019
rect 18248 28988 19165 29016
rect 19153 28985 19165 28988
rect 19199 28985 19211 29019
rect 19153 28979 19211 28985
rect 21266 28976 21272 29028
rect 21324 29016 21330 29028
rect 22094 29016 22100 29028
rect 21324 28988 22100 29016
rect 21324 28976 21330 28988
rect 22094 28976 22100 28988
rect 22152 28976 22158 29028
rect 22833 29019 22891 29025
rect 22833 28985 22845 29019
rect 22879 29016 22891 29019
rect 23293 29019 23351 29025
rect 23293 29016 23305 29019
rect 22879 28988 23305 29016
rect 22879 28985 22891 28988
rect 22833 28979 22891 28985
rect 23293 28985 23305 28988
rect 23339 28985 23351 29019
rect 23293 28979 23351 28985
rect 23385 29019 23443 29025
rect 23385 28985 23397 29019
rect 23431 29016 23443 29019
rect 24210 29016 24216 29028
rect 23431 28988 24216 29016
rect 23431 28985 23443 28988
rect 23385 28979 23443 28985
rect 24210 28976 24216 28988
rect 24268 28976 24274 29028
rect 25041 29019 25099 29025
rect 25041 28985 25053 29019
rect 25087 29016 25099 29019
rect 25222 29016 25228 29028
rect 25087 28988 25228 29016
rect 25087 28985 25099 28988
rect 25041 28979 25099 28985
rect 25222 28976 25228 28988
rect 25280 28976 25286 29028
rect 25314 28976 25320 29028
rect 25372 29016 25378 29028
rect 25884 29016 25912 29124
rect 25976 29084 26004 29192
rect 26988 29161 27016 29260
rect 26973 29155 27031 29161
rect 26973 29121 26985 29155
rect 27019 29121 27031 29155
rect 28552 29152 28580 29260
rect 28718 29248 28724 29260
rect 28776 29248 28782 29300
rect 29914 29248 29920 29300
rect 29972 29248 29978 29300
rect 30374 29248 30380 29300
rect 30432 29288 30438 29300
rect 31018 29288 31024 29300
rect 30432 29260 31024 29288
rect 30432 29248 30438 29260
rect 31018 29248 31024 29260
rect 31076 29288 31082 29300
rect 31294 29288 31300 29300
rect 31076 29260 31300 29288
rect 31076 29248 31082 29260
rect 31294 29248 31300 29260
rect 31352 29248 31358 29300
rect 31662 29248 31668 29300
rect 31720 29288 31726 29300
rect 32585 29291 32643 29297
rect 32585 29288 32597 29291
rect 31720 29260 32597 29288
rect 31720 29248 31726 29260
rect 32585 29257 32597 29260
rect 32631 29257 32643 29291
rect 32585 29251 32643 29257
rect 32950 29248 32956 29300
rect 33008 29288 33014 29300
rect 34698 29288 34704 29300
rect 33008 29260 34704 29288
rect 33008 29248 33014 29260
rect 34698 29248 34704 29260
rect 34756 29248 34762 29300
rect 34790 29248 34796 29300
rect 34848 29248 34854 29300
rect 28629 29223 28687 29229
rect 28629 29189 28641 29223
rect 28675 29220 28687 29223
rect 31754 29220 31760 29232
rect 28675 29192 31760 29220
rect 28675 29189 28687 29192
rect 28629 29183 28687 29189
rect 31754 29180 31760 29192
rect 31812 29180 31818 29232
rect 31938 29180 31944 29232
rect 31996 29220 32002 29232
rect 32490 29220 32496 29232
rect 31996 29192 32496 29220
rect 31996 29180 32002 29192
rect 32490 29180 32496 29192
rect 32548 29180 32554 29232
rect 34808 29220 34836 29248
rect 34348 29192 34836 29220
rect 31570 29152 31576 29164
rect 28552 29124 31576 29152
rect 26973 29115 27031 29121
rect 31570 29112 31576 29124
rect 31628 29112 31634 29164
rect 34348 29161 34376 29192
rect 34882 29180 34888 29232
rect 34940 29220 34946 29232
rect 34940 29192 35098 29220
rect 34940 29180 34946 29192
rect 36354 29180 36360 29232
rect 36412 29180 36418 29232
rect 34333 29155 34391 29161
rect 34333 29121 34345 29155
rect 34379 29121 34391 29155
rect 34333 29115 34391 29121
rect 36630 29112 36636 29164
rect 36688 29112 36694 29164
rect 36814 29112 36820 29164
rect 36872 29112 36878 29164
rect 28902 29084 28908 29096
rect 25976 29056 28908 29084
rect 28902 29044 28908 29056
rect 28960 29044 28966 29096
rect 32306 29044 32312 29096
rect 32364 29044 32370 29096
rect 32766 29044 32772 29096
rect 32824 29084 32830 29096
rect 33410 29084 33416 29096
rect 32824 29056 33416 29084
rect 32824 29044 32830 29056
rect 33410 29044 33416 29056
rect 33468 29044 33474 29096
rect 34609 29087 34667 29093
rect 34609 29053 34621 29087
rect 34655 29084 34667 29087
rect 34974 29084 34980 29096
rect 34655 29056 34980 29084
rect 34655 29053 34667 29056
rect 34609 29047 34667 29053
rect 34974 29044 34980 29056
rect 35032 29044 35038 29096
rect 25372 28988 25912 29016
rect 25372 28976 25378 28988
rect 4420 28951 4478 28957
rect 4420 28917 4432 28951
rect 4466 28948 4478 28951
rect 4982 28948 4988 28960
rect 4466 28920 4988 28948
rect 4466 28917 4478 28920
rect 4420 28911 4478 28917
rect 4982 28908 4988 28920
rect 5040 28908 5046 28960
rect 6362 28908 6368 28960
rect 6420 28908 6426 28960
rect 9122 28908 9128 28960
rect 9180 28948 9186 28960
rect 9217 28951 9275 28957
rect 9217 28948 9229 28951
rect 9180 28920 9229 28948
rect 9180 28908 9186 28920
rect 9217 28917 9229 28920
rect 9263 28917 9275 28951
rect 9217 28911 9275 28917
rect 9756 28951 9814 28957
rect 9756 28917 9768 28951
rect 9802 28948 9814 28951
rect 10226 28948 10232 28960
rect 9802 28920 10232 28948
rect 9802 28917 9814 28920
rect 9756 28911 9814 28917
rect 10226 28908 10232 28920
rect 10284 28908 10290 28960
rect 10410 28908 10416 28960
rect 10468 28948 10474 28960
rect 12161 28951 12219 28957
rect 12161 28948 12173 28951
rect 10468 28920 12173 28948
rect 10468 28908 10474 28920
rect 12161 28917 12173 28920
rect 12207 28917 12219 28951
rect 12161 28911 12219 28917
rect 13078 28908 13084 28960
rect 13136 28948 13142 28960
rect 13630 28948 13636 28960
rect 13136 28920 13636 28948
rect 13136 28908 13142 28920
rect 13630 28908 13636 28920
rect 13688 28908 13694 28960
rect 16022 28908 16028 28960
rect 16080 28948 16086 28960
rect 17218 28948 17224 28960
rect 16080 28920 17224 28948
rect 16080 28908 16086 28920
rect 17218 28908 17224 28920
rect 17276 28908 17282 28960
rect 18506 28908 18512 28960
rect 18564 28948 18570 28960
rect 18785 28951 18843 28957
rect 18785 28948 18797 28951
rect 18564 28920 18797 28948
rect 18564 28908 18570 28920
rect 18785 28917 18797 28920
rect 18831 28948 18843 28951
rect 20070 28948 20076 28960
rect 18831 28920 20076 28948
rect 18831 28917 18843 28920
rect 18785 28911 18843 28917
rect 20070 28908 20076 28920
rect 20128 28908 20134 28960
rect 20622 28908 20628 28960
rect 20680 28948 20686 28960
rect 22646 28948 22652 28960
rect 20680 28920 22652 28948
rect 20680 28908 20686 28920
rect 22646 28908 22652 28920
rect 22704 28908 22710 28960
rect 22925 28951 22983 28957
rect 22925 28917 22937 28951
rect 22971 28948 22983 28951
rect 23474 28948 23480 28960
rect 22971 28920 23480 28948
rect 22971 28917 22983 28920
rect 22925 28911 22983 28917
rect 23474 28908 23480 28920
rect 23532 28908 23538 28960
rect 25884 28948 25912 28988
rect 27982 28976 27988 29028
rect 28040 29016 28046 29028
rect 31938 29016 31944 29028
rect 28040 28988 31944 29016
rect 28040 28976 28046 28988
rect 31938 28976 31944 28988
rect 31996 28976 32002 29028
rect 32125 29019 32183 29025
rect 32125 28985 32137 29019
rect 32171 29016 32183 29019
rect 32324 29016 32352 29044
rect 32171 28988 32352 29016
rect 37001 29019 37059 29025
rect 32171 28985 32183 28988
rect 32125 28979 32183 28985
rect 37001 28985 37013 29019
rect 37047 29016 37059 29019
rect 37274 29016 37280 29028
rect 37047 28988 37280 29016
rect 37047 28985 37059 28988
rect 37001 28979 37059 28985
rect 37274 28976 37280 28988
rect 37332 28976 37338 29028
rect 26694 28948 26700 28960
rect 25884 28920 26700 28948
rect 26694 28908 26700 28920
rect 26752 28908 26758 28960
rect 27062 28908 27068 28960
rect 27120 28908 27126 28960
rect 28994 28908 29000 28960
rect 29052 28948 29058 28960
rect 29546 28948 29552 28960
rect 29052 28920 29552 28948
rect 29052 28908 29058 28920
rect 29546 28908 29552 28920
rect 29604 28908 29610 28960
rect 31478 28908 31484 28960
rect 31536 28948 31542 28960
rect 31665 28951 31723 28957
rect 31665 28948 31677 28951
rect 31536 28920 31677 28948
rect 31536 28908 31542 28920
rect 31665 28917 31677 28920
rect 31711 28917 31723 28951
rect 31665 28911 31723 28917
rect 1104 28858 38272 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38272 28858
rect 1104 28784 38272 28806
rect 4982 28704 4988 28756
rect 5040 28704 5046 28756
rect 7742 28704 7748 28756
rect 7800 28744 7806 28756
rect 8757 28747 8815 28753
rect 8757 28744 8769 28747
rect 7800 28716 8769 28744
rect 7800 28704 7806 28716
rect 8757 28713 8769 28716
rect 8803 28713 8815 28747
rect 8757 28707 8815 28713
rect 10226 28704 10232 28756
rect 10284 28744 10290 28756
rect 10689 28747 10747 28753
rect 10689 28744 10701 28747
rect 10284 28716 10701 28744
rect 10284 28704 10290 28716
rect 10689 28713 10701 28716
rect 10735 28713 10747 28747
rect 10689 28707 10747 28713
rect 12434 28704 12440 28756
rect 12492 28744 12498 28756
rect 13078 28744 13084 28756
rect 12492 28716 13084 28744
rect 12492 28704 12498 28716
rect 13078 28704 13084 28716
rect 13136 28744 13142 28756
rect 15562 28744 15568 28756
rect 13136 28716 15568 28744
rect 13136 28704 13142 28716
rect 15562 28704 15568 28716
rect 15620 28744 15626 28756
rect 20714 28744 20720 28756
rect 15620 28716 20720 28744
rect 15620 28704 15626 28716
rect 20714 28704 20720 28716
rect 20772 28704 20778 28756
rect 33686 28744 33692 28756
rect 22066 28716 33692 28744
rect 7834 28676 7840 28688
rect 1964 28648 7840 28676
rect 1964 28549 1992 28648
rect 7834 28636 7840 28648
rect 7892 28636 7898 28688
rect 8386 28636 8392 28688
rect 8444 28676 8450 28688
rect 10502 28676 10508 28688
rect 8444 28648 10508 28676
rect 8444 28636 8450 28648
rect 10502 28636 10508 28648
rect 10560 28636 10566 28688
rect 11146 28636 11152 28688
rect 11204 28636 11210 28688
rect 19426 28636 19432 28688
rect 19484 28676 19490 28688
rect 22066 28676 22094 28716
rect 33686 28704 33692 28716
rect 33744 28704 33750 28756
rect 19484 28648 22094 28676
rect 22848 28648 23793 28676
rect 19484 28636 19490 28648
rect 6362 28608 6368 28620
rect 5184 28580 6368 28608
rect 5184 28549 5212 28580
rect 6362 28568 6368 28580
rect 6420 28568 6426 28620
rect 8018 28608 8024 28620
rect 6840 28580 8024 28608
rect 1949 28543 2007 28549
rect 1949 28509 1961 28543
rect 1995 28509 2007 28543
rect 1949 28503 2007 28509
rect 4249 28543 4307 28549
rect 4249 28509 4261 28543
rect 4295 28509 4307 28543
rect 4249 28503 4307 28509
rect 5169 28543 5227 28549
rect 5169 28509 5181 28543
rect 5215 28509 5227 28543
rect 5169 28503 5227 28509
rect 4264 28472 4292 28503
rect 5350 28500 5356 28552
rect 5408 28500 5414 28552
rect 6840 28549 6868 28580
rect 8018 28568 8024 28580
rect 8076 28608 8082 28620
rect 11164 28608 11192 28636
rect 13725 28611 13783 28617
rect 8076 28580 11652 28608
rect 8076 28568 8082 28580
rect 6825 28543 6883 28549
rect 6825 28509 6837 28543
rect 6871 28509 6883 28543
rect 6825 28503 6883 28509
rect 8205 28543 8263 28549
rect 8205 28509 8217 28543
rect 8251 28509 8263 28543
rect 8205 28503 8263 28509
rect 5368 28472 5396 28500
rect 4264 28444 5396 28472
rect 1762 28364 1768 28416
rect 1820 28364 1826 28416
rect 4338 28364 4344 28416
rect 4396 28364 4402 28416
rect 6914 28364 6920 28416
rect 6972 28364 6978 28416
rect 8220 28404 8248 28503
rect 8386 28500 8392 28552
rect 8444 28500 8450 28552
rect 8573 28543 8631 28549
rect 8573 28509 8585 28543
rect 8619 28540 8631 28543
rect 8938 28540 8944 28552
rect 8619 28512 8944 28540
rect 8619 28509 8631 28512
rect 8573 28503 8631 28509
rect 8938 28500 8944 28512
rect 8996 28500 9002 28552
rect 9122 28500 9128 28552
rect 9180 28500 9186 28552
rect 10137 28543 10195 28549
rect 10137 28509 10149 28543
rect 10183 28509 10195 28543
rect 10137 28503 10195 28509
rect 8481 28475 8539 28481
rect 8481 28441 8493 28475
rect 8527 28472 8539 28475
rect 8846 28472 8852 28484
rect 8527 28444 8852 28472
rect 8527 28441 8539 28444
rect 8481 28435 8539 28441
rect 8846 28432 8852 28444
rect 8904 28432 8910 28484
rect 9677 28407 9735 28413
rect 9677 28404 9689 28407
rect 8220 28376 9689 28404
rect 9677 28373 9689 28376
rect 9723 28373 9735 28407
rect 10152 28404 10180 28503
rect 10410 28500 10416 28552
rect 10468 28500 10474 28552
rect 10502 28500 10508 28552
rect 10560 28500 10566 28552
rect 10870 28500 10876 28552
rect 10928 28500 10934 28552
rect 10962 28500 10968 28552
rect 11020 28500 11026 28552
rect 11149 28543 11207 28549
rect 11149 28509 11161 28543
rect 11195 28509 11207 28543
rect 11149 28503 11207 28509
rect 11241 28543 11299 28549
rect 11241 28509 11253 28543
rect 11287 28540 11299 28543
rect 11422 28540 11428 28552
rect 11287 28512 11428 28540
rect 11287 28509 11299 28512
rect 11241 28503 11299 28509
rect 10318 28432 10324 28484
rect 10376 28432 10382 28484
rect 10781 28475 10839 28481
rect 10781 28472 10793 28475
rect 10520 28444 10793 28472
rect 10520 28404 10548 28444
rect 10781 28441 10793 28444
rect 10827 28441 10839 28475
rect 10888 28472 10916 28500
rect 11164 28472 11192 28503
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 11624 28549 11652 28580
rect 13725 28577 13737 28611
rect 13771 28608 13783 28611
rect 14182 28608 14188 28620
rect 13771 28580 14188 28608
rect 13771 28577 13783 28580
rect 13725 28571 13783 28577
rect 14182 28568 14188 28580
rect 14240 28568 14246 28620
rect 20346 28608 20352 28620
rect 16868 28580 17724 28608
rect 16868 28552 16896 28580
rect 11609 28543 11667 28549
rect 11609 28509 11621 28543
rect 11655 28509 11667 28543
rect 11609 28503 11667 28509
rect 12894 28500 12900 28552
rect 12952 28500 12958 28552
rect 16850 28500 16856 28552
rect 16908 28500 16914 28552
rect 17218 28500 17224 28552
rect 17276 28500 17282 28552
rect 17696 28549 17724 28580
rect 19352 28580 20352 28608
rect 19352 28552 19380 28580
rect 20346 28568 20352 28580
rect 20404 28568 20410 28620
rect 17681 28543 17739 28549
rect 17681 28509 17693 28543
rect 17727 28540 17739 28543
rect 17954 28540 17960 28552
rect 17727 28512 17960 28540
rect 17727 28509 17739 28512
rect 17681 28503 17739 28509
rect 17954 28500 17960 28512
rect 18012 28500 18018 28552
rect 19334 28500 19340 28552
rect 19392 28500 19398 28552
rect 20254 28500 20260 28552
rect 20312 28500 20318 28552
rect 20441 28543 20499 28549
rect 20441 28509 20453 28543
rect 20487 28509 20499 28543
rect 20441 28503 20499 28509
rect 20346 28472 20352 28484
rect 10888 28444 11192 28472
rect 11256 28444 20352 28472
rect 10781 28435 10839 28441
rect 10152 28376 10548 28404
rect 9677 28367 9735 28373
rect 11054 28364 11060 28416
rect 11112 28404 11118 28416
rect 11256 28404 11284 28444
rect 20346 28432 20352 28444
rect 20404 28472 20410 28484
rect 20456 28472 20484 28503
rect 20530 28500 20536 28552
rect 20588 28500 20594 28552
rect 22848 28549 22876 28648
rect 23382 28568 23388 28620
rect 23440 28568 23446 28620
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28509 22891 28543
rect 23109 28543 23167 28549
rect 23109 28540 23121 28543
rect 22833 28503 22891 28509
rect 22940 28512 23121 28540
rect 22002 28472 22008 28484
rect 20404 28444 22008 28472
rect 20404 28432 20410 28444
rect 22002 28432 22008 28444
rect 22060 28472 22066 28484
rect 22940 28472 22968 28512
rect 23109 28509 23121 28512
rect 23155 28509 23167 28543
rect 23109 28503 23167 28509
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28540 23259 28543
rect 23400 28540 23428 28568
rect 23247 28512 23428 28540
rect 23661 28543 23719 28549
rect 23247 28509 23259 28512
rect 23201 28503 23259 28509
rect 23661 28509 23673 28543
rect 23707 28509 23719 28543
rect 23661 28503 23719 28509
rect 22060 28444 22968 28472
rect 22060 28432 22066 28444
rect 23014 28432 23020 28484
rect 23072 28432 23078 28484
rect 23216 28472 23244 28503
rect 23124 28444 23244 28472
rect 11112 28376 11284 28404
rect 11112 28364 11118 28376
rect 11698 28364 11704 28416
rect 11756 28364 11762 28416
rect 17862 28364 17868 28416
rect 17920 28364 17926 28416
rect 19978 28364 19984 28416
rect 20036 28404 20042 28416
rect 20073 28407 20131 28413
rect 20073 28404 20085 28407
rect 20036 28376 20085 28404
rect 20036 28364 20042 28376
rect 20073 28373 20085 28376
rect 20119 28373 20131 28407
rect 20073 28367 20131 28373
rect 22646 28364 22652 28416
rect 22704 28404 22710 28416
rect 23124 28404 23152 28444
rect 23290 28432 23296 28484
rect 23348 28472 23354 28484
rect 23676 28472 23704 28503
rect 23348 28444 23704 28472
rect 23765 28472 23793 28648
rect 24210 28636 24216 28688
rect 24268 28636 24274 28688
rect 26510 28636 26516 28688
rect 26568 28636 26574 28688
rect 28948 28676 28954 28688
rect 28184 28648 28954 28676
rect 26528 28608 26556 28636
rect 26789 28611 26847 28617
rect 23860 28580 24532 28608
rect 23860 28552 23888 28580
rect 24504 28552 24532 28580
rect 25332 28580 25728 28608
rect 26528 28580 26648 28608
rect 23842 28500 23848 28552
rect 23900 28500 23906 28552
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28540 24087 28543
rect 24210 28540 24216 28552
rect 24075 28512 24216 28540
rect 24075 28509 24087 28512
rect 24029 28503 24087 28509
rect 24210 28500 24216 28512
rect 24268 28500 24274 28552
rect 24486 28500 24492 28552
rect 24544 28500 24550 28552
rect 23937 28475 23995 28481
rect 23937 28472 23949 28475
rect 23765 28444 23949 28472
rect 23348 28432 23354 28444
rect 22704 28376 23152 28404
rect 22704 28364 22710 28376
rect 23198 28364 23204 28416
rect 23256 28404 23262 28416
rect 23385 28407 23443 28413
rect 23385 28404 23397 28407
rect 23256 28376 23397 28404
rect 23256 28364 23262 28376
rect 23385 28373 23397 28376
rect 23431 28373 23443 28407
rect 23676 28404 23704 28444
rect 23937 28441 23949 28444
rect 23983 28472 23995 28475
rect 25332 28472 25360 28580
rect 25409 28543 25467 28549
rect 25409 28509 25421 28543
rect 25455 28534 25467 28543
rect 25498 28534 25504 28552
rect 25455 28509 25504 28534
rect 25409 28506 25504 28509
rect 25409 28503 25467 28506
rect 23983 28444 25360 28472
rect 23983 28441 23995 28444
rect 23937 28435 23995 28441
rect 25424 28404 25452 28503
rect 25498 28500 25504 28506
rect 25556 28500 25562 28552
rect 25700 28484 25728 28580
rect 26620 28552 26648 28580
rect 26789 28577 26801 28611
rect 26835 28608 26847 28611
rect 27062 28608 27068 28620
rect 26835 28580 27068 28608
rect 26835 28577 26847 28580
rect 26789 28571 26847 28577
rect 27062 28568 27068 28580
rect 27120 28568 27126 28620
rect 25777 28543 25835 28549
rect 25777 28509 25789 28543
rect 25823 28540 25835 28543
rect 25866 28540 25872 28552
rect 25823 28512 25872 28540
rect 25823 28509 25835 28512
rect 25777 28503 25835 28509
rect 25866 28500 25872 28512
rect 25924 28500 25930 28552
rect 26234 28500 26240 28552
rect 26292 28500 26298 28552
rect 26326 28500 26332 28552
rect 26384 28500 26390 28552
rect 26513 28543 26571 28549
rect 26513 28509 26525 28543
rect 26559 28509 26571 28543
rect 26513 28503 26571 28509
rect 25593 28475 25651 28481
rect 25593 28441 25605 28475
rect 25639 28441 25651 28475
rect 25593 28435 25651 28441
rect 23676 28376 25452 28404
rect 25608 28404 25636 28435
rect 25682 28432 25688 28484
rect 25740 28432 25746 28484
rect 26528 28472 26556 28503
rect 26602 28500 26608 28552
rect 26660 28500 26666 28552
rect 25976 28444 26556 28472
rect 25774 28404 25780 28416
rect 25608 28376 25780 28404
rect 23385 28367 23443 28373
rect 25774 28364 25780 28376
rect 25832 28364 25838 28416
rect 25976 28413 26004 28444
rect 27062 28432 27068 28484
rect 27120 28432 27126 28484
rect 25961 28407 26019 28413
rect 25961 28373 25973 28407
rect 26007 28373 26019 28407
rect 25961 28367 26019 28373
rect 26050 28364 26056 28416
rect 26108 28364 26114 28416
rect 27890 28364 27896 28416
rect 27948 28404 27954 28416
rect 28184 28404 28212 28648
rect 28948 28636 28954 28648
rect 29006 28636 29012 28688
rect 29104 28648 29316 28676
rect 28813 28611 28871 28617
rect 28813 28577 28825 28611
rect 28859 28608 28871 28611
rect 29104 28608 29132 28648
rect 28859 28580 29132 28608
rect 29288 28608 29316 28648
rect 29288 28580 29408 28608
rect 28859 28577 28871 28580
rect 28813 28571 28871 28577
rect 29181 28559 29239 28565
rect 29181 28552 29193 28559
rect 29227 28552 29239 28559
rect 28721 28543 28779 28549
rect 28721 28509 28733 28543
rect 28767 28540 28779 28543
rect 29086 28540 29092 28552
rect 28767 28512 29092 28540
rect 28767 28509 28779 28512
rect 28721 28503 28779 28509
rect 29086 28500 29092 28512
rect 29144 28500 29150 28552
rect 29178 28500 29184 28552
rect 29236 28500 29242 28552
rect 29380 28536 29408 28580
rect 33134 28568 33140 28620
rect 33192 28608 33198 28620
rect 34790 28608 34796 28620
rect 33192 28580 34796 28608
rect 33192 28568 33198 28580
rect 34790 28568 34796 28580
rect 34848 28568 34854 28620
rect 29549 28543 29607 28549
rect 29549 28536 29561 28543
rect 29380 28509 29561 28536
rect 29595 28509 29607 28543
rect 29380 28508 29607 28509
rect 29549 28503 29607 28508
rect 31478 28500 31484 28552
rect 31536 28500 31542 28552
rect 33042 28500 33048 28552
rect 33100 28540 33106 28552
rect 34149 28543 34207 28549
rect 34149 28540 34161 28543
rect 33100 28512 34161 28540
rect 33100 28500 33106 28512
rect 34149 28509 34161 28512
rect 34195 28509 34207 28543
rect 34149 28503 34207 28509
rect 34885 28543 34943 28549
rect 34885 28509 34897 28543
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 29825 28475 29883 28481
rect 29825 28472 29837 28475
rect 29472 28444 29837 28472
rect 27948 28376 28212 28404
rect 27948 28364 27954 28376
rect 28534 28364 28540 28416
rect 28592 28364 28598 28416
rect 28997 28407 29055 28413
rect 28997 28373 29009 28407
rect 29043 28404 29055 28407
rect 29472 28404 29500 28444
rect 29825 28441 29837 28444
rect 29871 28441 29883 28475
rect 31386 28472 31392 28484
rect 31050 28444 31392 28472
rect 29825 28435 29883 28441
rect 31386 28432 31392 28444
rect 31444 28432 31450 28484
rect 31754 28432 31760 28484
rect 31812 28432 31818 28484
rect 32140 28444 32246 28472
rect 29043 28376 29500 28404
rect 29043 28373 29055 28376
rect 28997 28367 29055 28373
rect 29730 28364 29736 28416
rect 29788 28404 29794 28416
rect 31297 28407 31355 28413
rect 31297 28404 31309 28407
rect 29788 28376 31309 28404
rect 29788 28364 29794 28376
rect 31297 28373 31309 28376
rect 31343 28373 31355 28407
rect 31404 28404 31432 28432
rect 32140 28404 32168 28444
rect 33502 28432 33508 28484
rect 33560 28472 33566 28484
rect 34900 28472 34928 28503
rect 33560 28444 34928 28472
rect 33560 28432 33566 28444
rect 33134 28404 33140 28416
rect 31404 28376 33140 28404
rect 31297 28367 31355 28373
rect 33134 28364 33140 28376
rect 33192 28364 33198 28416
rect 33226 28364 33232 28416
rect 33284 28364 33290 28416
rect 34238 28364 34244 28416
rect 34296 28364 34302 28416
rect 34514 28364 34520 28416
rect 34572 28404 34578 28416
rect 34701 28407 34759 28413
rect 34701 28404 34713 28407
rect 34572 28376 34713 28404
rect 34572 28364 34578 28376
rect 34701 28373 34713 28376
rect 34747 28373 34759 28407
rect 34701 28367 34759 28373
rect 1104 28314 38272 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38272 28314
rect 1104 28240 38272 28262
rect 4338 28160 4344 28212
rect 4396 28160 4402 28212
rect 6914 28160 6920 28212
rect 6972 28160 6978 28212
rect 9122 28160 9128 28212
rect 9180 28200 9186 28212
rect 17681 28203 17739 28209
rect 9180 28172 17632 28200
rect 9180 28160 9186 28172
rect 4356 28132 4384 28160
rect 4172 28104 4384 28132
rect 4433 28135 4491 28141
rect 4172 28073 4200 28104
rect 4433 28101 4445 28135
rect 4479 28132 4491 28135
rect 4706 28132 4712 28144
rect 4479 28104 4712 28132
rect 4479 28101 4491 28104
rect 4433 28095 4491 28101
rect 4706 28092 4712 28104
rect 4764 28092 4770 28144
rect 6270 28132 6276 28144
rect 5658 28104 6276 28132
rect 6270 28092 6276 28104
rect 6328 28092 6334 28144
rect 6932 28132 6960 28160
rect 11698 28132 11704 28144
rect 6748 28104 6960 28132
rect 11532 28104 11704 28132
rect 6748 28073 6776 28104
rect 4157 28067 4215 28073
rect 4157 28033 4169 28067
rect 4203 28033 4215 28067
rect 4157 28027 4215 28033
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28033 6791 28067
rect 6733 28027 6791 28033
rect 8110 28024 8116 28076
rect 8168 28024 8174 28076
rect 11330 28024 11336 28076
rect 11388 28024 11394 28076
rect 11532 28073 11560 28104
rect 11698 28092 11704 28104
rect 11756 28092 11762 28144
rect 12250 28092 12256 28144
rect 12308 28092 12314 28144
rect 14550 28092 14556 28144
rect 14608 28092 14614 28144
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 14700 28104 15332 28132
rect 14700 28092 14706 28104
rect 11517 28067 11575 28073
rect 11517 28033 11529 28067
rect 11563 28033 11575 28067
rect 11517 28027 11575 28033
rect 14366 28024 14372 28076
rect 14424 28024 14430 28076
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28064 14519 28067
rect 14734 28064 14740 28076
rect 14507 28036 14740 28064
rect 14507 28033 14519 28036
rect 14461 28027 14519 28033
rect 14734 28024 14740 28036
rect 14792 28024 14798 28076
rect 14829 28067 14887 28073
rect 14829 28033 14841 28067
rect 14875 28064 14887 28067
rect 15194 28064 15200 28076
rect 14875 28036 15200 28064
rect 14875 28033 14887 28036
rect 14829 28027 14887 28033
rect 15194 28024 15200 28036
rect 15252 28024 15258 28076
rect 7006 27956 7012 28008
rect 7064 27956 7070 28008
rect 11793 27999 11851 28005
rect 11793 27996 11805 27999
rect 11624 27968 11805 27996
rect 11054 27928 11060 27940
rect 8036 27900 11060 27928
rect 5902 27820 5908 27872
rect 5960 27860 5966 27872
rect 8036 27860 8064 27900
rect 11054 27888 11060 27900
rect 11112 27888 11118 27940
rect 11149 27931 11207 27937
rect 11149 27897 11161 27931
rect 11195 27928 11207 27931
rect 11624 27928 11652 27968
rect 11793 27965 11805 27968
rect 11839 27965 11851 27999
rect 11793 27959 11851 27965
rect 13262 27956 13268 28008
rect 13320 27996 13326 28008
rect 15304 28005 15332 28104
rect 16482 28092 16488 28144
rect 16540 28132 16546 28144
rect 17313 28135 17371 28141
rect 17313 28132 17325 28135
rect 16540 28104 17325 28132
rect 16540 28092 16546 28104
rect 17313 28101 17325 28104
rect 17359 28101 17371 28135
rect 17313 28095 17371 28101
rect 15381 28067 15439 28073
rect 15381 28033 15393 28067
rect 15427 28033 15439 28067
rect 15381 28027 15439 28033
rect 15565 28067 15623 28073
rect 15565 28033 15577 28067
rect 15611 28064 15623 28067
rect 16114 28064 16120 28076
rect 15611 28036 16120 28064
rect 15611 28033 15623 28036
rect 15565 28027 15623 28033
rect 15289 27999 15347 28005
rect 13320 27968 14596 27996
rect 13320 27956 13326 27968
rect 14568 27940 14596 27968
rect 15289 27965 15301 27999
rect 15335 27965 15347 27999
rect 15396 27996 15424 28027
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 17129 28067 17187 28073
rect 17129 28033 17141 28067
rect 17175 28033 17187 28067
rect 17129 28027 17187 28033
rect 17144 27996 17172 28027
rect 17402 28024 17408 28076
rect 17460 28024 17466 28076
rect 17494 28024 17500 28076
rect 17552 28024 17558 28076
rect 17604 28064 17632 28172
rect 17681 28169 17693 28203
rect 17727 28169 17739 28203
rect 17681 28163 17739 28169
rect 17696 28132 17724 28163
rect 17954 28160 17960 28212
rect 18012 28200 18018 28212
rect 18782 28200 18788 28212
rect 18012 28172 18788 28200
rect 18012 28160 18018 28172
rect 18782 28160 18788 28172
rect 18840 28200 18846 28212
rect 19261 28203 19319 28209
rect 19261 28200 19273 28203
rect 18840 28172 19273 28200
rect 18840 28160 18846 28172
rect 19261 28169 19273 28172
rect 19307 28169 19319 28203
rect 19261 28163 19319 28169
rect 19429 28203 19487 28209
rect 19429 28169 19441 28203
rect 19475 28169 19487 28203
rect 20530 28200 20536 28212
rect 19429 28163 19487 28169
rect 20180 28172 20536 28200
rect 17770 28132 17776 28144
rect 17696 28104 17776 28132
rect 17770 28092 17776 28104
rect 17828 28092 17834 28144
rect 19061 28135 19119 28141
rect 19061 28132 19073 28135
rect 18064 28104 19073 28132
rect 18064 28064 18092 28104
rect 19061 28101 19073 28104
rect 19107 28101 19119 28135
rect 19061 28095 19119 28101
rect 17604 28036 18092 28064
rect 18138 28024 18144 28076
rect 18196 28024 18202 28076
rect 18156 27996 18184 28024
rect 15396 27968 18184 27996
rect 19076 27996 19104 28095
rect 19444 28064 19472 28163
rect 20180 28076 20208 28172
rect 20530 28160 20536 28172
rect 20588 28160 20594 28212
rect 20809 28203 20867 28209
rect 20809 28169 20821 28203
rect 20855 28169 20867 28203
rect 20809 28163 20867 28169
rect 20346 28132 20352 28144
rect 20272 28104 20352 28132
rect 19705 28067 19763 28073
rect 19705 28064 19717 28067
rect 19444 28036 19717 28064
rect 19705 28033 19717 28036
rect 19751 28033 19763 28067
rect 19705 28027 19763 28033
rect 19981 28067 20039 28073
rect 19981 28033 19993 28067
rect 20027 28064 20039 28067
rect 20070 28064 20076 28076
rect 20027 28036 20076 28064
rect 20027 28033 20039 28036
rect 19981 28027 20039 28033
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 20162 28024 20168 28076
rect 20220 28024 20226 28076
rect 20272 28073 20300 28104
rect 20346 28092 20352 28104
rect 20404 28092 20410 28144
rect 20441 28135 20499 28141
rect 20441 28101 20453 28135
rect 20487 28132 20499 28135
rect 20714 28132 20720 28144
rect 20487 28104 20720 28132
rect 20487 28101 20499 28104
rect 20441 28095 20499 28101
rect 20714 28092 20720 28104
rect 20772 28092 20778 28144
rect 20258 28067 20316 28073
rect 20258 28033 20270 28067
rect 20304 28033 20316 28067
rect 20258 28027 20316 28033
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28033 20591 28067
rect 20533 28027 20591 28033
rect 20630 28067 20688 28073
rect 20630 28033 20642 28067
rect 20676 28033 20688 28067
rect 20824 28064 20852 28163
rect 21082 28160 21088 28212
rect 21140 28200 21146 28212
rect 22002 28200 22008 28212
rect 21140 28172 22008 28200
rect 21140 28160 21146 28172
rect 22002 28160 22008 28172
rect 22060 28160 22066 28212
rect 22094 28160 22100 28212
rect 22152 28160 22158 28212
rect 22189 28203 22247 28209
rect 22189 28169 22201 28203
rect 22235 28200 22247 28203
rect 22738 28200 22744 28212
rect 22235 28172 22744 28200
rect 22235 28169 22247 28172
rect 22189 28163 22247 28169
rect 22738 28160 22744 28172
rect 22796 28160 22802 28212
rect 22922 28160 22928 28212
rect 22980 28200 22986 28212
rect 22980 28172 24072 28200
rect 22980 28160 22986 28172
rect 21818 28092 21824 28144
rect 21876 28132 21882 28144
rect 22554 28132 22560 28144
rect 21876 28104 22560 28132
rect 21876 28092 21882 28104
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 22812 28104 23336 28132
rect 21177 28067 21235 28073
rect 21177 28064 21189 28067
rect 20824 28036 21189 28064
rect 20630 28027 20688 28033
rect 21177 28033 21189 28036
rect 21223 28033 21235 28067
rect 21177 28027 21235 28033
rect 20548 27996 20576 28027
rect 19076 27968 20576 27996
rect 20645 27996 20673 28027
rect 21266 28024 21272 28076
rect 21324 28024 21330 28076
rect 22278 28064 22284 28076
rect 21376 28036 22284 28064
rect 21376 27996 21404 28036
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22812 28073 22840 28104
rect 23308 28076 23336 28104
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28064 22431 28067
rect 22649 28067 22707 28073
rect 22649 28064 22661 28067
rect 22419 28036 22661 28064
rect 22419 28033 22431 28036
rect 22373 28027 22431 28033
rect 22649 28033 22661 28036
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 22797 28067 22855 28073
rect 22797 28033 22809 28067
rect 22843 28033 22855 28067
rect 22797 28027 22855 28033
rect 22922 28024 22928 28076
rect 22980 28024 22986 28076
rect 23017 28067 23075 28073
rect 23017 28033 23029 28067
rect 23063 28033 23075 28067
rect 23017 28027 23075 28033
rect 20645 27968 21404 27996
rect 15289 27959 15347 27965
rect 11195 27900 11652 27928
rect 11195 27897 11207 27900
rect 11149 27891 11207 27897
rect 14182 27888 14188 27940
rect 14240 27888 14246 27940
rect 14550 27888 14556 27940
rect 14608 27888 14614 27940
rect 14737 27931 14795 27937
rect 14737 27897 14749 27931
rect 14783 27928 14795 27931
rect 15197 27931 15255 27937
rect 15197 27928 15209 27931
rect 14783 27900 15209 27928
rect 14783 27897 14795 27900
rect 14737 27891 14795 27897
rect 15197 27897 15209 27900
rect 15243 27897 15255 27931
rect 15197 27891 15255 27897
rect 15378 27888 15384 27940
rect 15436 27888 15442 27940
rect 16298 27888 16304 27940
rect 16356 27928 16362 27940
rect 19426 27928 19432 27940
rect 16356 27900 19432 27928
rect 16356 27888 16362 27900
rect 19426 27888 19432 27900
rect 19484 27888 19490 27940
rect 19794 27888 19800 27940
rect 19852 27888 19858 27940
rect 19889 27931 19947 27937
rect 19889 27897 19901 27931
rect 19935 27928 19947 27931
rect 19978 27928 19984 27940
rect 19935 27900 19984 27928
rect 19935 27897 19947 27900
rect 19889 27891 19947 27897
rect 19978 27888 19984 27900
rect 20036 27888 20042 27940
rect 20548 27928 20576 27968
rect 21450 27956 21456 28008
rect 21508 27996 21514 28008
rect 21545 27999 21603 28005
rect 21545 27996 21557 27999
rect 21508 27968 21557 27996
rect 21508 27956 21514 27968
rect 21545 27965 21557 27968
rect 21591 27996 21603 27999
rect 21726 27996 21732 28008
rect 21591 27968 21732 27996
rect 21591 27965 21603 27968
rect 21545 27959 21603 27965
rect 21726 27956 21732 27968
rect 21784 27956 21790 28008
rect 23032 27996 23060 28027
rect 23106 28024 23112 28076
rect 23164 28073 23170 28076
rect 23164 28064 23172 28073
rect 23164 28036 23209 28064
rect 23164 28027 23172 28036
rect 23164 28024 23170 28027
rect 23290 28024 23296 28076
rect 23348 28024 23354 28076
rect 23382 28024 23388 28076
rect 23440 28024 23446 28076
rect 23493 28073 23521 28172
rect 23566 28092 23572 28144
rect 23624 28092 23630 28144
rect 23661 28135 23719 28141
rect 23661 28101 23673 28135
rect 23707 28132 23719 28135
rect 23934 28132 23940 28144
rect 23707 28104 23940 28132
rect 23707 28101 23719 28104
rect 23661 28095 23719 28101
rect 23934 28092 23940 28104
rect 23992 28092 23998 28144
rect 23478 28067 23536 28073
rect 23478 28033 23490 28067
rect 23524 28033 23536 28067
rect 23584 28064 23612 28092
rect 23753 28067 23811 28073
rect 23753 28064 23765 28067
rect 23584 28036 23765 28064
rect 23478 28027 23536 28033
rect 23753 28033 23765 28036
rect 23799 28033 23811 28067
rect 23753 28027 23811 28033
rect 23850 28067 23908 28073
rect 23850 28033 23862 28067
rect 23896 28064 23908 28067
rect 23896 28036 23980 28064
rect 23896 28033 23908 28036
rect 23850 28027 23908 28033
rect 23952 27996 23980 28036
rect 22572 27968 23060 27996
rect 23216 27968 23980 27996
rect 22370 27928 22376 27940
rect 20548 27900 22376 27928
rect 22370 27888 22376 27900
rect 22428 27928 22434 27940
rect 22572 27928 22600 27968
rect 22428 27900 22600 27928
rect 22428 27888 22434 27900
rect 22646 27888 22652 27940
rect 22704 27928 22710 27940
rect 22922 27928 22928 27940
rect 22704 27900 22928 27928
rect 22704 27888 22710 27900
rect 22922 27888 22928 27900
rect 22980 27888 22986 27940
rect 5960 27832 8064 27860
rect 5960 27820 5966 27832
rect 8386 27820 8392 27872
rect 8444 27860 8450 27872
rect 8481 27863 8539 27869
rect 8481 27860 8493 27863
rect 8444 27832 8493 27860
rect 8444 27820 8450 27832
rect 8481 27829 8493 27832
rect 8527 27860 8539 27863
rect 11514 27860 11520 27872
rect 8527 27832 11520 27860
rect 8527 27829 8539 27832
rect 8481 27823 8539 27829
rect 11514 27820 11520 27832
rect 11572 27820 11578 27872
rect 15105 27863 15163 27869
rect 15105 27829 15117 27863
rect 15151 27860 15163 27863
rect 15396 27860 15424 27888
rect 15151 27832 15424 27860
rect 15151 27829 15163 27832
rect 15105 27823 15163 27829
rect 16758 27820 16764 27872
rect 16816 27860 16822 27872
rect 17218 27860 17224 27872
rect 16816 27832 17224 27860
rect 16816 27820 16822 27832
rect 17218 27820 17224 27832
rect 17276 27860 17282 27872
rect 19245 27863 19303 27869
rect 19245 27860 19257 27863
rect 17276 27832 19257 27860
rect 17276 27820 17282 27832
rect 19245 27829 19257 27832
rect 19291 27860 19303 27863
rect 19334 27860 19340 27872
rect 19291 27832 19340 27860
rect 19291 27829 19303 27832
rect 19245 27823 19303 27829
rect 19334 27820 19340 27832
rect 19392 27820 19398 27872
rect 19518 27820 19524 27872
rect 19576 27820 19582 27872
rect 20990 27820 20996 27872
rect 21048 27820 21054 27872
rect 21450 27820 21456 27872
rect 21508 27820 21514 27872
rect 21634 27820 21640 27872
rect 21692 27860 21698 27872
rect 23216 27860 23244 27968
rect 24044 27928 24072 28172
rect 25406 28160 25412 28212
rect 25464 28160 25470 28212
rect 26050 28160 26056 28212
rect 26108 28200 26114 28212
rect 26108 28172 26280 28200
rect 26108 28160 26114 28172
rect 25424 28132 25452 28160
rect 25424 28104 26188 28132
rect 26160 28076 26188 28104
rect 24118 28024 24124 28076
rect 24176 28064 24182 28076
rect 26053 28067 26111 28073
rect 26053 28064 26065 28067
rect 24176 28036 26065 28064
rect 24176 28024 24182 28036
rect 26053 28033 26065 28036
rect 26099 28033 26111 28067
rect 26053 28027 26111 28033
rect 26142 28024 26148 28076
rect 26200 28024 26206 28076
rect 26252 28073 26280 28172
rect 27062 28160 27068 28212
rect 27120 28160 27126 28212
rect 28721 28203 28779 28209
rect 28721 28169 28733 28203
rect 28767 28200 28779 28203
rect 29178 28200 29184 28212
rect 28767 28172 29184 28200
rect 28767 28169 28779 28172
rect 28721 28163 28779 28169
rect 29178 28160 29184 28172
rect 29236 28160 29242 28212
rect 30285 28203 30343 28209
rect 30285 28169 30297 28203
rect 30331 28169 30343 28203
rect 30285 28163 30343 28169
rect 26970 28092 26976 28144
rect 27028 28132 27034 28144
rect 27028 28104 28994 28132
rect 27028 28092 27034 28104
rect 28966 28100 28994 28104
rect 29380 28104 29776 28132
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28033 26295 28067
rect 26237 28027 26295 28033
rect 26421 28067 26479 28073
rect 26421 28033 26433 28067
rect 26467 28064 26479 28067
rect 26694 28064 26700 28076
rect 26467 28036 26700 28064
rect 26467 28033 26479 28036
rect 26421 28027 26479 28033
rect 26694 28024 26700 28036
rect 26752 28024 26758 28076
rect 26786 28024 26792 28076
rect 26844 28024 26850 28076
rect 27246 28024 27252 28076
rect 27304 28024 27310 28076
rect 28966 28060 29000 28100
rect 28994 28048 29000 28060
rect 29052 28048 29058 28100
rect 29086 28024 29092 28076
rect 29144 28024 29150 28076
rect 29181 28067 29239 28073
rect 29181 28033 29193 28067
rect 29227 28064 29239 28067
rect 29380 28064 29408 28104
rect 29748 28076 29776 28104
rect 29914 28092 29920 28144
rect 29972 28092 29978 28144
rect 30006 28092 30012 28144
rect 30064 28092 30070 28144
rect 29227 28036 29408 28064
rect 29227 28033 29239 28036
rect 29181 28027 29239 28033
rect 25777 27999 25835 28005
rect 25777 27965 25789 27999
rect 25823 27996 25835 27999
rect 26804 27996 26832 28024
rect 25823 27968 26832 27996
rect 25823 27965 25835 27968
rect 25777 27959 25835 27965
rect 28810 27956 28816 28008
rect 28868 27996 28874 28008
rect 29273 27999 29331 28005
rect 29273 27996 29285 27999
rect 28868 27968 29285 27996
rect 28868 27956 28874 27968
rect 29273 27965 29285 27968
rect 29319 27965 29331 27999
rect 29273 27959 29331 27965
rect 26326 27928 26332 27940
rect 24044 27900 26332 27928
rect 26326 27888 26332 27900
rect 26384 27928 26390 27940
rect 29380 27928 29408 28036
rect 29454 28024 29460 28076
rect 29512 28068 29518 28076
rect 29512 28064 29592 28068
rect 29641 28067 29699 28073
rect 29641 28064 29653 28067
rect 29512 28040 29653 28064
rect 29512 28024 29518 28040
rect 29564 28036 29653 28040
rect 29641 28033 29653 28036
rect 29687 28033 29699 28067
rect 29641 28027 29699 28033
rect 29730 28024 29736 28076
rect 29788 28064 29794 28076
rect 30024 28064 30052 28092
rect 29788 28036 29833 28064
rect 29932 28036 30052 28064
rect 29788 28024 29794 28036
rect 26384 27900 29408 27928
rect 29932 27928 29960 28036
rect 30098 28024 30104 28076
rect 30156 28073 30162 28076
rect 30156 28064 30164 28073
rect 30300 28064 30328 28163
rect 31754 28160 31760 28212
rect 31812 28160 31818 28212
rect 32125 28203 32183 28209
rect 32125 28169 32137 28203
rect 32171 28169 32183 28203
rect 32125 28163 32183 28169
rect 30374 28092 30380 28144
rect 30432 28132 30438 28144
rect 30745 28135 30803 28141
rect 30745 28132 30757 28135
rect 30432 28104 30757 28132
rect 30432 28092 30438 28104
rect 30745 28101 30757 28104
rect 30791 28101 30803 28135
rect 30745 28095 30803 28101
rect 30561 28067 30619 28073
rect 30561 28064 30573 28067
rect 30156 28036 30201 28064
rect 30300 28036 30573 28064
rect 30156 28027 30164 28036
rect 30561 28033 30573 28036
rect 30607 28033 30619 28067
rect 30561 28027 30619 28033
rect 30156 28024 30162 28027
rect 30760 27996 30788 28095
rect 30834 28024 30840 28076
rect 30892 28024 30898 28076
rect 31941 28067 31999 28073
rect 31941 28033 31953 28067
rect 31987 28064 31999 28067
rect 32140 28064 32168 28163
rect 34238 28160 34244 28212
rect 34296 28160 34302 28212
rect 34514 28200 34520 28212
rect 34348 28172 34520 28200
rect 33689 28135 33747 28141
rect 33689 28132 33701 28135
rect 32508 28104 33701 28132
rect 32508 28076 32536 28104
rect 33689 28101 33701 28104
rect 33735 28132 33747 28135
rect 33962 28132 33968 28144
rect 33735 28104 33968 28132
rect 33735 28101 33747 28104
rect 33689 28095 33747 28101
rect 33962 28092 33968 28104
rect 34020 28092 34026 28144
rect 34256 28132 34284 28160
rect 34348 28141 34376 28172
rect 34514 28160 34520 28172
rect 34572 28160 34578 28212
rect 34072 28104 34284 28132
rect 34333 28135 34391 28141
rect 31987 28036 32168 28064
rect 31987 28033 31999 28036
rect 31941 28027 31999 28033
rect 32490 28024 32496 28076
rect 32548 28024 32554 28076
rect 33226 28064 33232 28076
rect 32600 28036 33232 28064
rect 32600 28005 32628 28036
rect 33226 28024 33232 28036
rect 33284 28024 33290 28076
rect 33502 28024 33508 28076
rect 33560 28024 33566 28076
rect 34072 28073 34100 28104
rect 34333 28101 34345 28135
rect 34379 28101 34391 28135
rect 34333 28095 34391 28101
rect 34790 28092 34796 28144
rect 34848 28092 34854 28144
rect 33597 28067 33655 28073
rect 33597 28033 33609 28067
rect 33643 28064 33655 28067
rect 34057 28067 34115 28073
rect 33643 28036 33916 28064
rect 33643 28033 33655 28036
rect 33597 28027 33655 28033
rect 32585 27999 32643 28005
rect 32585 27996 32597 27999
rect 30760 27968 32597 27996
rect 32585 27965 32597 27968
rect 32631 27965 32643 27999
rect 32585 27959 32643 27965
rect 32766 27956 32772 28008
rect 32824 27956 32830 28008
rect 33229 27931 33287 27937
rect 29932 27900 30512 27928
rect 26384 27888 26390 27900
rect 21692 27832 23244 27860
rect 21692 27820 21698 27832
rect 23290 27820 23296 27872
rect 23348 27820 23354 27872
rect 23750 27820 23756 27872
rect 23808 27860 23814 27872
rect 24029 27863 24087 27869
rect 24029 27860 24041 27863
rect 23808 27832 24041 27860
rect 23808 27820 23814 27832
rect 24029 27829 24041 27832
rect 24075 27829 24087 27863
rect 24029 27823 24087 27829
rect 25682 27820 25688 27872
rect 25740 27860 25746 27872
rect 30282 27860 30288 27872
rect 25740 27832 30288 27860
rect 25740 27820 25746 27832
rect 30282 27820 30288 27832
rect 30340 27820 30346 27872
rect 30374 27820 30380 27872
rect 30432 27820 30438 27872
rect 30484 27860 30512 27900
rect 33229 27897 33241 27931
rect 33275 27928 33287 27931
rect 33520 27928 33548 28024
rect 33275 27900 33548 27928
rect 33275 27897 33287 27900
rect 33229 27891 33287 27897
rect 33612 27860 33640 28027
rect 33778 27956 33784 28008
rect 33836 27956 33842 28008
rect 33888 27996 33916 28036
rect 34057 28033 34069 28067
rect 34103 28033 34115 28067
rect 34057 28027 34115 28033
rect 35805 27999 35863 28005
rect 35805 27996 35817 27999
rect 33888 27968 35817 27996
rect 35805 27965 35817 27968
rect 35851 27965 35863 27999
rect 35805 27959 35863 27965
rect 30484 27832 33640 27860
rect 1104 27770 38272 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38272 27770
rect 1104 27696 38272 27718
rect 4706 27616 4712 27668
rect 4764 27616 4770 27668
rect 7006 27616 7012 27668
rect 7064 27656 7070 27668
rect 7193 27659 7251 27665
rect 7193 27656 7205 27659
rect 7064 27628 7205 27656
rect 7064 27616 7070 27628
rect 7193 27625 7205 27628
rect 7239 27625 7251 27659
rect 7193 27619 7251 27625
rect 8110 27616 8116 27668
rect 8168 27656 8174 27668
rect 8662 27656 8668 27668
rect 8168 27628 8668 27656
rect 8168 27616 8174 27628
rect 8662 27616 8668 27628
rect 8720 27616 8726 27668
rect 11330 27616 11336 27668
rect 11388 27656 11394 27668
rect 11609 27659 11667 27665
rect 11609 27656 11621 27659
rect 11388 27628 11621 27656
rect 11388 27616 11394 27628
rect 11609 27625 11621 27628
rect 11655 27625 11667 27659
rect 11609 27619 11667 27625
rect 11790 27616 11796 27668
rect 11848 27656 11854 27668
rect 11848 27628 19748 27656
rect 11848 27616 11854 27628
rect 7653 27591 7711 27597
rect 7653 27557 7665 27591
rect 7699 27557 7711 27591
rect 7653 27551 7711 27557
rect 8128 27560 8892 27588
rect 6089 27523 6147 27529
rect 6089 27489 6101 27523
rect 6135 27520 6147 27523
rect 6822 27520 6828 27532
rect 6135 27492 6828 27520
rect 6135 27489 6147 27492
rect 6089 27483 6147 27489
rect 6822 27480 6828 27492
rect 6880 27480 6886 27532
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27452 4951 27455
rect 5813 27455 5871 27461
rect 4939 27424 5488 27452
rect 4939 27421 4951 27424
rect 4893 27415 4951 27421
rect 5460 27325 5488 27424
rect 5813 27421 5825 27455
rect 5859 27452 5871 27455
rect 5902 27452 5908 27464
rect 5859 27424 5908 27452
rect 5859 27421 5871 27424
rect 5813 27415 5871 27421
rect 5902 27412 5908 27424
rect 5960 27412 5966 27464
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27452 7435 27455
rect 7668 27452 7696 27551
rect 8128 27529 8156 27560
rect 8864 27532 8892 27560
rect 10594 27548 10600 27600
rect 10652 27588 10658 27600
rect 11698 27588 11704 27600
rect 10652 27560 11704 27588
rect 10652 27548 10658 27560
rect 11698 27548 11704 27560
rect 11756 27588 11762 27600
rect 12066 27588 12072 27600
rect 11756 27560 12072 27588
rect 11756 27548 11762 27560
rect 12066 27548 12072 27560
rect 12124 27548 12130 27600
rect 13262 27588 13268 27600
rect 13096 27560 13268 27588
rect 8113 27523 8171 27529
rect 8113 27520 8125 27523
rect 7423 27424 7696 27452
rect 7760 27492 8125 27520
rect 7423 27421 7435 27424
rect 7377 27415 7435 27421
rect 6730 27344 6736 27396
rect 6788 27384 6794 27396
rect 7760 27384 7788 27492
rect 8113 27489 8125 27492
rect 8159 27489 8171 27523
rect 8113 27483 8171 27489
rect 8205 27523 8263 27529
rect 8205 27489 8217 27523
rect 8251 27520 8263 27523
rect 8251 27492 8800 27520
rect 8251 27489 8263 27492
rect 8205 27483 8263 27489
rect 8021 27455 8079 27461
rect 8021 27421 8033 27455
rect 8067 27452 8079 27455
rect 8386 27452 8392 27464
rect 8067 27424 8392 27452
rect 8067 27421 8079 27424
rect 8021 27415 8079 27421
rect 8386 27412 8392 27424
rect 8444 27412 8450 27464
rect 8478 27412 8484 27464
rect 8536 27412 8542 27464
rect 8772 27452 8800 27492
rect 8846 27480 8852 27532
rect 8904 27480 8910 27532
rect 10686 27520 10692 27532
rect 8956 27492 10692 27520
rect 8956 27452 8984 27492
rect 10686 27480 10692 27492
rect 10744 27520 10750 27532
rect 12253 27523 12311 27529
rect 12253 27520 12265 27523
rect 10744 27492 12265 27520
rect 10744 27480 10750 27492
rect 12253 27489 12265 27492
rect 12299 27520 12311 27523
rect 12342 27520 12348 27532
rect 12299 27492 12348 27520
rect 12299 27489 12311 27492
rect 12253 27483 12311 27489
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 13096 27461 13124 27560
rect 13262 27548 13268 27560
rect 13320 27548 13326 27600
rect 14550 27548 14556 27600
rect 14608 27548 14614 27600
rect 14642 27548 14648 27600
rect 14700 27588 14706 27600
rect 15105 27591 15163 27597
rect 15105 27588 15117 27591
rect 14700 27560 15117 27588
rect 14700 27548 14706 27560
rect 15105 27557 15117 27560
rect 15151 27557 15163 27591
rect 15105 27551 15163 27557
rect 15212 27560 16860 27588
rect 13814 27520 13820 27532
rect 13280 27492 13820 27520
rect 8772 27424 8984 27452
rect 11977 27455 12035 27461
rect 11977 27421 11989 27455
rect 12023 27452 12035 27455
rect 13081 27455 13139 27461
rect 13081 27452 13093 27455
rect 12023 27424 13093 27452
rect 12023 27421 12035 27424
rect 11977 27415 12035 27421
rect 13081 27421 13093 27424
rect 13127 27421 13139 27455
rect 13280 27452 13308 27492
rect 13814 27480 13820 27492
rect 13872 27520 13878 27532
rect 14182 27520 14188 27532
rect 13872 27492 14188 27520
rect 13872 27480 13878 27492
rect 14182 27480 14188 27492
rect 14240 27520 14246 27532
rect 15212 27520 15240 27560
rect 14240 27492 15240 27520
rect 14240 27480 14246 27492
rect 15654 27480 15660 27532
rect 15712 27520 15718 27532
rect 15712 27492 16160 27520
rect 15712 27480 15718 27492
rect 13357 27455 13415 27461
rect 13357 27452 13369 27455
rect 13280 27424 13369 27452
rect 13081 27415 13139 27421
rect 13357 27421 13369 27424
rect 13403 27421 13415 27455
rect 13357 27415 13415 27421
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 13630 27452 13636 27464
rect 13495 27424 13636 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 13630 27412 13636 27424
rect 13688 27452 13694 27464
rect 14458 27452 14464 27464
rect 13688 27424 14464 27452
rect 13688 27412 13694 27424
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27452 14979 27455
rect 15470 27452 15476 27464
rect 14967 27424 15476 27452
rect 14967 27421 14979 27424
rect 14921 27415 14979 27421
rect 15470 27412 15476 27424
rect 15528 27412 15534 27464
rect 15746 27412 15752 27464
rect 15804 27412 15810 27464
rect 16022 27452 16028 27464
rect 15856 27424 16028 27452
rect 6788 27356 7788 27384
rect 8496 27384 8524 27412
rect 8496 27356 9444 27384
rect 6788 27344 6794 27356
rect 5445 27319 5503 27325
rect 5445 27285 5457 27319
rect 5491 27285 5503 27319
rect 5445 27279 5503 27285
rect 5905 27319 5963 27325
rect 5905 27285 5917 27319
rect 5951 27316 5963 27319
rect 6748 27316 6776 27344
rect 9416 27328 9444 27356
rect 12618 27344 12624 27396
rect 12676 27384 12682 27396
rect 13265 27387 13323 27393
rect 13265 27384 13277 27387
rect 12676 27356 13277 27384
rect 12676 27344 12682 27356
rect 13265 27353 13277 27356
rect 13311 27353 13323 27387
rect 13265 27347 13323 27353
rect 15378 27344 15384 27396
rect 15436 27384 15442 27396
rect 15856 27384 15884 27424
rect 16022 27412 16028 27424
rect 16080 27412 16086 27464
rect 16132 27461 16160 27492
rect 16117 27455 16175 27461
rect 16117 27421 16129 27455
rect 16163 27452 16175 27455
rect 16482 27452 16488 27464
rect 16163 27424 16488 27452
rect 16163 27421 16175 27424
rect 16117 27415 16175 27421
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 16666 27412 16672 27464
rect 16724 27412 16730 27464
rect 16832 27461 16860 27560
rect 17052 27560 19564 27588
rect 17052 27532 17080 27560
rect 17034 27520 17040 27532
rect 16960 27492 17040 27520
rect 16960 27461 16988 27492
rect 17034 27480 17040 27492
rect 17092 27480 17098 27532
rect 17862 27520 17868 27532
rect 17328 27492 17868 27520
rect 16817 27455 16875 27461
rect 16817 27421 16829 27455
rect 16863 27421 16875 27455
rect 16817 27415 16875 27421
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27421 17003 27455
rect 16945 27415 17003 27421
rect 17175 27455 17233 27461
rect 17175 27421 17187 27455
rect 17221 27452 17233 27455
rect 17328 27452 17356 27492
rect 17862 27480 17868 27492
rect 17920 27520 17926 27532
rect 17920 27480 17954 27520
rect 17221 27424 17356 27452
rect 17221 27421 17233 27424
rect 17175 27415 17233 27421
rect 15436 27356 15884 27384
rect 15436 27344 15442 27356
rect 15930 27344 15936 27396
rect 15988 27344 15994 27396
rect 5951 27288 6776 27316
rect 5951 27285 5963 27288
rect 5905 27279 5963 27285
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 8573 27319 8631 27325
rect 8573 27316 8585 27319
rect 8352 27288 8585 27316
rect 8352 27276 8358 27288
rect 8573 27285 8585 27288
rect 8619 27285 8631 27319
rect 8573 27279 8631 27285
rect 9398 27276 9404 27328
rect 9456 27276 9462 27328
rect 10962 27276 10968 27328
rect 11020 27316 11026 27328
rect 11514 27316 11520 27328
rect 11020 27288 11520 27316
rect 11020 27276 11026 27288
rect 11514 27276 11520 27288
rect 11572 27276 11578 27328
rect 11790 27276 11796 27328
rect 11848 27316 11854 27328
rect 12069 27319 12127 27325
rect 12069 27316 12081 27319
rect 11848 27288 12081 27316
rect 11848 27276 11854 27288
rect 12069 27285 12081 27288
rect 12115 27285 12127 27319
rect 12069 27279 12127 27285
rect 13630 27276 13636 27328
rect 13688 27276 13694 27328
rect 14366 27276 14372 27328
rect 14424 27316 14430 27328
rect 14737 27319 14795 27325
rect 14737 27316 14749 27319
rect 14424 27288 14749 27316
rect 14424 27276 14430 27288
rect 14737 27285 14749 27288
rect 14783 27285 14795 27319
rect 14737 27279 14795 27285
rect 14826 27276 14832 27328
rect 14884 27276 14890 27328
rect 15654 27276 15660 27328
rect 15712 27316 15718 27328
rect 16301 27319 16359 27325
rect 16301 27316 16313 27319
rect 15712 27288 16313 27316
rect 15712 27276 15718 27288
rect 16301 27285 16313 27288
rect 16347 27285 16359 27319
rect 16832 27316 16860 27415
rect 17402 27412 17408 27464
rect 17460 27412 17466 27464
rect 17037 27387 17095 27393
rect 17037 27353 17049 27387
rect 17083 27384 17095 27387
rect 17420 27384 17448 27412
rect 17083 27356 17448 27384
rect 17926 27384 17954 27480
rect 19536 27464 19564 27560
rect 19720 27520 19748 27628
rect 19794 27616 19800 27668
rect 19852 27656 19858 27668
rect 19981 27659 20039 27665
rect 19981 27656 19993 27659
rect 19852 27628 19993 27656
rect 19852 27616 19858 27628
rect 19981 27625 19993 27628
rect 20027 27625 20039 27659
rect 19981 27619 20039 27625
rect 20070 27616 20076 27668
rect 20128 27656 20134 27668
rect 20622 27656 20628 27668
rect 20128 27628 20628 27656
rect 20128 27616 20134 27628
rect 20622 27616 20628 27628
rect 20680 27656 20686 27668
rect 21085 27659 21143 27665
rect 20680 27628 21036 27656
rect 20680 27616 20686 27628
rect 21008 27588 21036 27628
rect 21085 27625 21097 27659
rect 21131 27656 21143 27659
rect 21266 27656 21272 27668
rect 21131 27628 21272 27656
rect 21131 27625 21143 27628
rect 21085 27619 21143 27625
rect 21266 27616 21272 27628
rect 21324 27616 21330 27668
rect 24486 27656 24492 27668
rect 21376 27628 22232 27656
rect 21376 27588 21404 27628
rect 21008 27560 21404 27588
rect 22204 27588 22232 27628
rect 24044 27628 24492 27656
rect 24044 27588 24072 27628
rect 24486 27616 24492 27628
rect 24544 27656 24550 27668
rect 25038 27656 25044 27668
rect 24544 27628 25044 27656
rect 24544 27616 24550 27628
rect 25038 27616 25044 27628
rect 25096 27616 25102 27668
rect 26142 27616 26148 27668
rect 26200 27656 26206 27668
rect 26510 27656 26516 27668
rect 26200 27628 26516 27656
rect 26200 27616 26206 27628
rect 26510 27616 26516 27628
rect 26568 27616 26574 27668
rect 27157 27659 27215 27665
rect 27157 27625 27169 27659
rect 27203 27656 27215 27659
rect 27246 27656 27252 27668
rect 27203 27628 27252 27656
rect 27203 27625 27215 27628
rect 27157 27619 27215 27625
rect 27246 27616 27252 27628
rect 27304 27616 27310 27668
rect 29178 27616 29184 27668
rect 29236 27656 29242 27668
rect 32490 27656 32496 27668
rect 29236 27628 32496 27656
rect 29236 27616 29242 27628
rect 32490 27616 32496 27628
rect 32548 27616 32554 27668
rect 33686 27616 33692 27668
rect 33744 27616 33750 27668
rect 28902 27588 28908 27600
rect 22204 27560 24072 27588
rect 24412 27560 28908 27588
rect 19720 27492 21220 27520
rect 19426 27412 19432 27464
rect 19484 27412 19490 27464
rect 19518 27412 19524 27464
rect 19576 27452 19582 27464
rect 19720 27461 19748 27492
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 19576 27424 19625 27452
rect 19576 27412 19582 27424
rect 19613 27421 19625 27424
rect 19659 27421 19671 27455
rect 19613 27415 19671 27421
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 19812 27384 19840 27415
rect 20070 27412 20076 27464
rect 20128 27452 20134 27464
rect 20438 27452 20444 27464
rect 20128 27424 20444 27452
rect 20128 27412 20134 27424
rect 20438 27412 20444 27424
rect 20496 27412 20502 27464
rect 20548 27461 20576 27492
rect 20548 27455 20611 27461
rect 20548 27424 20565 27455
rect 20553 27421 20565 27424
rect 20599 27421 20611 27455
rect 20553 27415 20611 27421
rect 20806 27412 20812 27464
rect 20864 27412 20870 27464
rect 20901 27455 20959 27461
rect 20901 27421 20913 27455
rect 20947 27452 20959 27455
rect 21082 27452 21088 27464
rect 20947 27424 21088 27452
rect 20947 27421 20959 27424
rect 20901 27415 20959 27421
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 21192 27452 21220 27492
rect 21450 27480 21456 27532
rect 21508 27520 21514 27532
rect 23017 27523 23075 27529
rect 23017 27520 23029 27523
rect 21508 27492 23029 27520
rect 21508 27480 21514 27492
rect 23017 27489 23029 27492
rect 23063 27489 23075 27523
rect 23017 27483 23075 27489
rect 23290 27480 23296 27532
rect 23348 27480 23354 27532
rect 23385 27523 23443 27529
rect 23385 27489 23397 27523
rect 23431 27520 23443 27523
rect 23750 27520 23756 27532
rect 23431 27492 23756 27520
rect 23431 27489 23443 27492
rect 23385 27483 23443 27489
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 21818 27452 21824 27464
rect 21192 27424 21824 27452
rect 21818 27412 21824 27424
rect 21876 27412 21882 27464
rect 22186 27412 22192 27464
rect 22244 27452 22250 27464
rect 22373 27455 22431 27461
rect 22373 27452 22385 27455
rect 22244 27424 22385 27452
rect 22244 27412 22250 27424
rect 22373 27421 22385 27424
rect 22419 27421 22431 27455
rect 22373 27415 22431 27421
rect 19978 27384 19984 27396
rect 17926 27356 19984 27384
rect 17083 27353 17095 27356
rect 17037 27347 17095 27353
rect 19978 27344 19984 27356
rect 20036 27344 20042 27396
rect 20717 27387 20775 27393
rect 20717 27353 20729 27387
rect 20763 27353 20775 27387
rect 20717 27347 20775 27353
rect 17126 27316 17132 27328
rect 16832 27288 17132 27316
rect 16301 27279 16359 27285
rect 17126 27276 17132 27288
rect 17184 27276 17190 27328
rect 17313 27319 17371 27325
rect 17313 27285 17325 27319
rect 17359 27316 17371 27319
rect 18046 27316 18052 27328
rect 17359 27288 18052 27316
rect 17359 27285 17371 27288
rect 17313 27279 17371 27285
rect 18046 27276 18052 27288
rect 18104 27276 18110 27328
rect 20732 27316 20760 27347
rect 20990 27344 20996 27396
rect 21048 27344 21054 27396
rect 22388 27384 22416 27415
rect 22554 27412 22560 27464
rect 22612 27412 22618 27464
rect 23198 27412 23204 27464
rect 23256 27412 23262 27464
rect 23477 27455 23535 27461
rect 23477 27421 23489 27455
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 23382 27384 23388 27396
rect 22388 27356 23388 27384
rect 23382 27344 23388 27356
rect 23440 27344 23446 27396
rect 23492 27384 23520 27415
rect 23658 27412 23664 27464
rect 23716 27412 23722 27464
rect 24118 27412 24124 27464
rect 24176 27412 24182 27464
rect 24136 27384 24164 27412
rect 23492 27356 24164 27384
rect 21008 27316 21036 27344
rect 24412 27328 24440 27560
rect 28902 27548 28908 27560
rect 28960 27588 28966 27600
rect 29914 27588 29920 27600
rect 28960 27560 29920 27588
rect 28960 27548 28966 27560
rect 29914 27548 29920 27560
rect 29972 27548 29978 27600
rect 30374 27548 30380 27600
rect 30432 27588 30438 27600
rect 30561 27591 30619 27597
rect 30561 27588 30573 27591
rect 30432 27560 30573 27588
rect 30432 27548 30438 27560
rect 30561 27557 30573 27560
rect 30607 27557 30619 27591
rect 30561 27551 30619 27557
rect 30650 27548 30656 27600
rect 30708 27588 30714 27600
rect 30834 27588 30840 27600
rect 30708 27560 30840 27588
rect 30708 27548 30714 27560
rect 30834 27548 30840 27560
rect 30892 27548 30898 27600
rect 34698 27548 34704 27600
rect 34756 27548 34762 27600
rect 24578 27480 24584 27532
rect 24636 27520 24642 27532
rect 27709 27523 27767 27529
rect 27709 27520 27721 27523
rect 24636 27492 27721 27520
rect 24636 27480 24642 27492
rect 27709 27489 27721 27492
rect 27755 27520 27767 27523
rect 27755 27492 30972 27520
rect 27755 27489 27767 27492
rect 27709 27483 27767 27489
rect 27522 27412 27528 27464
rect 27580 27452 27586 27464
rect 27617 27455 27675 27461
rect 27617 27452 27629 27455
rect 27580 27424 27629 27452
rect 27580 27412 27586 27424
rect 27617 27421 27629 27424
rect 27663 27421 27675 27455
rect 27617 27415 27675 27421
rect 29086 27412 29092 27464
rect 29144 27452 29150 27464
rect 29362 27452 29368 27464
rect 29144 27424 29368 27452
rect 29144 27412 29150 27424
rect 29362 27412 29368 27424
rect 29420 27412 29426 27464
rect 30742 27412 30748 27464
rect 30800 27412 30806 27464
rect 27798 27384 27804 27396
rect 27540 27356 27804 27384
rect 20732 27288 21036 27316
rect 23014 27276 23020 27328
rect 23072 27316 23078 27328
rect 23566 27316 23572 27328
rect 23072 27288 23572 27316
rect 23072 27276 23078 27288
rect 23566 27276 23572 27288
rect 23624 27276 23630 27328
rect 24394 27276 24400 27328
rect 24452 27276 24458 27328
rect 25590 27276 25596 27328
rect 25648 27316 25654 27328
rect 27540 27325 27568 27356
rect 27798 27344 27804 27356
rect 27856 27344 27862 27396
rect 30653 27387 30711 27393
rect 30653 27353 30665 27387
rect 30699 27384 30711 27387
rect 30834 27384 30840 27396
rect 30699 27356 30840 27384
rect 30699 27353 30711 27356
rect 30653 27347 30711 27353
rect 30834 27344 30840 27356
rect 30892 27344 30898 27396
rect 27525 27319 27583 27325
rect 27525 27316 27537 27319
rect 25648 27288 27537 27316
rect 25648 27276 25654 27288
rect 27525 27285 27537 27288
rect 27571 27285 27583 27319
rect 27525 27279 27583 27285
rect 28626 27276 28632 27328
rect 28684 27316 28690 27328
rect 29454 27316 29460 27328
rect 28684 27288 29460 27316
rect 28684 27276 28690 27288
rect 29454 27276 29460 27288
rect 29512 27276 29518 27328
rect 30944 27316 30972 27492
rect 31018 27412 31024 27464
rect 31076 27452 31082 27464
rect 31202 27452 31208 27464
rect 31076 27424 31208 27452
rect 31076 27412 31082 27424
rect 31202 27412 31208 27424
rect 31260 27412 31266 27464
rect 32398 27452 32404 27464
rect 31726 27424 32404 27452
rect 31294 27344 31300 27396
rect 31352 27384 31358 27396
rect 31389 27387 31447 27393
rect 31389 27384 31401 27387
rect 31352 27356 31401 27384
rect 31352 27344 31358 27356
rect 31389 27353 31401 27356
rect 31435 27384 31447 27387
rect 31726 27384 31754 27424
rect 32398 27412 32404 27424
rect 32456 27412 32462 27464
rect 33505 27455 33563 27461
rect 33505 27421 33517 27455
rect 33551 27452 33563 27455
rect 34716 27452 34744 27548
rect 33551 27424 34744 27452
rect 33551 27421 33563 27424
rect 33505 27415 33563 27421
rect 31435 27356 31754 27384
rect 31435 27353 31447 27356
rect 31389 27347 31447 27353
rect 33778 27316 33784 27328
rect 30944 27288 33784 27316
rect 33778 27276 33784 27288
rect 33836 27276 33842 27328
rect 1104 27226 38272 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38272 27226
rect 1104 27152 38272 27174
rect 6822 27072 6828 27124
rect 6880 27112 6886 27124
rect 6880 27084 11376 27112
rect 6880 27072 6886 27084
rect 8294 27044 8300 27056
rect 8128 27016 8300 27044
rect 5902 26936 5908 26988
rect 5960 26936 5966 26988
rect 8128 26985 8156 27016
rect 8294 27004 8300 27016
rect 8352 27004 8358 27056
rect 8662 27004 8668 27056
rect 8720 27044 8726 27056
rect 10594 27044 10600 27056
rect 8720 27016 8878 27044
rect 10060 27016 10600 27044
rect 8720 27004 8726 27016
rect 8113 26979 8171 26985
rect 8113 26945 8125 26979
rect 8159 26945 8171 26979
rect 8113 26939 8171 26945
rect 8386 26868 8392 26920
rect 8444 26868 8450 26920
rect 10060 26908 10088 27016
rect 10594 27004 10600 27016
rect 10652 27004 10658 27056
rect 10134 26936 10140 26988
rect 10192 26976 10198 26988
rect 10321 26979 10379 26985
rect 10321 26976 10333 26979
rect 10192 26948 10333 26976
rect 10192 26936 10198 26948
rect 10321 26945 10333 26948
rect 10367 26976 10379 26979
rect 10367 26948 10916 26976
rect 10367 26945 10379 26948
rect 10321 26939 10379 26945
rect 9416 26880 10088 26908
rect 10413 26911 10471 26917
rect 5442 26732 5448 26784
rect 5500 26772 5506 26784
rect 5721 26775 5779 26781
rect 5721 26772 5733 26775
rect 5500 26744 5733 26772
rect 5500 26732 5506 26744
rect 5721 26741 5733 26744
rect 5767 26741 5779 26775
rect 5721 26735 5779 26741
rect 7374 26732 7380 26784
rect 7432 26772 7438 26784
rect 7742 26772 7748 26784
rect 7432 26744 7748 26772
rect 7432 26732 7438 26744
rect 7742 26732 7748 26744
rect 7800 26772 7806 26784
rect 9416 26772 9444 26880
rect 10413 26877 10425 26911
rect 10459 26877 10471 26911
rect 10413 26871 10471 26877
rect 9490 26800 9496 26852
rect 9548 26840 9554 26852
rect 9953 26843 10011 26849
rect 9953 26840 9965 26843
rect 9548 26812 9965 26840
rect 9548 26800 9554 26812
rect 9953 26809 9965 26812
rect 9999 26809 10011 26843
rect 9953 26803 10011 26809
rect 10428 26840 10456 26871
rect 10594 26868 10600 26920
rect 10652 26868 10658 26920
rect 10888 26908 10916 26948
rect 10962 26936 10968 26988
rect 11020 26936 11026 26988
rect 11348 26976 11376 27084
rect 11514 27072 11520 27124
rect 11572 27072 11578 27124
rect 15194 27072 15200 27124
rect 15252 27072 15258 27124
rect 16666 27072 16672 27124
rect 16724 27072 16730 27124
rect 16850 27072 16856 27124
rect 16908 27072 16914 27124
rect 16942 27072 16948 27124
rect 17000 27112 17006 27124
rect 17000 27084 17264 27112
rect 17000 27072 17006 27084
rect 11885 27047 11943 27053
rect 11885 27013 11897 27047
rect 11931 27044 11943 27047
rect 11974 27044 11980 27056
rect 11931 27016 11980 27044
rect 11931 27013 11943 27016
rect 11885 27007 11943 27013
rect 11974 27004 11980 27016
rect 12032 27044 12038 27056
rect 12802 27044 12808 27056
rect 12032 27016 12808 27044
rect 12032 27004 12038 27016
rect 12802 27004 12808 27016
rect 12860 27044 12866 27056
rect 12860 27016 13033 27044
rect 12860 27004 12866 27016
rect 11348 26948 12204 26976
rect 11790 26908 11796 26920
rect 10888 26880 11796 26908
rect 11790 26868 11796 26880
rect 11848 26908 11854 26920
rect 12176 26917 12204 26948
rect 12894 26936 12900 26988
rect 12952 26936 12958 26988
rect 13005 26985 13033 27016
rect 13078 27004 13084 27056
rect 13136 27044 13142 27056
rect 13173 27047 13231 27053
rect 13173 27044 13185 27047
rect 13136 27016 13185 27044
rect 13136 27004 13142 27016
rect 13173 27013 13185 27016
rect 13219 27013 13231 27047
rect 13173 27007 13231 27013
rect 13906 27004 13912 27056
rect 13964 27044 13970 27056
rect 13964 27016 15148 27044
rect 13964 27004 13970 27016
rect 12990 26979 13048 26985
rect 12990 26945 13002 26979
rect 13036 26945 13048 26979
rect 12990 26939 13048 26945
rect 13262 26936 13268 26988
rect 13320 26936 13326 26988
rect 13354 26936 13360 26988
rect 13412 26985 13418 26988
rect 13412 26976 13420 26985
rect 13538 26976 13544 26988
rect 13412 26948 13544 26976
rect 13412 26939 13420 26948
rect 13412 26936 13418 26939
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 13630 26936 13636 26988
rect 13688 26976 13694 26988
rect 15120 26985 15148 27016
rect 14645 26979 14703 26985
rect 14645 26976 14657 26979
rect 13688 26948 14657 26976
rect 13688 26936 13694 26948
rect 14645 26945 14657 26948
rect 14691 26945 14703 26979
rect 14645 26939 14703 26945
rect 15013 26979 15071 26985
rect 15013 26945 15025 26979
rect 15059 26945 15071 26979
rect 15013 26939 15071 26945
rect 15105 26979 15163 26985
rect 15105 26945 15117 26979
rect 15151 26945 15163 26979
rect 15212 26976 15240 27072
rect 16114 27044 16120 27056
rect 15764 27016 16120 27044
rect 15473 26979 15531 26985
rect 15473 26976 15485 26979
rect 15212 26948 15485 26976
rect 15105 26939 15163 26945
rect 15473 26945 15485 26948
rect 15519 26945 15531 26979
rect 15473 26939 15531 26945
rect 11977 26911 12035 26917
rect 11977 26908 11989 26911
rect 11848 26880 11989 26908
rect 11848 26868 11854 26880
rect 11977 26877 11989 26880
rect 12023 26877 12035 26911
rect 11977 26871 12035 26877
rect 12161 26911 12219 26917
rect 12161 26877 12173 26911
rect 12207 26908 12219 26911
rect 14182 26908 14188 26920
rect 12207 26880 14188 26908
rect 12207 26877 12219 26880
rect 12161 26871 12219 26877
rect 14182 26868 14188 26880
rect 14240 26868 14246 26920
rect 14461 26911 14519 26917
rect 14461 26877 14473 26911
rect 14507 26877 14519 26911
rect 15028 26908 15056 26939
rect 15654 26936 15660 26988
rect 15712 26936 15718 26988
rect 15764 26985 15792 27016
rect 16114 27004 16120 27016
rect 16172 27004 16178 27056
rect 16868 27044 16896 27072
rect 16868 27016 17080 27044
rect 15749 26979 15807 26985
rect 15749 26945 15761 26979
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 15933 26979 15991 26985
rect 15933 26976 15945 26979
rect 15896 26948 15945 26976
rect 15896 26936 15902 26948
rect 15933 26945 15945 26948
rect 15979 26945 15991 26979
rect 15933 26939 15991 26945
rect 16022 26936 16028 26988
rect 16080 26936 16086 26988
rect 16758 26936 16764 26988
rect 16816 26976 16822 26988
rect 17052 26985 17080 27016
rect 17236 26985 17264 27084
rect 18138 27072 18144 27124
rect 18196 27112 18202 27124
rect 18196 27084 19288 27112
rect 18196 27072 18202 27084
rect 17589 27047 17647 27053
rect 17589 27013 17601 27047
rect 17635 27044 17647 27047
rect 17635 27016 18920 27044
rect 17635 27013 17647 27016
rect 17589 27007 17647 27013
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16816 26948 16865 26976
rect 16816 26936 16822 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 17037 26979 17095 26985
rect 17037 26945 17049 26979
rect 17083 26945 17095 26979
rect 17037 26939 17095 26945
rect 17221 26979 17279 26985
rect 17221 26945 17233 26979
rect 17267 26945 17279 26979
rect 17221 26939 17279 26945
rect 17405 26979 17463 26985
rect 17405 26945 17417 26979
rect 17451 26945 17463 26979
rect 17405 26939 17463 26945
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 15289 26911 15347 26917
rect 15289 26908 15301 26911
rect 15028 26880 15301 26908
rect 14461 26871 14519 26877
rect 15289 26877 15301 26880
rect 15335 26877 15347 26911
rect 16040 26908 16068 26936
rect 17129 26911 17187 26917
rect 17129 26908 17141 26911
rect 16040 26880 17141 26908
rect 15289 26871 15347 26877
rect 17129 26877 17141 26880
rect 17175 26908 17187 26911
rect 17420 26908 17448 26939
rect 17175 26880 17448 26908
rect 18156 26908 18184 26939
rect 18322 26936 18328 26988
rect 18380 26936 18386 26988
rect 18414 26936 18420 26988
rect 18472 26936 18478 26988
rect 18509 26979 18567 26985
rect 18509 26945 18521 26979
rect 18555 26976 18567 26979
rect 18690 26976 18696 26988
rect 18555 26948 18696 26976
rect 18555 26945 18567 26948
rect 18509 26939 18567 26945
rect 18690 26936 18696 26948
rect 18748 26936 18754 26988
rect 18782 26936 18788 26988
rect 18840 26936 18846 26988
rect 18892 26974 18920 27016
rect 19058 27004 19064 27056
rect 19116 27004 19122 27056
rect 18969 26979 19027 26985
rect 18969 26974 18981 26979
rect 18892 26946 18981 26974
rect 18969 26945 18981 26946
rect 19015 26945 19027 26979
rect 19153 26979 19211 26985
rect 19153 26960 19165 26979
rect 18969 26939 19027 26945
rect 19076 26945 19165 26960
rect 19199 26945 19211 26979
rect 19260 26976 19288 27084
rect 20714 27072 20720 27124
rect 20772 27112 20778 27124
rect 23750 27112 23756 27124
rect 20772 27084 23756 27112
rect 20772 27072 20778 27084
rect 23750 27072 23756 27084
rect 23808 27072 23814 27124
rect 25866 27072 25872 27124
rect 25924 27072 25930 27124
rect 26421 27115 26479 27121
rect 26421 27081 26433 27115
rect 26467 27112 26479 27115
rect 29546 27112 29552 27124
rect 26467 27084 29552 27112
rect 26467 27081 26479 27084
rect 26421 27075 26479 27081
rect 29546 27072 29552 27084
rect 29604 27072 29610 27124
rect 34698 27072 34704 27124
rect 34756 27072 34762 27124
rect 34790 27072 34796 27124
rect 34848 27112 34854 27124
rect 35342 27112 35348 27124
rect 34848 27084 35348 27112
rect 34848 27072 34854 27084
rect 35342 27072 35348 27084
rect 35400 27072 35406 27124
rect 20990 27004 20996 27056
rect 21048 27044 21054 27056
rect 24394 27044 24400 27056
rect 21048 27016 24400 27044
rect 21048 27004 21054 27016
rect 24394 27004 24400 27016
rect 24452 27004 24458 27056
rect 24854 27004 24860 27056
rect 24912 27044 24918 27056
rect 25884 27044 25912 27072
rect 24912 27016 26004 27044
rect 24912 27004 24918 27016
rect 25590 26976 25596 26988
rect 19260 26948 25596 26976
rect 19076 26939 19211 26945
rect 19076 26932 19196 26939
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 25774 26936 25780 26988
rect 25832 26936 25838 26988
rect 25976 26985 26004 27016
rect 27798 27004 27804 27056
rect 27856 27044 27862 27056
rect 28534 27044 28540 27056
rect 27856 27016 28540 27044
rect 27856 27004 27862 27016
rect 28534 27004 28540 27016
rect 28592 27044 28598 27056
rect 28592 27016 29040 27044
rect 28592 27004 28598 27016
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26945 25927 26979
rect 25869 26939 25927 26945
rect 25961 26979 26019 26985
rect 25961 26945 25973 26979
rect 26007 26945 26019 26979
rect 25961 26939 26019 26945
rect 18156 26880 19012 26908
rect 17175 26877 17187 26880
rect 17129 26871 17187 26877
rect 13541 26843 13599 26849
rect 10428 26812 12388 26840
rect 7800 26744 9444 26772
rect 9861 26775 9919 26781
rect 7800 26732 7806 26744
rect 9861 26741 9873 26775
rect 9907 26772 9919 26775
rect 10428 26772 10456 26812
rect 9907 26744 10456 26772
rect 9907 26741 9919 26744
rect 9861 26735 9919 26741
rect 10594 26732 10600 26784
rect 10652 26772 10658 26784
rect 10781 26775 10839 26781
rect 10781 26772 10793 26775
rect 10652 26744 10793 26772
rect 10652 26732 10658 26744
rect 10781 26741 10793 26744
rect 10827 26741 10839 26775
rect 10781 26735 10839 26741
rect 10962 26732 10968 26784
rect 11020 26772 11026 26784
rect 12250 26772 12256 26784
rect 11020 26744 12256 26772
rect 11020 26732 11026 26744
rect 12250 26732 12256 26744
rect 12308 26732 12314 26784
rect 12360 26772 12388 26812
rect 13541 26809 13553 26843
rect 13587 26840 13599 26843
rect 14476 26840 14504 26871
rect 18984 26852 19012 26880
rect 19076 26852 19104 26932
rect 25884 26908 25912 26939
rect 26050 26936 26056 26988
rect 26108 26976 26114 26988
rect 26237 26979 26295 26985
rect 26237 26976 26249 26979
rect 26108 26948 26249 26976
rect 26108 26936 26114 26948
rect 26237 26945 26249 26948
rect 26283 26945 26295 26979
rect 26237 26939 26295 26945
rect 27614 26936 27620 26988
rect 27672 26936 27678 26988
rect 28626 26936 28632 26988
rect 28684 26936 28690 26988
rect 28718 26936 28724 26988
rect 28776 26976 28782 26988
rect 28776 26948 28821 26976
rect 28776 26936 28782 26948
rect 28902 26936 28908 26988
rect 28960 26936 28966 26988
rect 29012 26985 29040 27016
rect 28997 26979 29055 26985
rect 28997 26945 29009 26979
rect 29043 26945 29055 26979
rect 28997 26939 29055 26945
rect 29135 26979 29193 26985
rect 29135 26945 29147 26979
rect 29181 26976 29193 26979
rect 30098 26976 30104 26988
rect 29181 26948 30104 26976
rect 29181 26945 29193 26948
rect 29135 26939 29193 26945
rect 30098 26936 30104 26948
rect 30156 26936 30162 26988
rect 30742 26936 30748 26988
rect 30800 26976 30806 26988
rect 31018 26976 31024 26988
rect 30800 26948 31024 26976
rect 30800 26936 30806 26948
rect 31018 26936 31024 26948
rect 31076 26936 31082 26988
rect 34330 26936 34336 26988
rect 34388 26936 34394 26988
rect 34716 26976 34744 27072
rect 34793 26979 34851 26985
rect 34793 26976 34805 26979
rect 34716 26948 34805 26976
rect 34793 26945 34805 26948
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 30282 26908 30288 26920
rect 19276 26880 30288 26908
rect 13587 26812 14504 26840
rect 15565 26843 15623 26849
rect 13587 26809 13599 26812
rect 13541 26803 13599 26809
rect 15565 26809 15577 26843
rect 15611 26809 15623 26843
rect 18693 26843 18751 26849
rect 18693 26840 18705 26843
rect 15565 26803 15623 26809
rect 15856 26812 18705 26840
rect 13814 26772 13820 26784
rect 12360 26744 13820 26772
rect 13814 26732 13820 26744
rect 13872 26732 13878 26784
rect 14277 26775 14335 26781
rect 14277 26741 14289 26775
rect 14323 26772 14335 26775
rect 14550 26772 14556 26784
rect 14323 26744 14556 26772
rect 14323 26741 14335 26744
rect 14277 26735 14335 26741
rect 14550 26732 14556 26744
rect 14608 26732 14614 26784
rect 15580 26772 15608 26803
rect 15856 26772 15884 26812
rect 18693 26809 18705 26812
rect 18739 26809 18751 26843
rect 18693 26803 18751 26809
rect 18874 26800 18880 26852
rect 18932 26800 18938 26852
rect 18966 26800 18972 26852
rect 19024 26800 19030 26852
rect 19058 26800 19064 26852
rect 19116 26800 19122 26852
rect 19276 26840 19304 26880
rect 30282 26868 30288 26880
rect 30340 26908 30346 26920
rect 30340 26880 31754 26908
rect 30340 26868 30346 26880
rect 19260 26812 19304 26840
rect 15580 26744 15884 26772
rect 16482 26732 16488 26784
rect 16540 26772 16546 26784
rect 18892 26772 18920 26800
rect 16540 26744 18920 26772
rect 18984 26772 19012 26800
rect 19260 26772 19288 26812
rect 24118 26800 24124 26852
rect 24176 26840 24182 26852
rect 31294 26840 31300 26852
rect 24176 26812 31300 26840
rect 24176 26800 24182 26812
rect 31294 26800 31300 26812
rect 31352 26800 31358 26852
rect 18984 26744 19288 26772
rect 16540 26732 16546 26744
rect 19334 26732 19340 26784
rect 19392 26732 19398 26784
rect 21818 26732 21824 26784
rect 21876 26772 21882 26784
rect 22278 26772 22284 26784
rect 21876 26744 22284 26772
rect 21876 26732 21882 26744
rect 22278 26732 22284 26744
rect 22336 26772 22342 26784
rect 25590 26772 25596 26784
rect 22336 26744 25596 26772
rect 22336 26732 22342 26744
rect 25590 26732 25596 26744
rect 25648 26732 25654 26784
rect 26142 26732 26148 26784
rect 26200 26732 26206 26784
rect 27430 26732 27436 26784
rect 27488 26732 27494 26784
rect 29270 26732 29276 26784
rect 29328 26732 29334 26784
rect 31726 26772 31754 26880
rect 32582 26772 32588 26784
rect 31726 26744 32588 26772
rect 32582 26732 32588 26744
rect 32640 26732 32646 26784
rect 34149 26775 34207 26781
rect 34149 26741 34161 26775
rect 34195 26772 34207 26775
rect 34606 26772 34612 26784
rect 34195 26744 34612 26772
rect 34195 26741 34207 26744
rect 34149 26735 34207 26741
rect 34606 26732 34612 26744
rect 34664 26732 34670 26784
rect 34790 26732 34796 26784
rect 34848 26772 34854 26784
rect 34885 26775 34943 26781
rect 34885 26772 34897 26775
rect 34848 26744 34897 26772
rect 34848 26732 34854 26744
rect 34885 26741 34897 26744
rect 34931 26741 34943 26775
rect 34885 26735 34943 26741
rect 1104 26682 38272 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38272 26682
rect 1104 26608 38272 26630
rect 5350 26528 5356 26580
rect 5408 26568 5414 26580
rect 10492 26571 10550 26577
rect 5408 26540 9996 26568
rect 5408 26528 5414 26540
rect 8386 26460 8392 26512
rect 8444 26500 8450 26512
rect 8941 26503 8999 26509
rect 8941 26500 8953 26503
rect 8444 26472 8953 26500
rect 8444 26460 8450 26472
rect 8941 26469 8953 26472
rect 8987 26469 8999 26503
rect 8941 26463 8999 26469
rect 9490 26460 9496 26512
rect 9548 26460 9554 26512
rect 4062 26392 4068 26444
rect 4120 26432 4126 26444
rect 7098 26432 7104 26444
rect 4120 26404 7104 26432
rect 4120 26392 4126 26404
rect 7098 26392 7104 26404
rect 7156 26392 7162 26444
rect 8662 26392 8668 26444
rect 8720 26392 8726 26444
rect 4801 26367 4859 26373
rect 4801 26333 4813 26367
rect 4847 26333 4859 26367
rect 4801 26327 4859 26333
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26364 4951 26367
rect 5077 26367 5135 26373
rect 5077 26364 5089 26367
rect 4939 26336 5089 26364
rect 4939 26333 4951 26336
rect 4893 26327 4951 26333
rect 5077 26333 5089 26336
rect 5123 26333 5135 26367
rect 6638 26364 6644 26376
rect 6486 26336 6644 26364
rect 5077 26327 5135 26333
rect 4816 26296 4844 26327
rect 6638 26324 6644 26336
rect 6696 26364 6702 26376
rect 8680 26364 8708 26392
rect 6696 26336 8708 26364
rect 6696 26324 6702 26336
rect 5258 26296 5264 26308
rect 4816 26268 5264 26296
rect 5258 26256 5264 26268
rect 5316 26256 5322 26308
rect 5353 26299 5411 26305
rect 5353 26265 5365 26299
rect 5399 26296 5411 26299
rect 5442 26296 5448 26308
rect 5399 26268 5448 26296
rect 5399 26265 5411 26268
rect 5353 26259 5411 26265
rect 5442 26256 5448 26268
rect 5500 26256 5506 26308
rect 7101 26299 7159 26305
rect 7101 26265 7113 26299
rect 7147 26296 7159 26299
rect 7190 26296 7196 26308
rect 7147 26268 7196 26296
rect 7147 26265 7159 26268
rect 7101 26259 7159 26265
rect 7190 26256 7196 26268
rect 7248 26256 7254 26308
rect 8680 26296 8708 26336
rect 9125 26367 9183 26373
rect 9125 26333 9137 26367
rect 9171 26364 9183 26367
rect 9508 26364 9536 26460
rect 9968 26432 9996 26540
rect 10492 26537 10504 26571
rect 10538 26568 10550 26571
rect 10594 26568 10600 26580
rect 10538 26540 10600 26568
rect 10538 26537 10550 26540
rect 10492 26531 10550 26537
rect 10594 26528 10600 26540
rect 10652 26528 10658 26580
rect 11974 26528 11980 26580
rect 12032 26528 12038 26580
rect 12158 26528 12164 26580
rect 12216 26528 12222 26580
rect 12894 26528 12900 26580
rect 12952 26568 12958 26580
rect 17865 26571 17923 26577
rect 12952 26540 15700 26568
rect 12952 26528 12958 26540
rect 12176 26432 12204 26528
rect 15672 26512 15700 26540
rect 17865 26537 17877 26571
rect 17911 26568 17923 26571
rect 19334 26568 19340 26580
rect 17911 26540 19340 26568
rect 17911 26537 17923 26540
rect 17865 26531 17923 26537
rect 19334 26528 19340 26540
rect 19392 26528 19398 26580
rect 21821 26571 21879 26577
rect 21821 26568 21833 26571
rect 21100 26540 21833 26568
rect 14182 26460 14188 26512
rect 14240 26460 14246 26512
rect 15654 26460 15660 26512
rect 15712 26460 15718 26512
rect 17681 26503 17739 26509
rect 17681 26469 17693 26503
rect 17727 26500 17739 26503
rect 17727 26472 17908 26500
rect 17727 26469 17739 26472
rect 17681 26463 17739 26469
rect 9968 26404 12204 26432
rect 9968 26373 9996 26404
rect 13262 26392 13268 26444
rect 13320 26432 13326 26444
rect 17880 26441 17908 26472
rect 17865 26435 17923 26441
rect 13320 26404 17448 26432
rect 13320 26392 13326 26404
rect 9171 26336 9536 26364
rect 9953 26367 10011 26373
rect 9171 26333 9183 26336
rect 9125 26327 9183 26333
rect 9953 26333 9965 26367
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 10045 26367 10103 26373
rect 10045 26333 10057 26367
rect 10091 26364 10103 26367
rect 10229 26367 10287 26373
rect 10229 26364 10241 26367
rect 10091 26336 10241 26364
rect 10091 26333 10103 26336
rect 10045 26327 10103 26333
rect 10229 26333 10241 26336
rect 10275 26333 10287 26367
rect 10229 26327 10287 26333
rect 14090 26324 14096 26376
rect 14148 26324 14154 26376
rect 14642 26324 14648 26376
rect 14700 26324 14706 26376
rect 14918 26324 14924 26376
rect 14976 26324 14982 26376
rect 16390 26324 16396 26376
rect 16448 26324 16454 26376
rect 16574 26324 16580 26376
rect 16632 26324 16638 26376
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26364 16819 26367
rect 17037 26367 17095 26373
rect 17037 26364 17049 26367
rect 16807 26336 17049 26364
rect 16807 26333 16819 26336
rect 16761 26327 16819 26333
rect 17037 26333 17049 26336
rect 17083 26333 17095 26367
rect 17037 26327 17095 26333
rect 17126 26324 17132 26376
rect 17184 26324 17190 26376
rect 17310 26324 17316 26376
rect 17368 26324 17374 26376
rect 10962 26296 10968 26308
rect 8680 26268 10968 26296
rect 10962 26256 10968 26268
rect 11020 26256 11026 26308
rect 14936 26296 14964 26324
rect 13740 26268 14964 26296
rect 8938 26188 8944 26240
rect 8996 26228 9002 26240
rect 13078 26228 13084 26240
rect 8996 26200 13084 26228
rect 8996 26188 9002 26200
rect 13078 26188 13084 26200
rect 13136 26188 13142 26240
rect 13354 26188 13360 26240
rect 13412 26228 13418 26240
rect 13740 26228 13768 26268
rect 15746 26256 15752 26308
rect 15804 26296 15810 26308
rect 17420 26305 17448 26404
rect 17865 26401 17877 26435
rect 17911 26401 17923 26435
rect 17865 26395 17923 26401
rect 18782 26392 18788 26444
rect 18840 26392 18846 26444
rect 17543 26367 17601 26373
rect 17543 26333 17555 26367
rect 17589 26364 17601 26367
rect 17678 26364 17684 26376
rect 17589 26336 17684 26364
rect 17589 26333 17601 26336
rect 17543 26327 17601 26333
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 17770 26324 17776 26376
rect 17828 26324 17834 26376
rect 18414 26364 18420 26376
rect 17972 26336 18420 26364
rect 16209 26299 16267 26305
rect 16209 26296 16221 26299
rect 15804 26268 16221 26296
rect 15804 26256 15810 26268
rect 16209 26265 16221 26268
rect 16255 26296 16267 26299
rect 17405 26299 17463 26305
rect 16255 26268 16620 26296
rect 16255 26265 16267 26268
rect 16209 26259 16267 26265
rect 13412 26200 13768 26228
rect 13412 26188 13418 26200
rect 16298 26188 16304 26240
rect 16356 26228 16362 26240
rect 16485 26231 16543 26237
rect 16485 26228 16497 26231
rect 16356 26200 16497 26228
rect 16356 26188 16362 26200
rect 16485 26197 16497 26200
rect 16531 26197 16543 26231
rect 16592 26228 16620 26268
rect 17405 26265 17417 26299
rect 17451 26296 17463 26299
rect 17972 26296 18000 26336
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 18800 26364 18828 26392
rect 20809 26367 20867 26373
rect 20809 26364 20821 26367
rect 18800 26336 20821 26364
rect 20809 26333 20821 26336
rect 20855 26364 20867 26367
rect 20898 26364 20904 26376
rect 20855 26336 20904 26364
rect 20855 26333 20867 26336
rect 20809 26327 20867 26333
rect 20898 26324 20904 26336
rect 20956 26324 20962 26376
rect 20993 26367 21051 26373
rect 20993 26333 21005 26367
rect 21039 26364 21051 26367
rect 21100 26364 21128 26540
rect 21821 26537 21833 26540
rect 21867 26537 21879 26571
rect 21821 26531 21879 26537
rect 22186 26528 22192 26580
rect 22244 26568 22250 26580
rect 29917 26571 29975 26577
rect 22244 26540 28994 26568
rect 22244 26528 22250 26540
rect 22462 26460 22468 26512
rect 22520 26500 22526 26512
rect 22738 26500 22744 26512
rect 22520 26472 22744 26500
rect 22520 26460 22526 26472
rect 22738 26460 22744 26472
rect 22796 26460 22802 26512
rect 21450 26392 21456 26444
rect 21508 26432 21514 26444
rect 21508 26404 21772 26432
rect 21508 26392 21514 26404
rect 21039 26336 21128 26364
rect 21039 26333 21051 26336
rect 20993 26327 21051 26333
rect 21174 26324 21180 26376
rect 21232 26324 21238 26376
rect 17451 26268 18000 26296
rect 18064 26268 18276 26296
rect 17451 26265 17463 26268
rect 17405 26259 17463 26265
rect 18064 26228 18092 26268
rect 16592 26200 18092 26228
rect 16485 26191 16543 26197
rect 18138 26188 18144 26240
rect 18196 26188 18202 26240
rect 18248 26228 18276 26268
rect 18874 26256 18880 26308
rect 18932 26296 18938 26308
rect 20070 26296 20076 26308
rect 18932 26268 20076 26296
rect 18932 26256 18938 26268
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 20530 26256 20536 26308
rect 20588 26296 20594 26308
rect 21077 26299 21135 26305
rect 21077 26296 21089 26299
rect 20588 26268 21089 26296
rect 20588 26256 20594 26268
rect 21077 26265 21089 26268
rect 21123 26265 21135 26299
rect 21077 26259 21135 26265
rect 21453 26299 21511 26305
rect 21453 26265 21465 26299
rect 21499 26296 21511 26299
rect 21542 26296 21548 26308
rect 21499 26268 21548 26296
rect 21499 26265 21511 26268
rect 21453 26259 21511 26265
rect 21542 26256 21548 26268
rect 21600 26256 21606 26308
rect 21637 26299 21695 26305
rect 21637 26265 21649 26299
rect 21683 26296 21695 26299
rect 21744 26296 21772 26404
rect 25866 26392 25872 26444
rect 25924 26432 25930 26444
rect 25924 26404 26280 26432
rect 25924 26392 25930 26404
rect 23290 26324 23296 26376
rect 23348 26364 23354 26376
rect 23842 26364 23848 26376
rect 23348 26336 23848 26364
rect 23348 26324 23354 26336
rect 23842 26324 23848 26336
rect 23900 26324 23906 26376
rect 24026 26324 24032 26376
rect 24084 26324 24090 26376
rect 24121 26367 24179 26373
rect 24121 26333 24133 26367
rect 24167 26364 24179 26367
rect 24397 26367 24455 26373
rect 24397 26364 24409 26367
rect 24167 26336 24409 26364
rect 24167 26333 24179 26336
rect 24121 26327 24179 26333
rect 24397 26333 24409 26336
rect 24443 26333 24455 26367
rect 24397 26327 24455 26333
rect 21683 26268 21772 26296
rect 21683 26265 21695 26268
rect 21637 26259 21695 26265
rect 24670 26256 24676 26308
rect 24728 26256 24734 26308
rect 25406 26256 25412 26308
rect 25464 26256 25470 26308
rect 20806 26228 20812 26240
rect 18248 26200 20812 26228
rect 20806 26188 20812 26200
rect 20864 26188 20870 26240
rect 21361 26231 21419 26237
rect 21361 26197 21373 26231
rect 21407 26228 21419 26231
rect 22554 26228 22560 26240
rect 21407 26200 22560 26228
rect 21407 26197 21419 26200
rect 21361 26191 21419 26197
rect 22554 26188 22560 26200
rect 22612 26188 22618 26240
rect 25498 26188 25504 26240
rect 25556 26228 25562 26240
rect 26145 26231 26203 26237
rect 26145 26228 26157 26231
rect 25556 26200 26157 26228
rect 25556 26188 25562 26200
rect 26145 26197 26157 26200
rect 26191 26197 26203 26231
rect 26252 26228 26280 26404
rect 26436 26364 26464 26540
rect 26510 26460 26516 26512
rect 26568 26460 26574 26512
rect 26694 26460 26700 26512
rect 26752 26500 26758 26512
rect 26752 26472 26924 26500
rect 26752 26460 26758 26472
rect 26528 26432 26556 26460
rect 26528 26404 26740 26432
rect 26712 26373 26740 26404
rect 26605 26367 26663 26373
rect 26605 26364 26617 26367
rect 26436 26336 26617 26364
rect 26605 26333 26617 26336
rect 26651 26333 26663 26367
rect 26605 26327 26663 26333
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26333 26755 26367
rect 26697 26327 26755 26333
rect 26789 26367 26847 26373
rect 26789 26333 26801 26367
rect 26835 26333 26847 26367
rect 26896 26364 26924 26472
rect 27341 26435 27399 26441
rect 27341 26401 27353 26435
rect 27387 26432 27399 26435
rect 27430 26432 27436 26444
rect 27387 26404 27436 26432
rect 27387 26401 27399 26404
rect 27341 26395 27399 26401
rect 27430 26392 27436 26404
rect 27488 26392 27494 26444
rect 28966 26432 28994 26540
rect 29917 26537 29929 26571
rect 29963 26568 29975 26571
rect 33321 26571 33379 26577
rect 29963 26540 31156 26568
rect 29963 26537 29975 26540
rect 29917 26531 29975 26537
rect 30561 26503 30619 26509
rect 30561 26469 30573 26503
rect 30607 26500 30619 26503
rect 30650 26500 30656 26512
rect 30607 26472 30656 26500
rect 30607 26469 30619 26472
rect 30561 26463 30619 26469
rect 30650 26460 30656 26472
rect 30708 26460 30714 26512
rect 28966 26404 30604 26432
rect 26973 26367 27031 26373
rect 26973 26364 26985 26367
rect 26896 26336 26985 26364
rect 26789 26327 26847 26333
rect 26973 26333 26985 26336
rect 27019 26333 27031 26367
rect 26973 26327 27031 26333
rect 26326 26256 26332 26308
rect 26384 26256 26390 26308
rect 26804 26228 26832 26327
rect 27062 26324 27068 26376
rect 27120 26324 27126 26376
rect 29086 26324 29092 26376
rect 29144 26364 29150 26376
rect 29181 26367 29239 26373
rect 29181 26364 29193 26367
rect 29144 26336 29193 26364
rect 29144 26324 29150 26336
rect 29181 26333 29193 26336
rect 29227 26333 29239 26367
rect 29181 26327 29239 26333
rect 29270 26324 29276 26376
rect 29328 26364 29334 26376
rect 30101 26367 30159 26373
rect 30101 26364 30113 26367
rect 29328 26336 30113 26364
rect 29328 26324 29334 26336
rect 30101 26333 30113 26336
rect 30147 26333 30159 26367
rect 30101 26327 30159 26333
rect 30282 26324 30288 26376
rect 30340 26324 30346 26376
rect 30377 26367 30435 26373
rect 30377 26333 30389 26367
rect 30423 26364 30435 26367
rect 30466 26364 30472 26376
rect 30423 26336 30472 26364
rect 30423 26333 30435 26336
rect 30377 26327 30435 26333
rect 30466 26324 30472 26336
rect 30524 26324 30530 26376
rect 30576 26364 30604 26404
rect 30742 26364 30748 26376
rect 30576 26336 30748 26364
rect 30742 26324 30748 26336
rect 30800 26366 30806 26376
rect 30837 26367 30895 26373
rect 30837 26366 30849 26367
rect 30800 26338 30849 26366
rect 30800 26324 30806 26338
rect 30837 26333 30849 26338
rect 30883 26333 30895 26367
rect 30837 26327 30895 26333
rect 30929 26367 30987 26373
rect 30929 26333 30941 26367
rect 30975 26333 30987 26367
rect 30929 26327 30987 26333
rect 27798 26256 27804 26308
rect 27856 26256 27862 26308
rect 30944 26296 30972 26327
rect 31018 26324 31024 26376
rect 31076 26324 31082 26376
rect 31128 26364 31156 26540
rect 33321 26537 33333 26571
rect 33367 26568 33379 26571
rect 34330 26568 34336 26580
rect 33367 26540 34336 26568
rect 33367 26537 33379 26540
rect 33321 26531 33379 26537
rect 34330 26528 34336 26540
rect 34388 26528 34394 26580
rect 34698 26528 34704 26580
rect 34756 26528 34762 26580
rect 34790 26528 34796 26580
rect 34848 26528 34854 26580
rect 32674 26460 32680 26512
rect 32732 26500 32738 26512
rect 33137 26503 33195 26509
rect 33137 26500 33149 26503
rect 32732 26472 33149 26500
rect 32732 26460 32738 26472
rect 33137 26469 33149 26472
rect 33183 26469 33195 26503
rect 34716 26500 34744 26528
rect 33137 26463 33195 26469
rect 34348 26472 34744 26500
rect 33778 26392 33784 26444
rect 33836 26432 33842 26444
rect 33873 26435 33931 26441
rect 33873 26432 33885 26435
rect 33836 26404 33885 26432
rect 33836 26392 33842 26404
rect 33873 26401 33885 26404
rect 33919 26432 33931 26435
rect 34238 26432 34244 26444
rect 33919 26404 34244 26432
rect 33919 26401 33931 26404
rect 33873 26395 33931 26401
rect 34238 26392 34244 26404
rect 34296 26392 34302 26444
rect 31205 26367 31263 26373
rect 31205 26364 31217 26367
rect 31128 26336 31217 26364
rect 31205 26333 31217 26336
rect 31251 26333 31263 26367
rect 31205 26327 31263 26333
rect 31386 26324 31392 26376
rect 31444 26324 31450 26376
rect 34348 26373 34376 26472
rect 34606 26392 34612 26444
rect 34664 26392 34670 26444
rect 34701 26435 34759 26441
rect 34701 26401 34713 26435
rect 34747 26432 34759 26435
rect 34808 26432 34836 26528
rect 34747 26404 34836 26432
rect 34747 26401 34759 26404
rect 34701 26395 34759 26401
rect 34333 26367 34391 26373
rect 34333 26333 34345 26367
rect 34379 26333 34391 26367
rect 34333 26327 34391 26333
rect 30944 26268 31248 26296
rect 26252 26200 26832 26228
rect 26145 26191 26203 26197
rect 28350 26188 28356 26240
rect 28408 26228 28414 26240
rect 28718 26228 28724 26240
rect 28408 26200 28724 26228
rect 28408 26188 28414 26200
rect 28718 26188 28724 26200
rect 28776 26228 28782 26240
rect 28813 26231 28871 26237
rect 28813 26228 28825 26231
rect 28776 26200 28825 26228
rect 28776 26188 28782 26200
rect 28813 26197 28825 26200
rect 28859 26197 28871 26231
rect 28813 26191 28871 26197
rect 29086 26188 29092 26240
rect 29144 26228 29150 26240
rect 29273 26231 29331 26237
rect 29273 26228 29285 26231
rect 29144 26200 29285 26228
rect 29144 26188 29150 26200
rect 29273 26197 29285 26200
rect 29319 26197 29331 26231
rect 29273 26191 29331 26197
rect 30558 26188 30564 26240
rect 30616 26228 30622 26240
rect 30944 26228 30972 26268
rect 31220 26240 31248 26268
rect 31294 26256 31300 26308
rect 31352 26256 31358 26308
rect 31665 26299 31723 26305
rect 31665 26265 31677 26299
rect 31711 26296 31723 26299
rect 31754 26296 31760 26308
rect 31711 26268 31760 26296
rect 31711 26265 31723 26268
rect 31665 26259 31723 26265
rect 31754 26256 31760 26268
rect 31812 26256 31818 26308
rect 32048 26268 32154 26296
rect 30616 26200 30972 26228
rect 30616 26188 30622 26200
rect 31202 26188 31208 26240
rect 31260 26188 31266 26240
rect 31312 26228 31340 26256
rect 32048 26228 32076 26268
rect 33686 26256 33692 26308
rect 33744 26296 33750 26308
rect 34624 26296 34652 26392
rect 34977 26299 35035 26305
rect 34977 26296 34989 26299
rect 33744 26268 34560 26296
rect 34624 26268 34989 26296
rect 33744 26256 33750 26268
rect 31312 26200 32076 26228
rect 32490 26188 32496 26240
rect 32548 26228 32554 26240
rect 33781 26231 33839 26237
rect 33781 26228 33793 26231
rect 32548 26200 33793 26228
rect 32548 26188 32554 26200
rect 33781 26197 33793 26200
rect 33827 26197 33839 26231
rect 33781 26191 33839 26197
rect 34330 26188 34336 26240
rect 34388 26228 34394 26240
rect 34425 26231 34483 26237
rect 34425 26228 34437 26231
rect 34388 26200 34437 26228
rect 34388 26188 34394 26200
rect 34425 26197 34437 26200
rect 34471 26197 34483 26231
rect 34532 26228 34560 26268
rect 34977 26265 34989 26268
rect 35023 26265 35035 26299
rect 34977 26259 35035 26265
rect 35434 26256 35440 26308
rect 35492 26256 35498 26308
rect 36538 26256 36544 26308
rect 36596 26296 36602 26308
rect 36725 26299 36783 26305
rect 36725 26296 36737 26299
rect 36596 26268 36737 26296
rect 36596 26256 36602 26268
rect 36725 26265 36737 26268
rect 36771 26265 36783 26299
rect 36725 26259 36783 26265
rect 36556 26228 36584 26256
rect 34532 26200 36584 26228
rect 34425 26191 34483 26197
rect 1104 26138 38272 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38272 26138
rect 1104 26064 38272 26086
rect 5902 25984 5908 26036
rect 5960 26024 5966 26036
rect 6457 26027 6515 26033
rect 6457 26024 6469 26027
rect 5960 25996 6469 26024
rect 5960 25984 5966 25996
rect 6457 25993 6469 25996
rect 6503 25993 6515 26027
rect 6457 25987 6515 25993
rect 11054 25984 11060 26036
rect 11112 26024 11118 26036
rect 12158 26024 12164 26036
rect 11112 25996 12164 26024
rect 11112 25984 11118 25996
rect 12158 25984 12164 25996
rect 12216 25984 12222 26036
rect 15378 26024 15384 26036
rect 12912 25996 15384 26024
rect 6825 25959 6883 25965
rect 6825 25925 6837 25959
rect 6871 25956 6883 25959
rect 7190 25956 7196 25968
rect 6871 25928 7196 25956
rect 6871 25925 6883 25928
rect 6825 25919 6883 25925
rect 7190 25916 7196 25928
rect 7248 25956 7254 25968
rect 12912 25956 12940 25996
rect 15378 25984 15384 25996
rect 15436 25984 15442 26036
rect 23198 26024 23204 26036
rect 15764 25996 23204 26024
rect 7248 25928 12940 25956
rect 12989 25959 13047 25965
rect 7248 25916 7254 25928
rect 12989 25925 13001 25959
rect 13035 25956 13047 25959
rect 13722 25956 13728 25968
rect 13035 25928 13728 25956
rect 13035 25925 13047 25928
rect 12989 25919 13047 25925
rect 13722 25916 13728 25928
rect 13780 25916 13786 25968
rect 15764 25965 15792 25996
rect 23198 25984 23204 25996
rect 23256 25984 23262 26036
rect 23474 25984 23480 26036
rect 23532 25984 23538 26036
rect 23845 26027 23903 26033
rect 23845 25993 23857 26027
rect 23891 26024 23903 26027
rect 24397 26027 24455 26033
rect 24397 26024 24409 26027
rect 23891 25996 24409 26024
rect 23891 25993 23903 25996
rect 23845 25987 23903 25993
rect 24397 25993 24409 25996
rect 24443 25993 24455 26027
rect 24397 25987 24455 25993
rect 24489 26027 24547 26033
rect 24489 25993 24501 26027
rect 24535 26024 24547 26027
rect 24670 26024 24676 26036
rect 24535 25996 24676 26024
rect 24535 25993 24547 25996
rect 24489 25987 24547 25993
rect 24670 25984 24676 25996
rect 24728 25984 24734 26036
rect 24946 25984 24952 26036
rect 25004 26024 25010 26036
rect 25130 26024 25136 26036
rect 25004 25996 25136 26024
rect 25004 25984 25010 25996
rect 25130 25984 25136 25996
rect 25188 25984 25194 26036
rect 25777 26027 25835 26033
rect 25777 25993 25789 26027
rect 25823 26024 25835 26027
rect 25866 26024 25872 26036
rect 25823 25996 25872 26024
rect 25823 25993 25835 25996
rect 25777 25987 25835 25993
rect 25866 25984 25872 25996
rect 25924 25984 25930 26036
rect 26234 26024 26240 26036
rect 25976 25996 26240 26024
rect 15749 25959 15807 25965
rect 15749 25925 15761 25959
rect 15795 25925 15807 25959
rect 15749 25919 15807 25925
rect 16132 25928 18368 25956
rect 16132 25900 16160 25928
rect 5994 25848 6000 25900
rect 6052 25848 6058 25900
rect 6840 25860 7052 25888
rect 6840 25832 6868 25860
rect 6822 25780 6828 25832
rect 6880 25780 6886 25832
rect 7024 25829 7052 25860
rect 10410 25848 10416 25900
rect 10468 25848 10474 25900
rect 11793 25891 11851 25897
rect 11793 25857 11805 25891
rect 11839 25857 11851 25891
rect 11793 25851 11851 25857
rect 6917 25823 6975 25829
rect 6917 25789 6929 25823
rect 6963 25789 6975 25823
rect 6917 25783 6975 25789
rect 7009 25823 7067 25829
rect 7009 25789 7021 25823
rect 7055 25789 7067 25823
rect 11808 25820 11836 25851
rect 11882 25848 11888 25900
rect 11940 25848 11946 25900
rect 14642 25848 14648 25900
rect 14700 25888 14706 25900
rect 15013 25891 15071 25897
rect 15013 25888 15025 25891
rect 14700 25860 15025 25888
rect 14700 25848 14706 25860
rect 15013 25857 15025 25860
rect 15059 25857 15071 25891
rect 15013 25851 15071 25857
rect 15102 25848 15108 25900
rect 15160 25888 15166 25900
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 15160 25860 15485 25888
rect 15160 25848 15166 25860
rect 15473 25857 15485 25860
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 16114 25848 16120 25900
rect 16172 25848 16178 25900
rect 18230 25888 18236 25900
rect 17972 25860 18236 25888
rect 17972 25832 18000 25860
rect 18230 25848 18236 25860
rect 18288 25848 18294 25900
rect 11808 25792 17264 25820
rect 7009 25783 7067 25789
rect 5626 25644 5632 25696
rect 5684 25684 5690 25696
rect 5813 25687 5871 25693
rect 5813 25684 5825 25687
rect 5684 25656 5825 25684
rect 5684 25644 5690 25656
rect 5813 25653 5825 25656
rect 5859 25653 5871 25687
rect 6932 25684 6960 25783
rect 9398 25712 9404 25764
rect 9456 25752 9462 25764
rect 9456 25724 12434 25752
rect 9456 25712 9462 25724
rect 7926 25684 7932 25696
rect 6932 25656 7932 25684
rect 5813 25647 5871 25653
rect 7926 25644 7932 25656
rect 7984 25644 7990 25696
rect 10042 25644 10048 25696
rect 10100 25684 10106 25696
rect 10229 25687 10287 25693
rect 10229 25684 10241 25687
rect 10100 25656 10241 25684
rect 10100 25644 10106 25656
rect 10229 25653 10241 25656
rect 10275 25653 10287 25687
rect 10229 25647 10287 25653
rect 12066 25644 12072 25696
rect 12124 25644 12130 25696
rect 12406 25684 12434 25724
rect 12618 25712 12624 25764
rect 12676 25752 12682 25764
rect 16022 25752 16028 25764
rect 12676 25724 16028 25752
rect 12676 25712 12682 25724
rect 16022 25712 16028 25724
rect 16080 25712 16086 25764
rect 17236 25752 17264 25792
rect 17954 25780 17960 25832
rect 18012 25780 18018 25832
rect 18340 25829 18368 25928
rect 20346 25916 20352 25968
rect 20404 25956 20410 25968
rect 20404 25928 20944 25956
rect 20404 25916 20410 25928
rect 20622 25848 20628 25900
rect 20680 25848 20686 25900
rect 20916 25897 20944 25928
rect 22738 25916 22744 25968
rect 22796 25956 22802 25968
rect 23017 25959 23075 25965
rect 23017 25956 23029 25959
rect 22796 25928 23029 25956
rect 22796 25916 22802 25928
rect 23017 25925 23029 25928
rect 23063 25925 23075 25959
rect 23492 25956 23520 25984
rect 25682 25956 25688 25968
rect 23492 25928 23980 25956
rect 23017 25919 23075 25925
rect 20901 25891 20959 25897
rect 20901 25857 20913 25891
rect 20947 25857 20959 25891
rect 20901 25851 20959 25857
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 21450 25888 21456 25900
rect 21232 25860 21456 25888
rect 21232 25848 21238 25860
rect 21450 25848 21456 25860
rect 21508 25848 21514 25900
rect 22186 25848 22192 25900
rect 22244 25848 22250 25900
rect 22373 25891 22431 25897
rect 22373 25886 22385 25891
rect 22297 25858 22385 25886
rect 18325 25823 18383 25829
rect 18325 25789 18337 25823
rect 18371 25820 18383 25823
rect 22204 25820 22232 25848
rect 18371 25792 22232 25820
rect 18371 25789 18383 25792
rect 18325 25783 18383 25789
rect 19702 25752 19708 25764
rect 17236 25724 19708 25752
rect 19702 25712 19708 25724
rect 19760 25712 19766 25764
rect 19978 25712 19984 25764
rect 20036 25752 20042 25764
rect 20622 25752 20628 25764
rect 20036 25724 20628 25752
rect 20036 25712 20042 25724
rect 20622 25712 20628 25724
rect 20680 25712 20686 25764
rect 14461 25687 14519 25693
rect 14461 25684 14473 25687
rect 12406 25656 14473 25684
rect 14461 25653 14473 25656
rect 14507 25684 14519 25687
rect 16574 25684 16580 25696
rect 14507 25656 16580 25684
rect 14507 25653 14519 25656
rect 14461 25647 14519 25653
rect 16574 25644 16580 25656
rect 16632 25644 16638 25696
rect 18417 25687 18475 25693
rect 18417 25653 18429 25687
rect 18463 25684 18475 25687
rect 18506 25684 18512 25696
rect 18463 25656 18512 25684
rect 18463 25653 18475 25656
rect 18417 25647 18475 25653
rect 18506 25644 18512 25656
rect 18564 25644 18570 25696
rect 18598 25644 18604 25696
rect 18656 25644 18662 25696
rect 20438 25644 20444 25696
rect 20496 25644 20502 25696
rect 20806 25644 20812 25696
rect 20864 25644 20870 25696
rect 22186 25644 22192 25696
rect 22244 25644 22250 25696
rect 22297 25684 22325 25858
rect 22373 25857 22385 25858
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 22554 25848 22560 25900
rect 22612 25848 22618 25900
rect 22649 25891 22707 25897
rect 22649 25857 22661 25891
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 22833 25892 22891 25897
rect 22833 25891 22896 25892
rect 22833 25857 22845 25891
rect 22879 25888 22896 25891
rect 22879 25860 22968 25888
rect 22879 25857 22891 25860
rect 22833 25851 22891 25857
rect 22462 25712 22468 25764
rect 22520 25712 22526 25764
rect 22664 25752 22692 25851
rect 22940 25820 22968 25860
rect 23106 25848 23112 25900
rect 23164 25848 23170 25900
rect 23201 25891 23259 25897
rect 23201 25857 23213 25891
rect 23247 25888 23259 25891
rect 23290 25888 23296 25900
rect 23247 25860 23296 25888
rect 23247 25857 23259 25860
rect 23201 25851 23259 25857
rect 23290 25848 23296 25860
rect 23348 25848 23354 25900
rect 23658 25848 23664 25900
rect 23716 25848 23722 25900
rect 23952 25897 23980 25928
rect 24044 25928 25688 25956
rect 24044 25897 24072 25928
rect 25682 25916 25688 25928
rect 25740 25916 25746 25968
rect 23937 25891 23995 25897
rect 23937 25857 23949 25891
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 24029 25891 24087 25897
rect 24029 25857 24041 25891
rect 24075 25857 24087 25891
rect 24029 25851 24087 25857
rect 22940 25792 23336 25820
rect 23308 25764 23336 25792
rect 23842 25780 23848 25832
rect 23900 25820 23906 25832
rect 24044 25820 24072 25851
rect 24670 25848 24676 25900
rect 24728 25848 24734 25900
rect 24762 25848 24768 25900
rect 24820 25848 24826 25900
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 25976 25897 26004 25996
rect 26234 25984 26240 25996
rect 26292 25984 26298 26036
rect 26602 25984 26608 26036
rect 26660 25984 26666 26036
rect 27062 25984 27068 26036
rect 27120 26024 27126 26036
rect 27249 26027 27307 26033
rect 27249 26024 27261 26027
rect 27120 25996 27261 26024
rect 27120 25984 27126 25996
rect 27249 25993 27261 25996
rect 27295 25993 27307 26027
rect 27249 25987 27307 25993
rect 27525 26027 27583 26033
rect 27525 25993 27537 26027
rect 27571 26024 27583 26027
rect 27614 26024 27620 26036
rect 27571 25996 27620 26024
rect 27571 25993 27583 25996
rect 27525 25987 27583 25993
rect 27614 25984 27620 25996
rect 27672 25984 27678 26036
rect 28813 26027 28871 26033
rect 28813 25993 28825 26027
rect 28859 26024 28871 26027
rect 31294 26024 31300 26036
rect 28859 25996 29408 26024
rect 28859 25993 28871 25996
rect 28813 25987 28871 25993
rect 25961 25891 26019 25897
rect 25961 25888 25973 25891
rect 25004 25860 25973 25888
rect 25004 25848 25010 25860
rect 25961 25857 25973 25860
rect 26007 25857 26019 25891
rect 25961 25851 26019 25857
rect 26053 25891 26111 25897
rect 26053 25857 26065 25891
rect 26099 25857 26111 25891
rect 26053 25851 26111 25857
rect 23900 25792 24072 25820
rect 23900 25780 23906 25792
rect 24118 25780 24124 25832
rect 24176 25780 24182 25832
rect 24780 25820 24808 25848
rect 26068 25820 26096 25851
rect 26142 25848 26148 25900
rect 26200 25888 26206 25900
rect 26237 25891 26295 25897
rect 26237 25888 26249 25891
rect 26200 25860 26249 25888
rect 26200 25848 26206 25860
rect 26237 25857 26249 25860
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25888 26387 25891
rect 26620 25888 26648 25984
rect 28258 25956 28264 25968
rect 27172 25928 28264 25956
rect 27172 25897 27200 25928
rect 28258 25916 28264 25928
rect 28316 25956 28322 25968
rect 28902 25956 28908 25968
rect 28316 25928 28908 25956
rect 28316 25916 28322 25928
rect 28902 25916 28908 25928
rect 28960 25916 28966 25968
rect 29380 25965 29408 25996
rect 29749 25996 31300 26024
rect 29365 25959 29423 25965
rect 29365 25925 29377 25959
rect 29411 25925 29423 25959
rect 29365 25919 29423 25925
rect 29638 25916 29644 25968
rect 29696 25956 29702 25968
rect 29749 25956 29777 25996
rect 31294 25984 31300 25996
rect 31352 25984 31358 26036
rect 31386 25984 31392 26036
rect 31444 26024 31450 26036
rect 31573 26027 31631 26033
rect 31573 26024 31585 26027
rect 31444 25996 31585 26024
rect 31444 25984 31450 25996
rect 31573 25993 31585 25996
rect 31619 25993 31631 26027
rect 31573 25987 31631 25993
rect 31754 25984 31760 26036
rect 31812 25984 31818 26036
rect 32125 26027 32183 26033
rect 32125 25993 32137 26027
rect 32171 25993 32183 26027
rect 32125 25987 32183 25993
rect 29696 25928 29854 25956
rect 29696 25916 29702 25928
rect 26375 25860 26648 25888
rect 27157 25891 27215 25897
rect 26375 25857 26387 25860
rect 26329 25851 26387 25857
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27430 25848 27436 25900
rect 27488 25888 27494 25900
rect 27893 25891 27951 25897
rect 27893 25888 27905 25891
rect 27488 25860 27905 25888
rect 27488 25848 27494 25860
rect 27893 25857 27905 25860
rect 27939 25857 27951 25891
rect 28350 25888 28356 25900
rect 27893 25851 27951 25857
rect 28000 25860 28356 25888
rect 28000 25829 28028 25860
rect 28350 25848 28356 25860
rect 28408 25848 28414 25900
rect 28994 25848 29000 25900
rect 29052 25848 29058 25900
rect 31481 25891 31539 25897
rect 31481 25857 31493 25891
rect 31527 25857 31539 25891
rect 31481 25851 31539 25857
rect 31941 25891 31999 25897
rect 31941 25857 31953 25891
rect 31987 25888 31999 25891
rect 32140 25888 32168 25987
rect 32398 25984 32404 26036
rect 32456 25984 32462 26036
rect 32582 25984 32588 26036
rect 32640 25984 32646 26036
rect 33962 25984 33968 26036
rect 34020 25984 34026 26036
rect 34992 25996 36400 26024
rect 31987 25860 32168 25888
rect 32416 25888 32444 25984
rect 32490 25916 32496 25968
rect 32548 25916 32554 25968
rect 34992 25956 35020 25996
rect 33888 25928 35020 25956
rect 33888 25897 33916 25928
rect 35342 25916 35348 25968
rect 35400 25916 35406 25968
rect 36372 25965 36400 25996
rect 36357 25959 36415 25965
rect 36357 25925 36369 25959
rect 36403 25925 36415 25959
rect 36357 25919 36415 25925
rect 33873 25891 33931 25897
rect 33873 25888 33885 25891
rect 32416 25860 33885 25888
rect 31987 25857 31999 25860
rect 31941 25851 31999 25857
rect 33873 25857 33885 25860
rect 33919 25857 33931 25891
rect 33873 25851 33931 25857
rect 27985 25823 28043 25829
rect 27985 25820 27997 25823
rect 24780 25792 27997 25820
rect 27985 25789 27997 25792
rect 28031 25789 28043 25823
rect 27985 25783 28043 25789
rect 28169 25823 28227 25829
rect 28169 25789 28181 25823
rect 28215 25820 28227 25823
rect 28810 25820 28816 25832
rect 28215 25792 28816 25820
rect 28215 25789 28227 25792
rect 28169 25783 28227 25789
rect 28810 25780 28816 25792
rect 28868 25780 28874 25832
rect 29086 25780 29092 25832
rect 29144 25780 29150 25832
rect 30374 25780 30380 25832
rect 30432 25820 30438 25832
rect 31113 25823 31171 25829
rect 31113 25820 31125 25823
rect 30432 25792 31125 25820
rect 30432 25780 30438 25792
rect 31113 25789 31125 25792
rect 31159 25789 31171 25823
rect 31113 25783 31171 25789
rect 22738 25752 22744 25764
rect 22664 25724 22744 25752
rect 22738 25712 22744 25724
rect 22796 25712 22802 25764
rect 23290 25712 23296 25764
rect 23348 25712 23354 25764
rect 24762 25712 24768 25764
rect 24820 25752 24826 25764
rect 24820 25724 28948 25752
rect 24820 25712 24826 25724
rect 23385 25687 23443 25693
rect 23385 25684 23397 25687
rect 22297 25656 23397 25684
rect 23385 25653 23397 25656
rect 23431 25653 23443 25687
rect 23385 25647 23443 25653
rect 23474 25644 23480 25696
rect 23532 25644 23538 25696
rect 24026 25644 24032 25696
rect 24084 25644 24090 25696
rect 25682 25644 25688 25696
rect 25740 25684 25746 25696
rect 26510 25684 26516 25696
rect 25740 25656 26516 25684
rect 25740 25644 25746 25656
rect 26510 25644 26516 25656
rect 26568 25644 26574 25696
rect 28920 25684 28948 25724
rect 31496 25684 31524 25851
rect 32766 25780 32772 25832
rect 32824 25780 32830 25832
rect 32950 25780 32956 25832
rect 33008 25820 33014 25832
rect 33778 25820 33784 25832
rect 33008 25792 33784 25820
rect 33008 25780 33014 25792
rect 33778 25780 33784 25792
rect 33836 25820 33842 25832
rect 34057 25823 34115 25829
rect 34057 25820 34069 25823
rect 33836 25792 34069 25820
rect 33836 25780 33842 25792
rect 34057 25789 34069 25792
rect 34103 25789 34115 25823
rect 34057 25783 34115 25789
rect 34330 25780 34336 25832
rect 34388 25780 34394 25832
rect 34606 25780 34612 25832
rect 34664 25780 34670 25832
rect 28920 25656 31524 25684
rect 31754 25644 31760 25696
rect 31812 25684 31818 25696
rect 32490 25684 32496 25696
rect 31812 25656 32496 25684
rect 31812 25644 31818 25656
rect 32490 25644 32496 25656
rect 32548 25644 32554 25696
rect 33502 25644 33508 25696
rect 33560 25644 33566 25696
rect 1104 25594 38272 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38272 25594
rect 1104 25520 38272 25542
rect 5524 25483 5582 25489
rect 5524 25449 5536 25483
rect 5570 25480 5582 25483
rect 5626 25480 5632 25492
rect 5570 25452 5632 25480
rect 5570 25449 5582 25452
rect 5524 25443 5582 25449
rect 5626 25440 5632 25452
rect 5684 25440 5690 25492
rect 5994 25440 6000 25492
rect 6052 25480 6058 25492
rect 7193 25483 7251 25489
rect 7193 25480 7205 25483
rect 6052 25452 7205 25480
rect 6052 25440 6058 25452
rect 7193 25449 7205 25452
rect 7239 25449 7251 25483
rect 7193 25443 7251 25449
rect 7926 25440 7932 25492
rect 7984 25480 7990 25492
rect 9766 25480 9772 25492
rect 7984 25452 9772 25480
rect 7984 25440 7990 25452
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 10410 25440 10416 25492
rect 10468 25480 10474 25492
rect 11609 25483 11667 25489
rect 11609 25480 11621 25483
rect 10468 25452 11621 25480
rect 10468 25440 10474 25452
rect 11609 25449 11621 25452
rect 11655 25449 11667 25483
rect 13262 25480 13268 25492
rect 11609 25443 11667 25449
rect 11992 25452 13268 25480
rect 7009 25415 7067 25421
rect 7009 25381 7021 25415
rect 7055 25412 7067 25415
rect 7650 25412 7656 25424
rect 7055 25384 7656 25412
rect 7055 25381 7067 25384
rect 7009 25375 7067 25381
rect 7650 25372 7656 25384
rect 7708 25372 7714 25424
rect 7742 25304 7748 25356
rect 7800 25304 7806 25356
rect 1670 25236 1676 25288
rect 1728 25236 1734 25288
rect 4985 25279 5043 25285
rect 4985 25245 4997 25279
rect 5031 25245 5043 25279
rect 4985 25239 5043 25245
rect 5077 25279 5135 25285
rect 5077 25245 5089 25279
rect 5123 25276 5135 25279
rect 5261 25279 5319 25285
rect 5261 25276 5273 25279
rect 5123 25248 5273 25276
rect 5123 25245 5135 25248
rect 5077 25239 5135 25245
rect 5261 25245 5273 25248
rect 5307 25245 5319 25279
rect 5261 25239 5319 25245
rect 1946 25168 1952 25220
rect 2004 25168 2010 25220
rect 4062 25208 4068 25220
rect 3174 25180 4068 25208
rect 4062 25168 4068 25180
rect 4120 25168 4126 25220
rect 2774 25100 2780 25152
rect 2832 25140 2838 25152
rect 3421 25143 3479 25149
rect 3421 25140 3433 25143
rect 2832 25112 3433 25140
rect 2832 25100 2838 25112
rect 3421 25109 3433 25112
rect 3467 25109 3479 25143
rect 5000 25140 5028 25239
rect 6638 25236 6644 25288
rect 6696 25236 6702 25288
rect 7561 25279 7619 25285
rect 7561 25245 7573 25279
rect 7607 25276 7619 25279
rect 7944 25276 7972 25440
rect 8018 25372 8024 25424
rect 8076 25372 8082 25424
rect 9674 25412 9680 25424
rect 8588 25384 9680 25412
rect 8036 25285 8064 25372
rect 8588 25285 8616 25384
rect 9674 25372 9680 25384
rect 9732 25372 9738 25424
rect 11425 25415 11483 25421
rect 11425 25381 11437 25415
rect 11471 25412 11483 25415
rect 11992 25412 12020 25452
rect 13262 25440 13268 25452
rect 13320 25440 13326 25492
rect 15378 25440 15384 25492
rect 15436 25480 15442 25492
rect 20162 25480 20168 25492
rect 15436 25452 18552 25480
rect 15436 25440 15442 25452
rect 11471 25384 12020 25412
rect 11471 25381 11483 25384
rect 11425 25375 11483 25381
rect 9953 25347 10011 25353
rect 9953 25313 9965 25347
rect 9999 25344 10011 25347
rect 10042 25344 10048 25356
rect 9999 25316 10048 25344
rect 9999 25313 10011 25316
rect 9953 25307 10011 25313
rect 10042 25304 10048 25316
rect 10100 25304 10106 25356
rect 7607 25248 7972 25276
rect 8021 25279 8079 25285
rect 7607 25245 7619 25248
rect 7561 25239 7619 25245
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 8573 25279 8631 25285
rect 8573 25245 8585 25279
rect 8619 25245 8631 25279
rect 8573 25239 8631 25245
rect 9398 25236 9404 25288
rect 9456 25236 9462 25288
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25276 9551 25279
rect 9677 25279 9735 25285
rect 9677 25276 9689 25279
rect 9539 25248 9689 25276
rect 9539 25245 9551 25248
rect 9493 25239 9551 25245
rect 9677 25245 9689 25248
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 11330 25276 11336 25288
rect 11112 25248 11336 25276
rect 11112 25236 11118 25248
rect 11330 25236 11336 25248
rect 11388 25236 11394 25288
rect 11992 25285 12020 25384
rect 15102 25372 15108 25424
rect 15160 25372 15166 25424
rect 17034 25372 17040 25424
rect 17092 25412 17098 25424
rect 18524 25412 18552 25452
rect 19904 25452 20168 25480
rect 17092 25384 17356 25412
rect 18524 25384 19334 25412
rect 17092 25372 17098 25384
rect 12158 25304 12164 25356
rect 12216 25304 12222 25356
rect 12621 25347 12679 25353
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 12894 25344 12900 25356
rect 12667 25316 12900 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 12894 25304 12900 25316
rect 12952 25344 12958 25356
rect 13354 25344 13360 25356
rect 12952 25316 13360 25344
rect 12952 25304 12958 25316
rect 13354 25304 13360 25316
rect 13412 25304 13418 25356
rect 13722 25304 13728 25356
rect 13780 25304 13786 25356
rect 15120 25330 15148 25372
rect 17328 25353 17356 25384
rect 17313 25347 17371 25353
rect 17313 25313 17325 25347
rect 17359 25313 17371 25347
rect 17313 25307 17371 25313
rect 18598 25304 18604 25356
rect 18656 25304 18662 25356
rect 11977 25279 12035 25285
rect 11977 25245 11989 25279
rect 12023 25245 12035 25279
rect 12805 25279 12863 25285
rect 12805 25276 12817 25279
rect 11977 25239 12035 25245
rect 12728 25248 12817 25276
rect 9416 25208 9444 25236
rect 7576 25180 9444 25208
rect 7576 25140 7604 25180
rect 12728 25152 12756 25248
rect 12805 25245 12817 25248
rect 12851 25245 12863 25279
rect 12805 25239 12863 25245
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25245 13507 25279
rect 13449 25239 13507 25245
rect 13633 25279 13691 25285
rect 13633 25245 13645 25279
rect 13679 25276 13691 25279
rect 14090 25276 14096 25288
rect 13679 25248 14096 25276
rect 13679 25245 13691 25248
rect 13633 25239 13691 25245
rect 12989 25211 13047 25217
rect 12989 25177 13001 25211
rect 13035 25208 13047 25211
rect 13464 25208 13492 25239
rect 14090 25236 14096 25248
rect 14148 25236 14154 25288
rect 14182 25236 14188 25288
rect 14240 25236 14246 25288
rect 14642 25236 14648 25288
rect 14700 25236 14706 25288
rect 15105 25279 15163 25285
rect 15105 25245 15117 25279
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 16577 25279 16635 25285
rect 16577 25245 16589 25279
rect 16623 25245 16635 25279
rect 16577 25239 16635 25245
rect 15120 25208 15148 25239
rect 13035 25180 15148 25208
rect 16592 25208 16620 25239
rect 16666 25236 16672 25288
rect 16724 25276 16730 25288
rect 17221 25279 17279 25285
rect 17221 25276 17233 25279
rect 16724 25248 17233 25276
rect 16724 25236 16730 25248
rect 17221 25245 17233 25248
rect 17267 25245 17279 25279
rect 17221 25239 17279 25245
rect 18138 25236 18144 25288
rect 18196 25236 18202 25288
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25276 18475 25279
rect 18616 25276 18644 25304
rect 18463 25248 18644 25276
rect 18463 25245 18475 25248
rect 18417 25239 18475 25245
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 18785 25279 18843 25285
rect 18785 25276 18797 25279
rect 18748 25248 18797 25276
rect 18748 25236 18754 25248
rect 18785 25245 18797 25248
rect 18831 25245 18843 25279
rect 18785 25239 18843 25245
rect 18877 25279 18935 25285
rect 18877 25245 18889 25279
rect 18923 25276 18935 25279
rect 19306 25276 19334 25384
rect 19702 25276 19708 25288
rect 18923 25248 19196 25276
rect 19306 25248 19708 25276
rect 18923 25245 18935 25248
rect 18877 25239 18935 25245
rect 16758 25208 16764 25220
rect 16592 25180 16764 25208
rect 13035 25177 13047 25180
rect 12989 25171 13047 25177
rect 16758 25168 16764 25180
rect 16816 25208 16822 25220
rect 18156 25208 18184 25236
rect 19168 25220 19196 25248
rect 19702 25236 19708 25248
rect 19760 25276 19766 25288
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19760 25248 19809 25276
rect 19760 25236 19766 25248
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 18509 25211 18567 25217
rect 18509 25208 18521 25211
rect 16816 25180 17264 25208
rect 18156 25180 18521 25208
rect 16816 25168 16822 25180
rect 17236 25152 17264 25180
rect 18509 25177 18521 25180
rect 18555 25177 18567 25211
rect 18509 25171 18567 25177
rect 18601 25211 18659 25217
rect 18601 25177 18613 25211
rect 18647 25177 18659 25211
rect 18601 25171 18659 25177
rect 5000 25112 7604 25140
rect 3421 25103 3479 25109
rect 7650 25100 7656 25152
rect 7708 25100 7714 25152
rect 7834 25100 7840 25152
rect 7892 25140 7898 25152
rect 8113 25143 8171 25149
rect 8113 25140 8125 25143
rect 7892 25112 8125 25140
rect 7892 25100 7898 25112
rect 8113 25109 8125 25112
rect 8159 25109 8171 25143
rect 8113 25103 8171 25109
rect 8386 25100 8392 25152
rect 8444 25100 8450 25152
rect 12066 25100 12072 25152
rect 12124 25100 12130 25152
rect 12710 25100 12716 25152
rect 12768 25100 12774 25152
rect 13078 25100 13084 25152
rect 13136 25140 13142 25152
rect 14854 25143 14912 25149
rect 14854 25140 14866 25143
rect 13136 25112 14866 25140
rect 13136 25100 13142 25112
rect 14854 25109 14866 25112
rect 14900 25109 14912 25143
rect 14854 25103 14912 25109
rect 17218 25100 17224 25152
rect 17276 25100 17282 25152
rect 18230 25100 18236 25152
rect 18288 25100 18294 25152
rect 18616 25140 18644 25171
rect 19150 25168 19156 25220
rect 19208 25168 19214 25220
rect 19904 25140 19932 25452
rect 20162 25440 20168 25452
rect 20220 25440 20226 25492
rect 20346 25440 20352 25492
rect 20404 25440 20410 25492
rect 20714 25440 20720 25492
rect 20772 25480 20778 25492
rect 21726 25480 21732 25492
rect 20772 25452 21732 25480
rect 20772 25440 20778 25452
rect 21726 25440 21732 25452
rect 21784 25440 21790 25492
rect 22649 25483 22707 25489
rect 22649 25449 22661 25483
rect 22695 25449 22707 25483
rect 22649 25443 22707 25449
rect 22278 25412 22284 25424
rect 19996 25384 22284 25412
rect 19996 25285 20024 25384
rect 22278 25372 22284 25384
rect 22336 25372 22342 25424
rect 22554 25372 22560 25424
rect 22612 25412 22618 25424
rect 22664 25412 22692 25443
rect 22738 25440 22744 25492
rect 22796 25480 22802 25492
rect 23017 25483 23075 25489
rect 23017 25480 23029 25483
rect 22796 25452 23029 25480
rect 22796 25440 22802 25452
rect 23017 25449 23029 25452
rect 23063 25449 23075 25483
rect 23017 25443 23075 25449
rect 24026 25440 24032 25492
rect 24084 25440 24090 25492
rect 24397 25483 24455 25489
rect 24397 25449 24409 25483
rect 24443 25480 24455 25483
rect 24670 25480 24676 25492
rect 24443 25452 24676 25480
rect 24443 25449 24455 25452
rect 24397 25443 24455 25449
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 25314 25440 25320 25492
rect 25372 25480 25378 25492
rect 26142 25480 26148 25492
rect 25372 25452 26148 25480
rect 25372 25440 25378 25452
rect 26142 25440 26148 25452
rect 26200 25440 26206 25492
rect 26878 25440 26884 25492
rect 26936 25440 26942 25492
rect 28353 25483 28411 25489
rect 28353 25449 28365 25483
rect 28399 25480 28411 25483
rect 28994 25480 29000 25492
rect 28399 25452 29000 25480
rect 28399 25449 28411 25452
rect 28353 25443 28411 25449
rect 28994 25440 29000 25452
rect 29052 25440 29058 25492
rect 33502 25440 33508 25492
rect 33560 25440 33566 25492
rect 34057 25483 34115 25489
rect 34057 25449 34069 25483
rect 34103 25480 34115 25483
rect 34606 25480 34612 25492
rect 34103 25452 34612 25480
rect 34103 25449 34115 25452
rect 34057 25443 34115 25449
rect 34606 25440 34612 25452
rect 34664 25440 34670 25492
rect 24044 25412 24072 25440
rect 26896 25412 26924 25440
rect 32950 25412 32956 25424
rect 22612 25384 24072 25412
rect 24504 25384 26372 25412
rect 26896 25384 32956 25412
rect 22612 25372 22618 25384
rect 20438 25304 20444 25356
rect 20496 25304 20502 25356
rect 22741 25347 22799 25353
rect 22741 25344 22753 25347
rect 21008 25316 22232 25344
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25245 20039 25279
rect 19981 25239 20039 25245
rect 20165 25279 20223 25285
rect 20165 25245 20177 25279
rect 20211 25245 20223 25279
rect 20165 25239 20223 25245
rect 20073 25211 20131 25217
rect 20073 25177 20085 25211
rect 20119 25177 20131 25211
rect 20073 25171 20131 25177
rect 18616 25112 19932 25140
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 20088 25140 20116 25171
rect 20036 25112 20116 25140
rect 20180 25140 20208 25239
rect 20456 25208 20484 25304
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25276 20683 25279
rect 20714 25276 20720 25288
rect 20671 25248 20720 25276
rect 20671 25245 20683 25248
rect 20625 25239 20683 25245
rect 20714 25236 20720 25248
rect 20772 25236 20778 25288
rect 21008 25285 21036 25316
rect 22204 25288 22232 25316
rect 22388 25316 22753 25344
rect 22388 25288 22416 25316
rect 22741 25313 22753 25316
rect 22787 25313 22799 25347
rect 22741 25307 22799 25313
rect 22922 25304 22928 25356
rect 22980 25344 22986 25356
rect 23106 25344 23112 25356
rect 22980 25316 23112 25344
rect 22980 25304 22986 25316
rect 23106 25304 23112 25316
rect 23164 25304 23170 25356
rect 23842 25344 23848 25356
rect 23216 25316 23848 25344
rect 20993 25279 21051 25285
rect 20993 25245 21005 25279
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 21284 25208 21312 25239
rect 22186 25236 22192 25288
rect 22244 25236 22250 25288
rect 22370 25236 22376 25288
rect 22428 25236 22434 25288
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25276 22707 25279
rect 23216 25276 23244 25316
rect 23842 25304 23848 25316
rect 23900 25304 23906 25356
rect 22695 25248 23244 25276
rect 22695 25245 22707 25248
rect 22649 25239 22707 25245
rect 23290 25236 23296 25288
rect 23348 25276 23354 25288
rect 24504 25276 24532 25384
rect 24578 25304 24584 25356
rect 24636 25304 24642 25356
rect 24670 25304 24676 25356
rect 24728 25344 24734 25356
rect 24857 25347 24915 25353
rect 24857 25344 24869 25347
rect 24728 25316 24869 25344
rect 24728 25304 24734 25316
rect 24857 25313 24869 25316
rect 24903 25313 24915 25347
rect 24857 25307 24915 25313
rect 24949 25347 25007 25353
rect 24949 25313 24961 25347
rect 24995 25313 25007 25347
rect 26344 25344 26372 25384
rect 26878 25344 26884 25356
rect 24949 25307 25007 25313
rect 25332 25316 26280 25344
rect 23348 25248 24532 25276
rect 24596 25276 24624 25304
rect 24964 25276 24992 25307
rect 24596 25248 24992 25276
rect 23348 25236 23354 25248
rect 20456 25180 21312 25208
rect 21542 25168 21548 25220
rect 21600 25168 21606 25220
rect 24946 25208 24952 25220
rect 22848 25180 24952 25208
rect 20622 25140 20628 25152
rect 20180 25112 20628 25140
rect 20036 25100 20042 25112
rect 20622 25100 20628 25112
rect 20680 25140 20686 25152
rect 22848 25140 22876 25180
rect 24946 25168 24952 25180
rect 25004 25208 25010 25220
rect 25332 25208 25360 25316
rect 25593 25279 25651 25285
rect 25593 25276 25605 25279
rect 25424 25248 25605 25276
rect 25424 25220 25452 25248
rect 25593 25245 25605 25248
rect 25639 25245 25651 25279
rect 25593 25239 25651 25245
rect 25682 25236 25688 25288
rect 25740 25236 25746 25288
rect 26252 25285 26280 25316
rect 26344 25316 26884 25344
rect 26344 25285 26372 25316
rect 26878 25304 26884 25316
rect 26936 25304 26942 25356
rect 29012 25353 29040 25384
rect 32950 25372 32956 25384
rect 33008 25372 33014 25424
rect 28997 25347 29055 25353
rect 28997 25313 29009 25347
rect 29043 25313 29055 25347
rect 28997 25307 29055 25313
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 25961 25279 26019 25285
rect 25961 25245 25973 25279
rect 26007 25276 26019 25279
rect 26237 25279 26295 25285
rect 26007 25248 26188 25276
rect 26007 25245 26019 25248
rect 25961 25239 26019 25245
rect 25004 25180 25360 25208
rect 25004 25168 25010 25180
rect 25406 25168 25412 25220
rect 25464 25208 25470 25220
rect 25792 25208 25820 25239
rect 26053 25211 26111 25217
rect 26053 25208 26065 25211
rect 25464 25180 25728 25208
rect 25792 25180 26065 25208
rect 25464 25168 25470 25180
rect 20680 25112 22876 25140
rect 20680 25100 20686 25112
rect 22922 25100 22928 25152
rect 22980 25140 22986 25152
rect 24765 25143 24823 25149
rect 24765 25140 24777 25143
rect 22980 25112 24777 25140
rect 22980 25100 22986 25112
rect 24765 25109 24777 25112
rect 24811 25140 24823 25143
rect 25498 25140 25504 25152
rect 24811 25112 25504 25140
rect 24811 25109 24823 25112
rect 24765 25103 24823 25109
rect 25498 25100 25504 25112
rect 25556 25100 25562 25152
rect 25700 25140 25728 25180
rect 26053 25177 26065 25180
rect 26099 25177 26111 25211
rect 26160 25208 26188 25248
rect 26237 25245 26249 25279
rect 26283 25245 26295 25279
rect 26237 25239 26295 25245
rect 26329 25279 26387 25285
rect 26329 25245 26341 25279
rect 26375 25245 26387 25279
rect 26329 25239 26387 25245
rect 26510 25236 26516 25288
rect 26568 25236 26574 25288
rect 26602 25236 26608 25288
rect 26660 25236 26666 25288
rect 26694 25236 26700 25288
rect 26752 25236 26758 25288
rect 28721 25279 28779 25285
rect 28721 25276 28733 25279
rect 26804 25248 28733 25276
rect 26712 25208 26740 25236
rect 26160 25180 26740 25208
rect 26053 25171 26111 25177
rect 26804 25140 26832 25248
rect 28721 25245 28733 25248
rect 28767 25276 28779 25279
rect 30190 25276 30196 25288
rect 28767 25248 30196 25276
rect 28767 25245 28779 25248
rect 28721 25239 28779 25245
rect 30190 25236 30196 25248
rect 30248 25276 30254 25288
rect 30374 25276 30380 25288
rect 30248 25248 30380 25276
rect 30248 25236 30254 25248
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 32030 25236 32036 25288
rect 32088 25276 32094 25288
rect 32490 25276 32496 25288
rect 32088 25248 32496 25276
rect 32088 25236 32094 25248
rect 32490 25236 32496 25248
rect 32548 25236 32554 25288
rect 33520 25276 33548 25440
rect 34241 25279 34299 25285
rect 34241 25276 34253 25279
rect 33520 25248 34253 25276
rect 34241 25245 34253 25248
rect 34287 25245 34299 25279
rect 34241 25239 34299 25245
rect 28813 25211 28871 25217
rect 28813 25208 28825 25211
rect 28552 25180 28825 25208
rect 28552 25152 28580 25180
rect 28813 25177 28825 25180
rect 28859 25177 28871 25211
rect 28813 25171 28871 25177
rect 25700 25112 26832 25140
rect 28534 25100 28540 25152
rect 28592 25100 28598 25152
rect 1104 25050 38272 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38272 25050
rect 1104 24976 38272 24998
rect 1578 24896 1584 24948
rect 1636 24896 1642 24948
rect 1946 24896 1952 24948
rect 2004 24936 2010 24948
rect 2133 24939 2191 24945
rect 2133 24936 2145 24939
rect 2004 24908 2145 24936
rect 2004 24896 2010 24908
rect 2133 24905 2145 24908
rect 2179 24905 2191 24939
rect 2133 24899 2191 24905
rect 7650 24896 7656 24948
rect 7708 24936 7714 24948
rect 7708 24908 9444 24936
rect 7708 24896 7714 24908
rect 1670 24828 1676 24880
rect 1728 24868 1734 24880
rect 1728 24840 2728 24868
rect 1728 24828 1734 24840
rect 1486 24760 1492 24812
rect 1544 24760 1550 24812
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24800 2375 24803
rect 2700 24800 2728 24840
rect 2774 24828 2780 24880
rect 2832 24828 2838 24880
rect 6638 24828 6644 24880
rect 6696 24828 6702 24880
rect 8113 24871 8171 24877
rect 8113 24837 8125 24871
rect 8159 24868 8171 24871
rect 8386 24868 8392 24880
rect 8159 24840 8392 24868
rect 8159 24837 8171 24840
rect 8113 24831 8171 24837
rect 8386 24828 8392 24840
rect 8444 24828 8450 24880
rect 8662 24828 8668 24880
rect 8720 24828 8726 24880
rect 9416 24868 9444 24908
rect 9674 24896 9680 24948
rect 9732 24936 9738 24948
rect 9769 24939 9827 24945
rect 9769 24936 9781 24939
rect 9732 24908 9781 24936
rect 9732 24896 9738 24908
rect 9769 24905 9781 24908
rect 9815 24905 9827 24939
rect 9769 24899 9827 24905
rect 10042 24896 10048 24948
rect 10100 24936 10106 24948
rect 10137 24939 10195 24945
rect 10137 24936 10149 24939
rect 10100 24908 10149 24936
rect 10100 24896 10106 24908
rect 10137 24905 10149 24908
rect 10183 24936 10195 24939
rect 12250 24936 12256 24948
rect 10183 24908 12256 24936
rect 10183 24905 10195 24908
rect 10137 24899 10195 24905
rect 12250 24896 12256 24908
rect 12308 24896 12314 24948
rect 15930 24936 15936 24948
rect 12406 24908 15936 24936
rect 12406 24868 12434 24908
rect 15930 24896 15936 24908
rect 15988 24896 15994 24948
rect 18414 24896 18420 24948
rect 18472 24896 18478 24948
rect 20806 24896 20812 24948
rect 20864 24936 20870 24948
rect 20993 24939 21051 24945
rect 20993 24936 21005 24939
rect 20864 24908 21005 24936
rect 20864 24896 20870 24908
rect 20993 24905 21005 24908
rect 21039 24905 21051 24939
rect 20993 24899 21051 24905
rect 22462 24896 22468 24948
rect 22520 24936 22526 24948
rect 22741 24939 22799 24945
rect 22741 24936 22753 24939
rect 22520 24908 22753 24936
rect 22520 24896 22526 24908
rect 22741 24905 22753 24908
rect 22787 24905 22799 24939
rect 25774 24936 25780 24948
rect 22741 24899 22799 24905
rect 25700 24908 25780 24936
rect 18432 24868 18460 24896
rect 9416 24840 12434 24868
rect 13740 24840 13952 24868
rect 6178 24800 6184 24812
rect 2363 24772 2452 24800
rect 2700 24772 2774 24800
rect 4830 24786 6184 24800
rect 2363 24769 2375 24772
rect 2317 24763 2375 24769
rect 2424 24673 2452 24772
rect 2409 24667 2467 24673
rect 2409 24633 2421 24667
rect 2455 24633 2467 24667
rect 2746 24664 2774 24772
rect 4816 24772 6184 24786
rect 2866 24692 2872 24744
rect 2924 24692 2930 24744
rect 3053 24735 3111 24741
rect 3053 24701 3065 24735
rect 3099 24732 3111 24735
rect 3142 24732 3148 24744
rect 3099 24704 3148 24732
rect 3099 24701 3111 24704
rect 3053 24695 3111 24701
rect 3142 24692 3148 24704
rect 3200 24692 3206 24744
rect 3421 24735 3479 24741
rect 3421 24701 3433 24735
rect 3467 24732 3479 24735
rect 3467 24704 3556 24732
rect 3467 24701 3479 24704
rect 3421 24695 3479 24701
rect 3528 24664 3556 24704
rect 3694 24692 3700 24744
rect 3752 24692 3758 24744
rect 4062 24692 4068 24744
rect 4120 24732 4126 24744
rect 4816 24732 4844 24772
rect 6178 24760 6184 24772
rect 6236 24800 6242 24812
rect 6656 24800 6684 24828
rect 6236 24772 6684 24800
rect 6236 24760 6242 24772
rect 11698 24760 11704 24812
rect 11756 24760 11762 24812
rect 12161 24803 12219 24809
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12526 24800 12532 24812
rect 12207 24772 12532 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 12621 24803 12679 24809
rect 12621 24769 12633 24803
rect 12667 24800 12679 24803
rect 13357 24803 13415 24809
rect 12667 24772 13308 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 4120 24704 4844 24732
rect 4120 24692 4126 24704
rect 5442 24692 5448 24744
rect 5500 24692 5506 24744
rect 7834 24692 7840 24744
rect 7892 24692 7898 24744
rect 9766 24692 9772 24744
rect 9824 24732 9830 24744
rect 10226 24732 10232 24744
rect 9824 24704 10232 24732
rect 9824 24692 9830 24704
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 10413 24735 10471 24741
rect 10413 24701 10425 24735
rect 10459 24701 10471 24735
rect 10413 24695 10471 24701
rect 5460 24664 5488 24692
rect 2746 24636 3556 24664
rect 2409 24627 2467 24633
rect 3528 24596 3556 24636
rect 4724 24636 5488 24664
rect 4724 24596 4752 24636
rect 3528 24568 4752 24596
rect 4798 24556 4804 24608
rect 4856 24596 4862 24608
rect 5169 24599 5227 24605
rect 5169 24596 5181 24599
rect 4856 24568 5181 24596
rect 4856 24556 4862 24568
rect 5169 24565 5181 24568
rect 5215 24596 5227 24599
rect 5258 24596 5264 24608
rect 5215 24568 5264 24596
rect 5215 24565 5227 24568
rect 5169 24559 5227 24565
rect 5258 24556 5264 24568
rect 5316 24556 5322 24608
rect 9585 24599 9643 24605
rect 9585 24565 9597 24599
rect 9631 24596 9643 24599
rect 10042 24596 10048 24608
rect 9631 24568 10048 24596
rect 9631 24565 9643 24568
rect 9585 24559 9643 24565
rect 10042 24556 10048 24568
rect 10100 24556 10106 24608
rect 10428 24596 10456 24695
rect 11716 24664 11744 24760
rect 13280 24741 13308 24772
rect 13357 24769 13369 24803
rect 13403 24769 13415 24803
rect 13357 24763 13415 24769
rect 12713 24735 12771 24741
rect 12713 24701 12725 24735
rect 12759 24701 12771 24735
rect 12713 24695 12771 24701
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24701 13323 24735
rect 13372 24732 13400 24763
rect 13538 24760 13544 24812
rect 13596 24800 13602 24812
rect 13740 24809 13768 24840
rect 13725 24803 13783 24809
rect 13725 24800 13737 24803
rect 13596 24772 13737 24800
rect 13596 24760 13602 24772
rect 13725 24769 13737 24772
rect 13771 24769 13783 24803
rect 13725 24763 13783 24769
rect 13814 24760 13820 24812
rect 13872 24760 13878 24812
rect 13924 24800 13952 24840
rect 17880 24840 18460 24868
rect 14369 24803 14427 24809
rect 14369 24800 14381 24803
rect 13924 24772 14381 24800
rect 14369 24769 14381 24772
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 14734 24760 14740 24812
rect 14792 24800 14798 24812
rect 14829 24803 14887 24809
rect 14829 24800 14841 24803
rect 14792 24772 14841 24800
rect 14792 24760 14798 24772
rect 14829 24769 14841 24772
rect 14875 24769 14887 24803
rect 14829 24763 14887 24769
rect 16114 24760 16120 24812
rect 16172 24760 16178 24812
rect 16298 24760 16304 24812
rect 16356 24760 16362 24812
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 17880 24809 17908 24840
rect 19426 24828 19432 24880
rect 19484 24868 19490 24880
rect 20622 24868 20628 24880
rect 19484 24840 20628 24868
rect 19484 24828 19490 24840
rect 20622 24828 20628 24840
rect 20680 24828 20686 24880
rect 20717 24871 20775 24877
rect 20717 24837 20729 24871
rect 20763 24868 20775 24871
rect 20763 24840 22233 24868
rect 20763 24837 20775 24840
rect 20717 24831 20775 24837
rect 21284 24812 21312 24840
rect 17037 24803 17095 24809
rect 17037 24800 17049 24803
rect 16724 24772 17049 24800
rect 16724 24760 16730 24772
rect 17037 24769 17049 24772
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24769 17923 24803
rect 17865 24763 17923 24769
rect 17954 24760 17960 24812
rect 18012 24760 18018 24812
rect 18046 24760 18052 24812
rect 18104 24760 18110 24812
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 18233 24803 18291 24809
rect 18233 24800 18245 24803
rect 18196 24772 18245 24800
rect 18196 24760 18202 24772
rect 18233 24769 18245 24772
rect 18279 24769 18291 24803
rect 18233 24763 18291 24769
rect 18414 24760 18420 24812
rect 18472 24800 18478 24812
rect 18601 24803 18659 24809
rect 18601 24800 18613 24803
rect 18472 24772 18613 24800
rect 18472 24760 18478 24772
rect 18601 24769 18613 24772
rect 18647 24769 18659 24803
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 18601 24763 18659 24769
rect 18800 24772 19165 24800
rect 13832 24732 13860 24760
rect 13372 24704 13860 24732
rect 13909 24735 13967 24741
rect 13265 24695 13323 24701
rect 13909 24701 13921 24735
rect 13955 24701 13967 24735
rect 13909 24695 13967 24701
rect 11977 24667 12035 24673
rect 11977 24664 11989 24667
rect 11716 24636 11989 24664
rect 11977 24633 11989 24636
rect 12023 24633 12035 24667
rect 11977 24627 12035 24633
rect 12342 24596 12348 24608
rect 10428 24568 12348 24596
rect 12342 24556 12348 24568
rect 12400 24596 12406 24608
rect 12728 24596 12756 24695
rect 13280 24608 13308 24695
rect 13354 24624 13360 24676
rect 13412 24664 13418 24676
rect 13924 24664 13952 24695
rect 14090 24692 14096 24744
rect 14148 24692 14154 24744
rect 14182 24692 14188 24744
rect 14240 24692 14246 24744
rect 15105 24735 15163 24741
rect 15105 24701 15117 24735
rect 15151 24732 15163 24735
rect 17126 24732 17132 24744
rect 15151 24704 17132 24732
rect 15151 24701 15163 24704
rect 15105 24695 15163 24701
rect 17126 24692 17132 24704
rect 17184 24692 17190 24744
rect 17313 24735 17371 24741
rect 17313 24701 17325 24735
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 17589 24735 17647 24741
rect 17589 24701 17601 24735
rect 17635 24732 17647 24735
rect 18690 24732 18696 24744
rect 17635 24704 18696 24732
rect 17635 24701 17647 24704
rect 17589 24695 17647 24701
rect 13412 24636 13952 24664
rect 13412 24624 13418 24636
rect 12400 24568 12756 24596
rect 12400 24556 12406 24568
rect 13262 24556 13268 24608
rect 13320 24556 13326 24608
rect 13630 24556 13636 24608
rect 13688 24596 13694 24608
rect 14108 24596 14136 24692
rect 16022 24624 16028 24676
rect 16080 24664 16086 24676
rect 17328 24664 17356 24695
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 18322 24664 18328 24676
rect 16080 24636 17264 24664
rect 17328 24636 18328 24664
rect 16080 24624 16086 24636
rect 13688 24568 14136 24596
rect 13688 24556 13694 24568
rect 16482 24556 16488 24608
rect 16540 24556 16546 24608
rect 17236 24596 17264 24636
rect 18322 24624 18328 24636
rect 18380 24624 18386 24676
rect 18800 24596 18828 24772
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 20530 24809 20536 24812
rect 20349 24803 20407 24809
rect 20349 24800 20361 24803
rect 20220 24772 20361 24800
rect 20220 24760 20226 24772
rect 20349 24769 20361 24772
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20497 24803 20536 24809
rect 20497 24769 20509 24803
rect 20497 24763 20536 24769
rect 20530 24760 20536 24763
rect 20588 24760 20594 24812
rect 20898 24809 20904 24812
rect 20855 24803 20904 24809
rect 20855 24769 20867 24803
rect 20901 24769 20904 24803
rect 20855 24763 20904 24769
rect 20898 24760 20904 24763
rect 20956 24760 20962 24812
rect 21266 24760 21272 24812
rect 21324 24760 21330 24812
rect 22094 24760 22100 24812
rect 22152 24760 22158 24812
rect 22205 24809 22233 24840
rect 24578 24828 24584 24880
rect 24636 24868 24642 24880
rect 25700 24877 25728 24908
rect 25774 24896 25780 24908
rect 25832 24896 25838 24948
rect 27982 24896 27988 24948
rect 28040 24936 28046 24948
rect 28261 24939 28319 24945
rect 28261 24936 28273 24939
rect 28040 24908 28273 24936
rect 28040 24896 28046 24908
rect 28261 24905 28273 24908
rect 28307 24905 28319 24939
rect 28261 24899 28319 24905
rect 28350 24896 28356 24948
rect 28408 24936 28414 24948
rect 28445 24939 28503 24945
rect 28445 24936 28457 24939
rect 28408 24908 28457 24936
rect 28408 24896 28414 24908
rect 28445 24905 28457 24908
rect 28491 24905 28503 24939
rect 28445 24899 28503 24905
rect 30650 24896 30656 24948
rect 30708 24936 30714 24948
rect 33870 24936 33876 24948
rect 30708 24908 33876 24936
rect 30708 24896 30714 24908
rect 33870 24896 33876 24908
rect 33928 24896 33934 24948
rect 25685 24871 25743 24877
rect 25685 24868 25697 24871
rect 24636 24840 25697 24868
rect 24636 24828 24642 24840
rect 25685 24837 25697 24840
rect 25731 24837 25743 24871
rect 25685 24831 25743 24837
rect 26694 24828 26700 24880
rect 26752 24828 26758 24880
rect 27430 24828 27436 24880
rect 27488 24868 27494 24880
rect 31754 24868 31760 24880
rect 27488 24840 31760 24868
rect 27488 24828 27494 24840
rect 31754 24828 31760 24840
rect 31812 24828 31818 24880
rect 32490 24828 32496 24880
rect 32548 24868 32554 24880
rect 32548 24840 32628 24868
rect 32548 24828 32554 24840
rect 22190 24803 22248 24809
rect 22190 24769 22202 24803
rect 22236 24769 22248 24803
rect 22190 24763 22248 24769
rect 22278 24760 22284 24812
rect 22336 24800 22342 24812
rect 22373 24803 22431 24809
rect 22373 24800 22385 24803
rect 22336 24772 22385 24800
rect 22336 24760 22342 24772
rect 22373 24769 22385 24772
rect 22419 24769 22431 24803
rect 22373 24763 22431 24769
rect 22462 24760 22468 24812
rect 22520 24760 22526 24812
rect 22562 24803 22620 24809
rect 22562 24769 22574 24803
rect 22608 24800 22620 24803
rect 24210 24800 24216 24812
rect 22608 24772 24216 24800
rect 22608 24769 22620 24772
rect 22562 24763 22620 24769
rect 18877 24735 18935 24741
rect 18877 24701 18889 24735
rect 18923 24701 18935 24735
rect 18877 24695 18935 24701
rect 19429 24735 19487 24741
rect 19429 24701 19441 24735
rect 19475 24732 19487 24735
rect 20990 24732 20996 24744
rect 19475 24704 20996 24732
rect 19475 24701 19487 24704
rect 19429 24695 19487 24701
rect 17236 24568 18828 24596
rect 18892 24596 18920 24695
rect 20990 24692 20996 24704
rect 21048 24692 21054 24744
rect 19058 24624 19064 24676
rect 19116 24664 19122 24676
rect 22572 24664 22600 24763
rect 24210 24760 24216 24772
rect 24268 24760 24274 24812
rect 24946 24760 24952 24812
rect 25004 24760 25010 24812
rect 25498 24760 25504 24812
rect 25556 24760 25562 24812
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24769 25835 24803
rect 25777 24763 25835 24769
rect 25869 24803 25927 24809
rect 25869 24769 25881 24803
rect 25915 24800 25927 24803
rect 26050 24800 26056 24812
rect 25915 24772 26056 24800
rect 25915 24769 25927 24772
rect 25869 24763 25927 24769
rect 24964 24732 24992 24760
rect 25792 24732 25820 24763
rect 26050 24760 26056 24772
rect 26108 24760 26114 24812
rect 26712 24800 26740 24828
rect 27522 24800 27528 24812
rect 26712 24772 27528 24800
rect 27522 24760 27528 24772
rect 27580 24760 27586 24812
rect 28169 24803 28227 24809
rect 28169 24769 28181 24803
rect 28215 24800 28227 24803
rect 28258 24800 28264 24812
rect 28215 24772 28264 24800
rect 28215 24769 28227 24772
rect 28169 24763 28227 24769
rect 28258 24760 28264 24772
rect 28316 24760 28322 24812
rect 28626 24760 28632 24812
rect 28684 24760 28690 24812
rect 29365 24803 29423 24809
rect 29365 24800 29377 24803
rect 28736 24772 29377 24800
rect 26510 24732 26516 24744
rect 24964 24704 25820 24732
rect 26068 24704 26516 24732
rect 26068 24673 26096 24704
rect 26510 24692 26516 24704
rect 26568 24692 26574 24744
rect 26694 24692 26700 24744
rect 26752 24732 26758 24744
rect 28736 24732 28764 24772
rect 29365 24769 29377 24772
rect 29411 24769 29423 24803
rect 29365 24763 29423 24769
rect 29549 24803 29607 24809
rect 29549 24769 29561 24803
rect 29595 24769 29607 24803
rect 29549 24763 29607 24769
rect 29641 24803 29699 24809
rect 29641 24769 29653 24803
rect 29687 24800 29699 24803
rect 29914 24800 29920 24812
rect 29687 24772 29920 24800
rect 29687 24769 29699 24772
rect 29641 24763 29699 24769
rect 26752 24704 28764 24732
rect 26752 24692 26758 24704
rect 28902 24692 28908 24744
rect 28960 24732 28966 24744
rect 29564 24732 29592 24763
rect 29914 24760 29920 24772
rect 29972 24760 29978 24812
rect 32122 24760 32128 24812
rect 32180 24760 32186 24812
rect 32306 24760 32312 24812
rect 32364 24760 32370 24812
rect 32398 24760 32404 24812
rect 32456 24760 32462 24812
rect 32600 24809 32628 24840
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24769 32643 24803
rect 32585 24763 32643 24769
rect 32677 24803 32735 24809
rect 32677 24769 32689 24803
rect 32723 24769 32735 24803
rect 32677 24763 32735 24769
rect 28960 24704 29592 24732
rect 28960 24692 28966 24704
rect 19116 24636 22600 24664
rect 26053 24667 26111 24673
rect 19116 24624 19122 24636
rect 26053 24633 26065 24667
rect 26099 24633 26111 24667
rect 26053 24627 26111 24633
rect 26602 24624 26608 24676
rect 26660 24664 26666 24676
rect 30466 24664 30472 24676
rect 26660 24636 30472 24664
rect 26660 24624 26666 24636
rect 30466 24624 30472 24636
rect 30524 24624 30530 24676
rect 32030 24624 32036 24676
rect 32088 24664 32094 24676
rect 32401 24667 32459 24673
rect 32088 24636 32352 24664
rect 32088 24624 32094 24636
rect 21082 24596 21088 24608
rect 18892 24568 21088 24596
rect 21082 24556 21088 24568
rect 21140 24596 21146 24608
rect 22186 24596 22192 24608
rect 21140 24568 22192 24596
rect 21140 24556 21146 24568
rect 22186 24556 22192 24568
rect 22244 24556 22250 24608
rect 29181 24599 29239 24605
rect 29181 24565 29193 24599
rect 29227 24596 29239 24599
rect 30650 24596 30656 24608
rect 29227 24568 30656 24596
rect 29227 24565 29239 24568
rect 29181 24559 29239 24565
rect 30650 24556 30656 24568
rect 30708 24556 30714 24608
rect 32214 24556 32220 24608
rect 32272 24556 32278 24608
rect 32324 24596 32352 24636
rect 32401 24633 32413 24667
rect 32447 24664 32459 24667
rect 32582 24664 32588 24676
rect 32447 24636 32588 24664
rect 32447 24633 32459 24636
rect 32401 24627 32459 24633
rect 32582 24624 32588 24636
rect 32640 24664 32646 24676
rect 32692 24664 32720 24763
rect 32858 24760 32864 24812
rect 32916 24760 32922 24812
rect 32950 24760 32956 24812
rect 33008 24800 33014 24812
rect 34793 24803 34851 24809
rect 34793 24800 34805 24803
rect 33008 24772 34805 24800
rect 33008 24760 33014 24772
rect 34793 24769 34805 24772
rect 34839 24769 34851 24803
rect 34793 24763 34851 24769
rect 32640 24636 32720 24664
rect 32640 24624 32646 24636
rect 32677 24599 32735 24605
rect 32677 24596 32689 24599
rect 32324 24568 32689 24596
rect 32677 24565 32689 24568
rect 32723 24565 32735 24599
rect 32677 24559 32735 24565
rect 34885 24599 34943 24605
rect 34885 24565 34897 24599
rect 34931 24596 34943 24599
rect 35342 24596 35348 24608
rect 34931 24568 35348 24596
rect 34931 24565 34943 24568
rect 34885 24559 34943 24565
rect 35342 24556 35348 24568
rect 35400 24556 35406 24608
rect 1104 24506 38272 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38272 24506
rect 1104 24432 38272 24454
rect 3694 24352 3700 24404
rect 3752 24392 3758 24404
rect 3973 24395 4031 24401
rect 3973 24392 3985 24395
rect 3752 24364 3985 24392
rect 3752 24352 3758 24364
rect 3973 24361 3985 24364
rect 4019 24361 4031 24395
rect 3973 24355 4031 24361
rect 8662 24352 8668 24404
rect 8720 24352 8726 24404
rect 11241 24395 11299 24401
rect 11241 24361 11253 24395
rect 11287 24392 11299 24395
rect 12066 24392 12072 24404
rect 11287 24364 12072 24392
rect 11287 24361 11299 24364
rect 11241 24355 11299 24361
rect 12066 24352 12072 24364
rect 12124 24352 12130 24404
rect 12526 24352 12532 24404
rect 12584 24392 12590 24404
rect 12584 24364 14596 24392
rect 12584 24352 12590 24364
rect 4433 24327 4491 24333
rect 4433 24293 4445 24327
rect 4479 24293 4491 24327
rect 4433 24287 4491 24293
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4448 24188 4476 24287
rect 4985 24259 5043 24265
rect 4985 24256 4997 24259
rect 4203 24160 4476 24188
rect 4724 24228 4997 24256
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 3142 24080 3148 24132
rect 3200 24120 3206 24132
rect 4724 24120 4752 24228
rect 4985 24225 4997 24228
rect 5031 24225 5043 24259
rect 4985 24219 5043 24225
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 5000 24188 5028 24219
rect 5442 24216 5448 24268
rect 5500 24256 5506 24268
rect 6457 24259 6515 24265
rect 6457 24256 6469 24259
rect 5500 24228 6469 24256
rect 5500 24216 5506 24228
rect 6457 24225 6469 24228
rect 6503 24256 6515 24259
rect 8294 24256 8300 24268
rect 6503 24228 8300 24256
rect 6503 24225 6515 24228
rect 6457 24219 6515 24225
rect 8294 24216 8300 24228
rect 8352 24216 8358 24268
rect 8680 24188 8708 24352
rect 12621 24327 12679 24333
rect 12621 24293 12633 24327
rect 12667 24324 12679 24327
rect 12710 24324 12716 24336
rect 12667 24296 12716 24324
rect 12667 24293 12679 24296
rect 12621 24287 12679 24293
rect 12710 24284 12716 24296
rect 12768 24284 12774 24336
rect 13630 24284 13636 24336
rect 13688 24284 13694 24336
rect 14568 24333 14596 24364
rect 14642 24352 14648 24404
rect 14700 24392 14706 24404
rect 14829 24395 14887 24401
rect 14829 24392 14841 24395
rect 14700 24364 14841 24392
rect 14700 24352 14706 24364
rect 14829 24361 14841 24364
rect 14875 24361 14887 24395
rect 14829 24355 14887 24361
rect 16298 24352 16304 24404
rect 16356 24392 16362 24404
rect 16393 24395 16451 24401
rect 16393 24392 16405 24395
rect 16356 24364 16405 24392
rect 16356 24352 16362 24364
rect 16393 24361 16405 24364
rect 16439 24361 16451 24395
rect 16393 24355 16451 24361
rect 17681 24395 17739 24401
rect 17681 24361 17693 24395
rect 17727 24361 17739 24395
rect 17681 24355 17739 24361
rect 14553 24327 14611 24333
rect 14553 24293 14565 24327
rect 14599 24324 14611 24327
rect 14734 24324 14740 24336
rect 14599 24296 14740 24324
rect 14599 24293 14611 24296
rect 14553 24287 14611 24293
rect 14734 24284 14740 24296
rect 14792 24284 14798 24336
rect 15470 24284 15476 24336
rect 15528 24324 15534 24336
rect 17696 24324 17724 24355
rect 17862 24352 17868 24404
rect 17920 24352 17926 24404
rect 18322 24352 18328 24404
rect 18380 24352 18386 24404
rect 19978 24392 19984 24404
rect 19628 24364 19984 24392
rect 15528 24296 16257 24324
rect 15528 24284 15534 24296
rect 11422 24216 11428 24268
rect 11480 24256 11486 24268
rect 11793 24259 11851 24265
rect 11793 24256 11805 24259
rect 11480 24228 11805 24256
rect 11480 24216 11486 24228
rect 11793 24225 11805 24228
rect 11839 24225 11851 24259
rect 11793 24219 11851 24225
rect 13556 24228 13860 24256
rect 5000 24160 6500 24188
rect 7866 24160 8708 24188
rect 12529 24191 12587 24197
rect 3200 24092 4752 24120
rect 3200 24080 3206 24092
rect 4890 24012 4896 24064
rect 4948 24012 4954 24064
rect 6472 24052 6500 24160
rect 12529 24157 12541 24191
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 6730 24080 6736 24132
rect 6788 24080 6794 24132
rect 12544 24120 12572 24151
rect 12710 24148 12716 24200
rect 12768 24148 12774 24200
rect 12894 24148 12900 24200
rect 12952 24148 12958 24200
rect 13354 24148 13360 24200
rect 13412 24148 13418 24200
rect 13556 24178 13584 24228
rect 13832 24200 13860 24228
rect 14090 24216 14096 24268
rect 14148 24216 14154 24268
rect 14645 24259 14703 24265
rect 14645 24225 14657 24259
rect 14691 24256 14703 24259
rect 15102 24256 15108 24268
rect 14691 24228 15108 24256
rect 14691 24225 14703 24228
rect 14645 24219 14703 24225
rect 15102 24216 15108 24228
rect 15160 24216 15166 24268
rect 15396 24228 16160 24256
rect 15396 24200 15424 24228
rect 13633 24191 13691 24197
rect 13633 24178 13645 24191
rect 13556 24157 13645 24178
rect 13679 24157 13691 24191
rect 13556 24151 13691 24157
rect 13556 24150 13676 24151
rect 13814 24148 13820 24200
rect 13872 24148 13878 24200
rect 14182 24148 14188 24200
rect 14240 24188 14246 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 14240 24160 14289 24188
rect 14240 24148 14246 24160
rect 14277 24157 14289 24160
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 13722 24120 13728 24132
rect 12544 24092 13728 24120
rect 13722 24080 13728 24092
rect 13780 24120 13786 24132
rect 13998 24120 14004 24132
rect 13780 24092 14004 24120
rect 13780 24080 13786 24092
rect 13998 24080 14004 24092
rect 14056 24120 14062 24132
rect 14752 24120 14780 24151
rect 15286 24148 15292 24200
rect 15344 24148 15350 24200
rect 15378 24148 15384 24200
rect 15436 24148 15442 24200
rect 15746 24148 15752 24200
rect 15804 24148 15810 24200
rect 15842 24191 15900 24197
rect 15842 24157 15854 24191
rect 15888 24157 15900 24191
rect 15842 24151 15900 24157
rect 14056 24092 14780 24120
rect 14056 24080 14062 24092
rect 15856 24064 15884 24151
rect 16022 24148 16028 24200
rect 16080 24148 16086 24200
rect 16132 24197 16160 24228
rect 16229 24197 16257 24296
rect 16316 24296 17724 24324
rect 16316 24268 16344 24296
rect 16298 24216 16304 24268
rect 16356 24216 16362 24268
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 16942 24256 16948 24268
rect 16899 24228 16948 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17696 24256 17724 24296
rect 17696 24228 18276 24256
rect 16117 24191 16175 24197
rect 16117 24157 16129 24191
rect 16163 24157 16175 24191
rect 16117 24151 16175 24157
rect 16214 24191 16272 24197
rect 16214 24157 16226 24191
rect 16260 24157 16272 24191
rect 16214 24151 16272 24157
rect 16390 24148 16396 24200
rect 16448 24188 16454 24200
rect 16761 24191 16819 24197
rect 16761 24188 16773 24191
rect 16448 24160 16773 24188
rect 16448 24148 16454 24160
rect 16761 24157 16773 24160
rect 16807 24157 16819 24191
rect 16761 24151 16819 24157
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24188 17279 24191
rect 18046 24188 18052 24200
rect 17267 24160 18052 24188
rect 17267 24157 17279 24160
rect 17221 24151 17279 24157
rect 16776 24120 16804 24151
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18248 24197 18276 24228
rect 18340 24197 18368 24352
rect 18598 24284 18604 24336
rect 18656 24324 18662 24336
rect 19628 24333 19656 24364
rect 19978 24352 19984 24364
rect 20036 24392 20042 24404
rect 20036 24364 20668 24392
rect 20036 24352 20042 24364
rect 19613 24327 19671 24333
rect 19613 24324 19625 24327
rect 18656 24296 19625 24324
rect 18656 24284 18662 24296
rect 19613 24293 19625 24296
rect 19659 24293 19671 24327
rect 19613 24287 19671 24293
rect 20254 24284 20260 24336
rect 20312 24284 20318 24336
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 19058 24256 19064 24268
rect 18831 24228 19064 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 20272 24256 20300 24284
rect 19996 24228 20300 24256
rect 19996 24200 20024 24228
rect 20530 24216 20536 24268
rect 20588 24216 20594 24268
rect 20640 24256 20668 24364
rect 20990 24352 20996 24404
rect 21048 24392 21054 24404
rect 21266 24392 21272 24404
rect 21048 24364 21272 24392
rect 21048 24352 21054 24364
rect 21266 24352 21272 24364
rect 21324 24352 21330 24404
rect 21545 24395 21603 24401
rect 21545 24361 21557 24395
rect 21591 24392 21603 24395
rect 22094 24392 22100 24404
rect 21591 24364 22100 24392
rect 21591 24361 21603 24364
rect 21545 24355 21603 24361
rect 22094 24352 22100 24364
rect 22152 24352 22158 24404
rect 22646 24352 22652 24404
rect 22704 24392 22710 24404
rect 22741 24395 22799 24401
rect 22741 24392 22753 24395
rect 22704 24364 22753 24392
rect 22704 24352 22710 24364
rect 22741 24361 22753 24364
rect 22787 24361 22799 24395
rect 22741 24355 22799 24361
rect 24394 24352 24400 24404
rect 24452 24392 24458 24404
rect 24452 24364 25084 24392
rect 24452 24352 24458 24364
rect 22665 24296 22876 24324
rect 20993 24259 21051 24265
rect 20993 24256 21005 24259
rect 20640 24228 21005 24256
rect 20993 24225 21005 24228
rect 21039 24225 21051 24259
rect 20993 24219 21051 24225
rect 22002 24216 22008 24268
rect 22060 24256 22066 24268
rect 22665 24256 22693 24296
rect 22060 24228 22693 24256
rect 22060 24216 22066 24228
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24157 18291 24191
rect 18233 24151 18291 24157
rect 18325 24191 18383 24197
rect 18325 24157 18337 24191
rect 18371 24188 18383 24191
rect 19426 24188 19432 24200
rect 18371 24160 19432 24188
rect 18371 24157 18383 24160
rect 18325 24151 18383 24157
rect 17310 24120 17316 24132
rect 16776 24092 17316 24120
rect 17310 24080 17316 24092
rect 17368 24080 17374 24132
rect 17497 24123 17555 24129
rect 17497 24089 17509 24123
rect 17543 24120 17555 24123
rect 18156 24120 18184 24151
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 19978 24148 19984 24200
rect 20036 24148 20042 24200
rect 20438 24197 20444 24200
rect 20165 24191 20223 24197
rect 20165 24157 20177 24191
rect 20211 24188 20223 24191
rect 20257 24191 20315 24197
rect 20257 24188 20269 24191
rect 20211 24160 20269 24188
rect 20211 24157 20223 24160
rect 20165 24151 20223 24157
rect 20257 24157 20269 24160
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 20405 24191 20444 24197
rect 20405 24157 20417 24191
rect 20405 24151 20444 24157
rect 20438 24148 20444 24151
rect 20496 24148 20502 24200
rect 20548 24188 20576 24216
rect 20625 24191 20683 24197
rect 20625 24188 20637 24191
rect 20548 24160 20637 24188
rect 20625 24157 20637 24160
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 20763 24191 20821 24197
rect 20763 24157 20775 24191
rect 20809 24188 20821 24191
rect 21177 24191 21235 24197
rect 20809 24160 21128 24188
rect 20809 24157 20821 24160
rect 20763 24151 20821 24157
rect 17543 24092 18184 24120
rect 17543 24089 17555 24092
rect 17497 24083 17555 24089
rect 6914 24052 6920 24064
rect 6472 24024 6920 24052
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 7558 24012 7564 24064
rect 7616 24052 7622 24064
rect 8205 24055 8263 24061
rect 8205 24052 8217 24055
rect 7616 24024 8217 24052
rect 7616 24012 7622 24024
rect 8205 24021 8217 24024
rect 8251 24021 8263 24055
rect 8205 24015 8263 24021
rect 10134 24012 10140 24064
rect 10192 24052 10198 24064
rect 11238 24052 11244 24064
rect 10192 24024 11244 24052
rect 10192 24012 10198 24024
rect 11238 24012 11244 24024
rect 11296 24052 11302 24064
rect 11609 24055 11667 24061
rect 11609 24052 11621 24055
rect 11296 24024 11621 24052
rect 11296 24012 11302 24024
rect 11609 24021 11621 24024
rect 11655 24021 11667 24055
rect 11609 24015 11667 24021
rect 11701 24055 11759 24061
rect 11701 24021 11713 24055
rect 11747 24052 11759 24055
rect 12066 24052 12072 24064
rect 11747 24024 12072 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 12250 24012 12256 24064
rect 12308 24052 12314 24064
rect 15838 24052 15844 24064
rect 12308 24024 15844 24052
rect 12308 24012 12314 24024
rect 15838 24012 15844 24024
rect 15896 24012 15902 24064
rect 16850 24012 16856 24064
rect 16908 24052 16914 24064
rect 17681 24055 17739 24061
rect 17681 24052 17693 24055
rect 16908 24024 17693 24052
rect 16908 24012 16914 24024
rect 17681 24021 17693 24024
rect 17727 24021 17739 24055
rect 18156 24052 18184 24092
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 20533 24123 20591 24129
rect 19392 24092 19932 24120
rect 19392 24080 19398 24092
rect 18414 24052 18420 24064
rect 18156 24024 18420 24052
rect 17681 24015 17739 24021
rect 18414 24012 18420 24024
rect 18472 24012 18478 24064
rect 19242 24012 19248 24064
rect 19300 24052 19306 24064
rect 19904 24061 19932 24092
rect 20533 24089 20545 24123
rect 20579 24089 20591 24123
rect 21100 24120 21128 24160
rect 21177 24157 21189 24191
rect 21223 24188 21235 24191
rect 22094 24188 22100 24200
rect 21223 24160 22100 24188
rect 21223 24157 21235 24160
rect 21177 24151 21235 24157
rect 22094 24148 22100 24160
rect 22152 24188 22158 24200
rect 22554 24188 22560 24200
rect 22152 24160 22560 24188
rect 22152 24148 22158 24160
rect 22554 24148 22560 24160
rect 22612 24148 22618 24200
rect 22738 24148 22744 24200
rect 22796 24148 22802 24200
rect 22848 24197 22876 24296
rect 23382 24284 23388 24336
rect 23440 24324 23446 24336
rect 23477 24327 23535 24333
rect 23477 24324 23489 24327
rect 23440 24296 23489 24324
rect 23440 24284 23446 24296
rect 23477 24293 23489 24296
rect 23523 24293 23535 24327
rect 23477 24287 23535 24293
rect 24489 24327 24547 24333
rect 24489 24293 24501 24327
rect 24535 24324 24547 24327
rect 24854 24324 24860 24336
rect 24535 24296 24860 24324
rect 24535 24293 24547 24296
rect 24489 24287 24547 24293
rect 24854 24284 24860 24296
rect 24912 24284 24918 24336
rect 25056 24265 25084 24364
rect 25498 24352 25504 24404
rect 25556 24352 25562 24404
rect 26421 24395 26479 24401
rect 26421 24361 26433 24395
rect 26467 24392 26479 24395
rect 26694 24392 26700 24404
rect 26467 24364 26700 24392
rect 26467 24361 26479 24364
rect 26421 24355 26479 24361
rect 26694 24352 26700 24364
rect 26752 24352 26758 24404
rect 28261 24395 28319 24401
rect 28261 24361 28273 24395
rect 28307 24392 28319 24395
rect 28626 24392 28632 24404
rect 28307 24364 28632 24392
rect 28307 24361 28319 24364
rect 28261 24355 28319 24361
rect 28626 24352 28632 24364
rect 28684 24352 28690 24404
rect 28718 24352 28724 24404
rect 28776 24392 28782 24404
rect 30558 24392 30564 24404
rect 28776 24364 30564 24392
rect 28776 24352 28782 24364
rect 30558 24352 30564 24364
rect 30616 24352 30622 24404
rect 31389 24395 31447 24401
rect 31389 24392 31401 24395
rect 31220 24364 31401 24392
rect 25516 24324 25544 24352
rect 28902 24324 28908 24336
rect 25516 24296 25913 24324
rect 25041 24259 25099 24265
rect 25041 24225 25053 24259
rect 25087 24256 25099 24259
rect 25590 24256 25596 24268
rect 25087 24228 25596 24256
rect 25087 24225 25099 24228
rect 25041 24219 25099 24225
rect 25590 24216 25596 24228
rect 25648 24216 25654 24268
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24188 22891 24191
rect 23106 24188 23112 24200
rect 22879 24160 23112 24188
rect 22879 24157 22891 24160
rect 22833 24151 22891 24157
rect 23106 24148 23112 24160
rect 23164 24148 23170 24200
rect 24029 24191 24087 24197
rect 24029 24157 24041 24191
rect 24075 24188 24087 24191
rect 24762 24188 24768 24200
rect 24075 24160 24768 24188
rect 24075 24157 24087 24160
rect 24029 24151 24087 24157
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 25682 24148 25688 24200
rect 25740 24190 25746 24200
rect 25885 24197 25913 24296
rect 26896 24296 28908 24324
rect 26896 24268 26924 24296
rect 26878 24216 26884 24268
rect 26936 24216 26942 24268
rect 28736 24265 28764 24296
rect 28902 24284 28908 24296
rect 28960 24324 28966 24336
rect 29178 24324 29184 24336
rect 28960 24296 29184 24324
rect 28960 24284 28966 24296
rect 29178 24284 29184 24296
rect 29236 24284 29242 24336
rect 31018 24324 31024 24336
rect 30392 24296 31024 24324
rect 28721 24259 28779 24265
rect 27356 24228 27936 24256
rect 27356 24200 27384 24228
rect 25777 24191 25835 24197
rect 25777 24190 25789 24191
rect 25740 24162 25789 24190
rect 25740 24148 25746 24162
rect 25777 24157 25789 24162
rect 25823 24157 25835 24191
rect 25777 24151 25835 24157
rect 25870 24191 25928 24197
rect 25870 24157 25882 24191
rect 25916 24157 25928 24191
rect 25870 24151 25928 24157
rect 26283 24191 26341 24197
rect 26283 24157 26295 24191
rect 26329 24188 26341 24191
rect 26602 24188 26608 24200
rect 26329 24160 26608 24188
rect 26329 24157 26341 24160
rect 26283 24151 26341 24157
rect 26602 24148 26608 24160
rect 26660 24148 26666 24200
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24188 26755 24191
rect 26786 24188 26792 24200
rect 26743 24160 26792 24188
rect 26743 24157 26755 24160
rect 26697 24151 26755 24157
rect 26786 24148 26792 24160
rect 26844 24148 26850 24200
rect 27065 24191 27123 24197
rect 27065 24157 27077 24191
rect 27111 24188 27123 24191
rect 27338 24188 27344 24200
rect 27111 24160 27344 24188
rect 27111 24157 27123 24160
rect 27065 24151 27123 24157
rect 27338 24148 27344 24160
rect 27396 24148 27402 24200
rect 27709 24191 27767 24197
rect 27709 24157 27721 24191
rect 27755 24188 27767 24191
rect 27798 24188 27804 24200
rect 27755 24160 27804 24188
rect 27755 24157 27767 24160
rect 27709 24151 27767 24157
rect 27798 24148 27804 24160
rect 27856 24148 27862 24200
rect 27908 24197 27936 24228
rect 28721 24225 28733 24259
rect 28767 24225 28779 24259
rect 28721 24219 28779 24225
rect 28810 24216 28816 24268
rect 28868 24216 28874 24268
rect 30392 24256 30420 24296
rect 28966 24228 30420 24256
rect 27893 24191 27951 24197
rect 27893 24157 27905 24191
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 28169 24191 28227 24197
rect 28169 24157 28181 24191
rect 28215 24188 28227 24191
rect 28966 24188 28994 24228
rect 28215 24160 28994 24188
rect 28215 24157 28227 24160
rect 28169 24151 28227 24157
rect 30190 24148 30196 24200
rect 30248 24185 30254 24200
rect 30285 24191 30343 24197
rect 30285 24185 30297 24191
rect 30248 24157 30297 24185
rect 30331 24157 30343 24191
rect 30248 24148 30254 24157
rect 30285 24151 30343 24157
rect 30374 24148 30380 24200
rect 30432 24148 30438 24200
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24188 30527 24191
rect 30576 24188 30604 24296
rect 31018 24284 31024 24296
rect 31076 24284 31082 24336
rect 31220 24256 31248 24364
rect 31389 24361 31401 24364
rect 31435 24361 31447 24395
rect 31389 24355 31447 24361
rect 32858 24352 32864 24404
rect 32916 24392 32922 24404
rect 33229 24395 33287 24401
rect 33229 24392 33241 24395
rect 32916 24364 33241 24392
rect 32916 24352 32922 24364
rect 33229 24361 33241 24364
rect 33275 24361 33287 24395
rect 33229 24355 33287 24361
rect 32122 24284 32128 24336
rect 32180 24284 32186 24336
rect 32490 24284 32496 24336
rect 32548 24284 32554 24336
rect 30944 24228 31248 24256
rect 30515 24160 30604 24188
rect 30515 24157 30527 24160
rect 30469 24151 30527 24157
rect 30650 24148 30656 24200
rect 30708 24148 30714 24200
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24157 30803 24191
rect 30745 24151 30803 24157
rect 21634 24120 21640 24132
rect 21100 24092 21640 24120
rect 20533 24083 20591 24089
rect 19797 24055 19855 24061
rect 19797 24052 19809 24055
rect 19300 24024 19809 24052
rect 19300 24012 19306 24024
rect 19797 24021 19809 24024
rect 19843 24021 19855 24055
rect 19797 24015 19855 24021
rect 19889 24055 19947 24061
rect 19889 24021 19901 24055
rect 19935 24052 19947 24055
rect 20162 24052 20168 24064
rect 19935 24024 20168 24052
rect 19935 24021 19947 24024
rect 19889 24015 19947 24021
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 20548 24052 20576 24083
rect 21634 24080 21640 24092
rect 21692 24080 21698 24132
rect 22002 24080 22008 24132
rect 22060 24120 22066 24132
rect 23293 24123 23351 24129
rect 23293 24120 23305 24123
rect 22060 24092 23305 24120
rect 22060 24080 22066 24092
rect 23293 24089 23305 24092
rect 23339 24089 23351 24123
rect 23293 24083 23351 24089
rect 23750 24080 23756 24132
rect 23808 24120 23814 24132
rect 26053 24123 26111 24129
rect 26053 24120 26065 24123
rect 23808 24092 26065 24120
rect 23808 24080 23814 24092
rect 26053 24089 26065 24092
rect 26099 24089 26111 24123
rect 26053 24083 26111 24089
rect 26145 24123 26203 24129
rect 26145 24089 26157 24123
rect 26191 24089 26203 24123
rect 26145 24083 26203 24089
rect 20622 24052 20628 24064
rect 20548 24024 20628 24052
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 20898 24012 20904 24064
rect 20956 24012 20962 24064
rect 21266 24012 21272 24064
rect 21324 24012 21330 24064
rect 21358 24012 21364 24064
rect 21416 24012 21422 24064
rect 22186 24012 22192 24064
rect 22244 24052 22250 24064
rect 22738 24052 22744 24064
rect 22244 24024 22744 24052
rect 22244 24012 22250 24024
rect 22738 24012 22744 24024
rect 22796 24012 22802 24064
rect 23109 24055 23167 24061
rect 23109 24021 23121 24055
rect 23155 24052 23167 24055
rect 23382 24052 23388 24064
rect 23155 24024 23388 24052
rect 23155 24021 23167 24024
rect 23109 24015 23167 24021
rect 23382 24012 23388 24024
rect 23440 24012 23446 24064
rect 24118 24012 24124 24064
rect 24176 24012 24182 24064
rect 24762 24012 24768 24064
rect 24820 24052 24826 24064
rect 24857 24055 24915 24061
rect 24857 24052 24869 24055
rect 24820 24024 24869 24052
rect 24820 24012 24826 24024
rect 24857 24021 24869 24024
rect 24903 24021 24915 24055
rect 24857 24015 24915 24021
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 26160 24052 26188 24083
rect 26510 24080 26516 24132
rect 26568 24120 26574 24132
rect 26881 24123 26939 24129
rect 26881 24120 26893 24123
rect 26568 24092 26893 24120
rect 26568 24080 26574 24092
rect 26881 24089 26893 24092
rect 26927 24089 26939 24123
rect 26881 24083 26939 24089
rect 26970 24080 26976 24132
rect 27028 24080 27034 24132
rect 30760 24120 30788 24151
rect 30834 24148 30840 24200
rect 30892 24188 30898 24200
rect 30944 24197 30972 24228
rect 31220 24197 31248 24228
rect 31478 24216 31484 24268
rect 31536 24256 31542 24268
rect 32140 24256 32168 24284
rect 32309 24259 32367 24265
rect 32309 24256 32321 24259
rect 31536 24228 32321 24256
rect 31536 24216 31542 24228
rect 32309 24225 32321 24228
rect 32355 24225 32367 24259
rect 32309 24219 32367 24225
rect 32968 24228 34100 24256
rect 32968 24200 32996 24228
rect 30929 24191 30987 24197
rect 30929 24188 30941 24191
rect 30892 24160 30941 24188
rect 30892 24148 30898 24160
rect 30929 24157 30941 24160
rect 30975 24157 30987 24191
rect 30929 24151 30987 24157
rect 31021 24191 31079 24197
rect 31021 24157 31033 24191
rect 31067 24157 31079 24191
rect 31021 24151 31079 24157
rect 31205 24191 31263 24197
rect 31205 24157 31217 24191
rect 31251 24157 31263 24191
rect 31205 24151 31263 24157
rect 31297 24191 31355 24197
rect 31297 24157 31309 24191
rect 31343 24157 31355 24191
rect 31297 24151 31355 24157
rect 31036 24120 31064 24151
rect 31312 24120 31340 24151
rect 32030 24148 32036 24200
rect 32088 24148 32094 24200
rect 32122 24148 32128 24200
rect 32180 24148 32186 24200
rect 32398 24148 32404 24200
rect 32456 24148 32462 24200
rect 32493 24191 32551 24197
rect 32493 24157 32505 24191
rect 32539 24188 32551 24191
rect 32582 24188 32588 24200
rect 32539 24160 32588 24188
rect 32539 24157 32551 24160
rect 32493 24151 32551 24157
rect 32582 24148 32588 24160
rect 32640 24148 32646 24200
rect 32769 24191 32827 24197
rect 32769 24157 32781 24191
rect 32815 24188 32827 24191
rect 32861 24191 32919 24197
rect 32861 24188 32873 24191
rect 32815 24160 32873 24188
rect 32815 24157 32827 24160
rect 32769 24151 32827 24157
rect 32861 24157 32873 24160
rect 32907 24157 32919 24191
rect 32861 24151 32919 24157
rect 32784 24120 32812 24151
rect 32950 24148 32956 24200
rect 33008 24148 33014 24200
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24157 33195 24191
rect 33137 24151 33195 24157
rect 33152 24120 33180 24151
rect 33870 24148 33876 24200
rect 33928 24148 33934 24200
rect 33962 24148 33968 24200
rect 34020 24148 34026 24200
rect 34072 24188 34100 24228
rect 34238 24216 34244 24268
rect 34296 24256 34302 24268
rect 34296 24228 34376 24256
rect 34296 24216 34302 24228
rect 34348 24197 34376 24228
rect 34333 24191 34391 24197
rect 34072 24160 34284 24188
rect 27264 24092 31340 24120
rect 31772 24092 32812 24120
rect 32876 24092 33180 24120
rect 33888 24120 33916 24148
rect 34256 24129 34284 24160
rect 34333 24157 34345 24191
rect 34379 24188 34391 24191
rect 34793 24191 34851 24197
rect 34793 24188 34805 24191
rect 34379 24160 34805 24188
rect 34379 24157 34391 24160
rect 34333 24151 34391 24157
rect 34793 24157 34805 24160
rect 34839 24157 34851 24191
rect 34793 24151 34851 24157
rect 34977 24191 35035 24197
rect 34977 24157 34989 24191
rect 35023 24157 35035 24191
rect 34977 24151 35035 24157
rect 34149 24123 34207 24129
rect 34149 24120 34161 24123
rect 33888 24092 34161 24120
rect 26234 24052 26240 24064
rect 25004 24024 26240 24052
rect 25004 24012 25010 24024
rect 26234 24012 26240 24024
rect 26292 24012 26298 24064
rect 27264 24061 27292 24092
rect 27249 24055 27307 24061
rect 27249 24021 27261 24055
rect 27295 24021 27307 24055
rect 27249 24015 27307 24021
rect 27614 24012 27620 24064
rect 27672 24052 27678 24064
rect 28534 24052 28540 24064
rect 27672 24024 28540 24052
rect 27672 24012 27678 24024
rect 28534 24012 28540 24024
rect 28592 24052 28598 24064
rect 28629 24055 28687 24061
rect 28629 24052 28641 24055
rect 28592 24024 28641 24052
rect 28592 24012 28598 24024
rect 28629 24021 28641 24024
rect 28675 24021 28687 24055
rect 28629 24015 28687 24021
rect 30009 24055 30067 24061
rect 30009 24021 30021 24055
rect 30055 24052 30067 24055
rect 30742 24052 30748 24064
rect 30055 24024 30748 24052
rect 30055 24021 30067 24024
rect 30009 24015 30067 24021
rect 30742 24012 30748 24024
rect 30800 24012 30806 24064
rect 30834 24012 30840 24064
rect 30892 24012 30898 24064
rect 31202 24012 31208 24064
rect 31260 24012 31266 24064
rect 31772 24061 31800 24092
rect 31757 24055 31815 24061
rect 31757 24021 31769 24055
rect 31803 24021 31815 24055
rect 31757 24015 31815 24021
rect 31846 24012 31852 24064
rect 31904 24012 31910 24064
rect 32214 24012 32220 24064
rect 32272 24052 32278 24064
rect 32677 24055 32735 24061
rect 32677 24052 32689 24055
rect 32272 24024 32689 24052
rect 32272 24012 32278 24024
rect 32677 24021 32689 24024
rect 32723 24052 32735 24055
rect 32876 24052 32904 24092
rect 34149 24089 34161 24092
rect 34195 24089 34207 24123
rect 34149 24083 34207 24089
rect 34241 24123 34299 24129
rect 34241 24089 34253 24123
rect 34287 24120 34299 24123
rect 34992 24120 35020 24151
rect 35066 24120 35072 24132
rect 34287 24092 35072 24120
rect 34287 24089 34299 24092
rect 34241 24083 34299 24089
rect 35066 24080 35072 24092
rect 35124 24080 35130 24132
rect 32723 24024 32904 24052
rect 32723 24021 32735 24024
rect 32677 24015 32735 24021
rect 32950 24012 32956 24064
rect 33008 24012 33014 24064
rect 34514 24012 34520 24064
rect 34572 24012 34578 24064
rect 34698 24012 34704 24064
rect 34756 24052 34762 24064
rect 35805 24055 35863 24061
rect 35805 24052 35817 24055
rect 34756 24024 35817 24052
rect 34756 24012 34762 24024
rect 35805 24021 35817 24024
rect 35851 24021 35863 24055
rect 35805 24015 35863 24021
rect 1104 23962 38272 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38272 23962
rect 1104 23888 38272 23910
rect 6730 23808 6736 23860
rect 6788 23848 6794 23860
rect 6917 23851 6975 23857
rect 6917 23848 6929 23851
rect 6788 23820 6929 23848
rect 6788 23808 6794 23820
rect 6917 23817 6929 23820
rect 6963 23817 6975 23851
rect 6917 23811 6975 23817
rect 7193 23851 7251 23857
rect 7193 23817 7205 23851
rect 7239 23817 7251 23851
rect 7193 23811 7251 23817
rect 1670 23780 1676 23792
rect 1412 23752 1676 23780
rect 1412 23721 1440 23752
rect 1670 23740 1676 23752
rect 1728 23740 1734 23792
rect 4062 23780 4068 23792
rect 2898 23752 4068 23780
rect 4062 23740 4068 23752
rect 4120 23740 4126 23792
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 7101 23715 7159 23721
rect 7101 23681 7113 23715
rect 7147 23712 7159 23715
rect 7208 23712 7236 23811
rect 10318 23808 10324 23860
rect 10376 23848 10382 23860
rect 10781 23851 10839 23857
rect 10781 23848 10793 23851
rect 10376 23820 10793 23848
rect 10376 23808 10382 23820
rect 10781 23817 10793 23820
rect 10827 23817 10839 23851
rect 10781 23811 10839 23817
rect 12710 23808 12716 23860
rect 12768 23808 12774 23860
rect 13354 23848 13360 23860
rect 12912 23820 13360 23848
rect 11606 23780 11612 23792
rect 7147 23684 7236 23712
rect 7484 23752 7788 23780
rect 7147 23681 7159 23684
rect 7101 23675 7159 23681
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23644 1731 23647
rect 1762 23644 1768 23656
rect 1719 23616 1768 23644
rect 1719 23613 1731 23616
rect 1673 23607 1731 23613
rect 1762 23604 1768 23616
rect 1820 23604 1826 23656
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 7484 23644 7512 23752
rect 7558 23672 7564 23724
rect 7616 23672 7622 23724
rect 6972 23616 7512 23644
rect 6972 23604 6978 23616
rect 7650 23604 7656 23656
rect 7708 23604 7714 23656
rect 7760 23653 7788 23752
rect 10704 23752 11612 23780
rect 10704 23721 10732 23752
rect 11606 23740 11612 23752
rect 11664 23740 11670 23792
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 10689 23715 10747 23721
rect 10689 23681 10701 23715
rect 10735 23681 10747 23715
rect 10689 23675 10747 23681
rect 7745 23647 7803 23653
rect 7745 23613 7757 23647
rect 7791 23613 7803 23647
rect 10520 23644 10548 23675
rect 10778 23672 10784 23724
rect 10836 23712 10842 23724
rect 10873 23715 10931 23721
rect 10873 23712 10885 23715
rect 10836 23684 10885 23712
rect 10836 23672 10842 23684
rect 10873 23681 10885 23684
rect 10919 23712 10931 23715
rect 11422 23712 11428 23724
rect 10919 23684 11428 23712
rect 10919 23681 10931 23684
rect 10873 23675 10931 23681
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11514 23644 11520 23656
rect 10520 23616 11520 23644
rect 7745 23607 7803 23613
rect 11514 23604 11520 23616
rect 11572 23604 11578 23656
rect 12728 23644 12756 23808
rect 12912 23789 12940 23820
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 13817 23851 13875 23857
rect 13817 23848 13829 23851
rect 13556 23820 13829 23848
rect 13556 23792 13584 23820
rect 13817 23817 13829 23820
rect 13863 23817 13875 23851
rect 13817 23811 13875 23817
rect 13906 23808 13912 23860
rect 13964 23848 13970 23860
rect 14093 23851 14151 23857
rect 14093 23848 14105 23851
rect 13964 23820 14105 23848
rect 13964 23808 13970 23820
rect 14093 23817 14105 23820
rect 14139 23817 14151 23851
rect 14093 23811 14151 23817
rect 14458 23808 14464 23860
rect 14516 23848 14522 23860
rect 18322 23848 18328 23860
rect 14516 23820 18328 23848
rect 14516 23808 14522 23820
rect 12897 23783 12955 23789
rect 12897 23749 12909 23783
rect 12943 23749 12955 23783
rect 12897 23743 12955 23749
rect 13262 23740 13268 23792
rect 13320 23740 13326 23792
rect 13538 23740 13544 23792
rect 13596 23740 13602 23792
rect 15286 23780 15292 23792
rect 13648 23752 15292 23780
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13354 23712 13360 23724
rect 13127 23684 13360 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 13354 23672 13360 23684
rect 13412 23672 13418 23724
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 13648 23712 13676 23752
rect 13495 23684 13676 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 13722 23672 13728 23724
rect 13780 23672 13786 23724
rect 13832 23712 13860 23752
rect 14292 23724 14320 23752
rect 15286 23740 15292 23752
rect 15344 23740 15350 23792
rect 15930 23740 15936 23792
rect 15988 23780 15994 23792
rect 15988 23752 16160 23780
rect 15988 23740 15994 23752
rect 13903 23715 13961 23721
rect 13903 23712 13915 23715
rect 13832 23684 13915 23712
rect 13903 23681 13915 23684
rect 13949 23681 13961 23715
rect 13903 23675 13961 23681
rect 13998 23672 14004 23724
rect 14056 23672 14062 23724
rect 14185 23715 14243 23721
rect 14185 23681 14197 23715
rect 14231 23681 14243 23715
rect 14185 23675 14243 23681
rect 13541 23647 13599 23653
rect 13541 23644 13553 23647
rect 12728 23616 13553 23644
rect 13541 23613 13553 23616
rect 13587 23644 13599 23647
rect 14200 23644 14228 23675
rect 14274 23672 14280 23724
rect 14332 23672 14338 23724
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15838 23712 15844 23724
rect 15252 23684 15844 23712
rect 15252 23672 15258 23684
rect 15838 23672 15844 23684
rect 15896 23672 15902 23724
rect 16132 23721 16160 23752
rect 16224 23721 16252 23820
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 18417 23851 18475 23857
rect 18417 23817 18429 23851
rect 18463 23848 18475 23851
rect 18506 23848 18512 23860
rect 18463 23820 18512 23848
rect 18463 23817 18475 23820
rect 18417 23811 18475 23817
rect 18506 23808 18512 23820
rect 18564 23848 18570 23860
rect 22094 23848 22100 23860
rect 18564 23820 22100 23848
rect 18564 23808 18570 23820
rect 22094 23808 22100 23820
rect 22152 23808 22158 23860
rect 22186 23808 22192 23860
rect 22244 23848 22250 23860
rect 22244 23820 23336 23848
rect 22244 23808 22250 23820
rect 17144 23752 18184 23780
rect 17144 23721 17172 23752
rect 16025 23715 16083 23721
rect 16025 23681 16037 23715
rect 16071 23681 16083 23715
rect 16025 23675 16083 23681
rect 16117 23715 16175 23721
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 16209 23715 16267 23721
rect 16209 23681 16221 23715
rect 16255 23681 16267 23715
rect 17129 23715 17187 23721
rect 17129 23712 17141 23715
rect 16209 23675 16267 23681
rect 16684 23684 17141 23712
rect 13587 23616 14228 23644
rect 13587 23613 13599 23616
rect 13541 23607 13599 23613
rect 15562 23604 15568 23656
rect 15620 23644 15626 23656
rect 16040 23644 16068 23675
rect 15620 23616 16068 23644
rect 15620 23604 15626 23616
rect 7098 23536 7104 23588
rect 7156 23576 7162 23588
rect 13906 23576 13912 23588
rect 7156 23548 13912 23576
rect 7156 23536 7162 23548
rect 13906 23536 13912 23548
rect 13964 23536 13970 23588
rect 16114 23536 16120 23588
rect 16172 23536 16178 23588
rect 16206 23536 16212 23588
rect 16264 23576 16270 23588
rect 16684 23576 16712 23684
rect 17129 23681 17141 23684
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23681 17371 23715
rect 17313 23675 17371 23681
rect 17034 23604 17040 23656
rect 17092 23644 17098 23656
rect 17328 23644 17356 23675
rect 17402 23672 17408 23724
rect 17460 23712 17466 23724
rect 18156 23721 18184 23752
rect 18524 23752 19334 23780
rect 18524 23724 18552 23752
rect 17497 23715 17555 23721
rect 17497 23712 17509 23715
rect 17460 23684 17509 23712
rect 17460 23672 17466 23684
rect 17497 23681 17509 23684
rect 17543 23681 17555 23715
rect 17497 23675 17555 23681
rect 18141 23715 18199 23721
rect 18141 23681 18153 23715
rect 18187 23681 18199 23715
rect 18141 23675 18199 23681
rect 18414 23672 18420 23724
rect 18472 23672 18478 23724
rect 18506 23672 18512 23724
rect 18564 23672 18570 23724
rect 18598 23672 18604 23724
rect 18656 23672 18662 23724
rect 17092 23616 17356 23644
rect 19306 23644 19334 23752
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 20346 23780 20352 23792
rect 19484 23752 20352 23780
rect 19484 23740 19490 23752
rect 20346 23740 20352 23752
rect 20404 23780 20410 23792
rect 21358 23780 21364 23792
rect 20404 23752 21364 23780
rect 20404 23740 20410 23752
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 21468 23752 22508 23780
rect 21468 23724 21496 23752
rect 20530 23672 20536 23724
rect 20588 23712 20594 23724
rect 20806 23712 20812 23724
rect 20588 23684 20812 23712
rect 20588 23672 20594 23684
rect 20806 23672 20812 23684
rect 20864 23672 20870 23724
rect 21450 23672 21456 23724
rect 21508 23672 21514 23724
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 22480 23721 22508 23752
rect 22572 23721 22600 23820
rect 22738 23740 22744 23792
rect 22796 23780 22802 23792
rect 23106 23780 23112 23792
rect 22796 23752 23112 23780
rect 22796 23740 22802 23752
rect 23106 23740 23112 23752
rect 23164 23740 23170 23792
rect 22281 23715 22339 23721
rect 22281 23712 22293 23715
rect 21784 23684 22293 23712
rect 21784 23672 21790 23684
rect 22281 23681 22293 23684
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 22465 23715 22523 23721
rect 22465 23681 22477 23715
rect 22511 23681 22523 23715
rect 22465 23675 22523 23681
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 19429 23647 19487 23653
rect 19429 23644 19441 23647
rect 19306 23616 19441 23644
rect 17092 23604 17098 23616
rect 19429 23613 19441 23616
rect 19475 23644 19487 23647
rect 21818 23644 21824 23656
rect 19475 23616 21824 23644
rect 19475 23613 19487 23616
rect 19429 23607 19487 23613
rect 21818 23604 21824 23616
rect 21876 23604 21882 23656
rect 22480 23644 22508 23675
rect 22646 23672 22652 23724
rect 22704 23712 22710 23724
rect 23017 23715 23075 23721
rect 22704 23684 22749 23712
rect 22704 23672 22710 23684
rect 23017 23681 23029 23715
rect 23063 23712 23075 23715
rect 23124 23712 23152 23740
rect 23308 23721 23336 23820
rect 23382 23808 23388 23860
rect 23440 23808 23446 23860
rect 26053 23851 26111 23857
rect 24044 23820 26004 23848
rect 23400 23780 23428 23808
rect 24044 23789 24072 23820
rect 24029 23783 24087 23789
rect 23400 23752 23796 23780
rect 23063 23684 23152 23712
rect 23201 23715 23259 23721
rect 23063 23681 23075 23684
rect 23017 23675 23075 23681
rect 23201 23681 23213 23715
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 23293 23715 23351 23721
rect 23293 23681 23305 23715
rect 23339 23681 23351 23715
rect 23293 23675 23351 23681
rect 23386 23715 23444 23721
rect 23386 23681 23398 23715
rect 23432 23681 23444 23715
rect 23386 23675 23444 23681
rect 23216 23644 23244 23675
rect 22480 23616 23244 23644
rect 16264 23548 16712 23576
rect 16945 23579 17003 23585
rect 16264 23536 16270 23548
rect 16945 23545 16957 23579
rect 16991 23576 17003 23579
rect 17218 23576 17224 23588
rect 16991 23548 17224 23576
rect 16991 23545 17003 23548
rect 16945 23539 17003 23545
rect 17218 23536 17224 23548
rect 17276 23576 17282 23588
rect 21266 23576 21272 23588
rect 17276 23548 21272 23576
rect 17276 23536 17282 23548
rect 21266 23536 21272 23548
rect 21324 23536 21330 23588
rect 21910 23576 21916 23588
rect 21560 23548 21916 23576
rect 3145 23511 3203 23517
rect 3145 23477 3157 23511
rect 3191 23508 3203 23511
rect 3326 23508 3332 23520
rect 3191 23480 3332 23508
rect 3191 23477 3203 23480
rect 3145 23471 3203 23477
rect 3326 23468 3332 23480
rect 3384 23468 3390 23520
rect 10226 23468 10232 23520
rect 10284 23508 10290 23520
rect 10321 23511 10379 23517
rect 10321 23508 10333 23511
rect 10284 23480 10333 23508
rect 10284 23468 10290 23480
rect 10321 23477 10333 23480
rect 10367 23477 10379 23511
rect 10321 23471 10379 23477
rect 13354 23468 13360 23520
rect 13412 23508 13418 23520
rect 13630 23508 13636 23520
rect 13412 23480 13636 23508
rect 13412 23468 13418 23480
rect 13630 23468 13636 23480
rect 13688 23508 13694 23520
rect 14182 23508 14188 23520
rect 13688 23480 14188 23508
rect 13688 23468 13694 23480
rect 14182 23468 14188 23480
rect 14240 23468 14246 23520
rect 16132 23508 16160 23536
rect 16393 23511 16451 23517
rect 16393 23508 16405 23511
rect 16132 23480 16405 23508
rect 16393 23477 16405 23480
rect 16439 23477 16451 23511
rect 16393 23471 16451 23477
rect 18138 23468 18144 23520
rect 18196 23508 18202 23520
rect 18966 23508 18972 23520
rect 18196 23480 18972 23508
rect 18196 23468 18202 23480
rect 18966 23468 18972 23480
rect 19024 23468 19030 23520
rect 19242 23468 19248 23520
rect 19300 23508 19306 23520
rect 21560 23508 21588 23548
rect 21910 23536 21916 23548
rect 21968 23536 21974 23588
rect 22925 23579 22983 23585
rect 22925 23545 22937 23579
rect 22971 23576 22983 23579
rect 23014 23576 23020 23588
rect 22971 23548 23020 23576
rect 22971 23545 22983 23548
rect 22925 23539 22983 23545
rect 23014 23536 23020 23548
rect 23072 23536 23078 23588
rect 23106 23536 23112 23588
rect 23164 23576 23170 23588
rect 23400 23576 23428 23675
rect 23566 23672 23572 23724
rect 23624 23712 23630 23724
rect 23768 23721 23796 23752
rect 24029 23749 24041 23783
rect 24075 23749 24087 23783
rect 24029 23743 24087 23749
rect 25314 23740 25320 23792
rect 25372 23740 25378 23792
rect 25976 23780 26004 23820
rect 26053 23817 26065 23851
rect 26099 23848 26111 23851
rect 26234 23848 26240 23860
rect 26099 23820 26240 23848
rect 26099 23817 26111 23820
rect 26053 23811 26111 23817
rect 26234 23808 26240 23820
rect 26292 23808 26298 23860
rect 28718 23848 28724 23860
rect 26436 23820 28724 23848
rect 26436 23780 26464 23820
rect 28718 23808 28724 23820
rect 28776 23808 28782 23860
rect 29178 23808 29184 23860
rect 29236 23848 29242 23860
rect 29825 23851 29883 23857
rect 29825 23848 29837 23851
rect 29236 23820 29837 23848
rect 29236 23808 29242 23820
rect 29825 23817 29837 23820
rect 29871 23817 29883 23851
rect 29825 23811 29883 23817
rect 30834 23808 30840 23860
rect 30892 23808 30898 23860
rect 31757 23851 31815 23857
rect 31757 23817 31769 23851
rect 31803 23848 31815 23851
rect 32122 23848 32128 23860
rect 31803 23820 32128 23848
rect 31803 23817 31815 23820
rect 31757 23811 31815 23817
rect 32122 23808 32128 23820
rect 32180 23808 32186 23860
rect 32306 23808 32312 23860
rect 32364 23808 32370 23860
rect 32398 23808 32404 23860
rect 32456 23808 32462 23860
rect 34514 23808 34520 23860
rect 34572 23808 34578 23860
rect 35342 23808 35348 23860
rect 35400 23808 35406 23860
rect 25976 23752 26464 23780
rect 26510 23740 26516 23792
rect 26568 23780 26574 23792
rect 27157 23783 27215 23789
rect 27157 23780 27169 23783
rect 26568 23752 27169 23780
rect 26568 23740 26574 23752
rect 27157 23749 27169 23752
rect 27203 23749 27215 23783
rect 27157 23743 27215 23749
rect 27982 23740 27988 23792
rect 28040 23740 28046 23792
rect 28258 23740 28264 23792
rect 28316 23780 28322 23792
rect 28353 23783 28411 23789
rect 28353 23780 28365 23783
rect 28316 23752 28365 23780
rect 28316 23740 28322 23752
rect 28353 23749 28365 23752
rect 28399 23749 28411 23783
rect 29638 23780 29644 23792
rect 29578 23752 29644 23780
rect 28353 23743 28411 23749
rect 29638 23740 29644 23752
rect 29696 23740 29702 23792
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23624 23684 23673 23712
rect 23624 23672 23630 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 23753 23715 23811 23721
rect 23753 23681 23765 23715
rect 23799 23681 23811 23715
rect 23753 23675 23811 23681
rect 24118 23672 24124 23724
rect 24176 23712 24182 23724
rect 24305 23715 24363 23721
rect 24305 23712 24317 23715
rect 24176 23684 24317 23712
rect 24176 23672 24182 23684
rect 24305 23681 24317 23684
rect 24351 23681 24363 23715
rect 24305 23675 24363 23681
rect 26973 23715 27031 23721
rect 26973 23681 26985 23715
rect 27019 23712 27031 23715
rect 27062 23712 27068 23724
rect 27019 23684 27068 23712
rect 27019 23681 27031 23684
rect 26973 23675 27031 23681
rect 27062 23672 27068 23684
rect 27120 23672 27126 23724
rect 27246 23672 27252 23724
rect 27304 23672 27310 23724
rect 27338 23672 27344 23724
rect 27396 23672 27402 23724
rect 27614 23712 27620 23724
rect 27448 23684 27620 23712
rect 23934 23604 23940 23656
rect 23992 23604 23998 23656
rect 24578 23604 24584 23656
rect 24636 23604 24642 23656
rect 24670 23604 24676 23656
rect 24728 23644 24734 23656
rect 27448 23644 27476 23684
rect 27614 23672 27620 23684
rect 27672 23672 27678 23724
rect 28000 23712 28028 23740
rect 28077 23715 28135 23721
rect 28077 23712 28089 23715
rect 28000 23684 28089 23712
rect 28077 23681 28089 23684
rect 28123 23681 28135 23715
rect 30852 23712 30880 23808
rect 31018 23740 31024 23792
rect 31076 23780 31082 23792
rect 31076 23752 32260 23780
rect 31076 23740 31082 23752
rect 31665 23715 31723 23721
rect 31665 23712 31677 23715
rect 30852 23684 31677 23712
rect 28077 23675 28135 23681
rect 31665 23681 31677 23684
rect 31711 23681 31723 23715
rect 31665 23675 31723 23681
rect 31478 23644 31484 23656
rect 24728 23616 27476 23644
rect 27540 23616 31484 23644
rect 24728 23604 24734 23616
rect 23164 23548 23428 23576
rect 23164 23536 23170 23548
rect 19300 23480 21588 23508
rect 19300 23468 19306 23480
rect 21634 23468 21640 23520
rect 21692 23508 21698 23520
rect 22370 23508 22376 23520
rect 21692 23480 22376 23508
rect 21692 23468 21698 23480
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 22646 23468 22652 23520
rect 22704 23508 22710 23520
rect 23952 23508 23980 23604
rect 27540 23585 27568 23616
rect 31478 23604 31484 23616
rect 31536 23604 31542 23656
rect 32232 23644 32260 23752
rect 32324 23721 32352 23808
rect 32309 23715 32367 23721
rect 32309 23681 32321 23715
rect 32355 23681 32367 23715
rect 34532 23712 34560 23808
rect 35360 23721 35388 23808
rect 34793 23715 34851 23721
rect 34793 23712 34805 23715
rect 34532 23684 34805 23712
rect 32309 23675 32367 23681
rect 34793 23681 34805 23684
rect 34839 23681 34851 23715
rect 35161 23715 35219 23721
rect 35161 23712 35173 23715
rect 34793 23675 34851 23681
rect 34992 23684 35173 23712
rect 33962 23644 33968 23656
rect 32232 23616 33968 23644
rect 33962 23604 33968 23616
rect 34020 23604 34026 23656
rect 34992 23653 35020 23684
rect 35161 23681 35173 23684
rect 35207 23681 35219 23715
rect 35161 23675 35219 23681
rect 35345 23715 35403 23721
rect 35345 23681 35357 23715
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 34977 23647 35035 23653
rect 34977 23644 34989 23647
rect 34256 23616 34989 23644
rect 27525 23579 27583 23585
rect 27525 23545 27537 23579
rect 27571 23545 27583 23579
rect 27525 23539 27583 23545
rect 31110 23536 31116 23588
rect 31168 23576 31174 23588
rect 33226 23576 33232 23588
rect 31168 23548 33232 23576
rect 31168 23536 31174 23548
rect 33226 23536 33232 23548
rect 33284 23536 33290 23588
rect 34256 23520 34284 23616
rect 34977 23613 34989 23616
rect 35023 23613 35035 23647
rect 34977 23607 35035 23613
rect 35066 23604 35072 23656
rect 35124 23604 35130 23656
rect 34790 23536 34796 23588
rect 34848 23576 34854 23588
rect 35161 23579 35219 23585
rect 35161 23576 35173 23579
rect 34848 23548 35173 23576
rect 34848 23536 34854 23548
rect 35161 23545 35173 23548
rect 35207 23545 35219 23579
rect 35161 23539 35219 23545
rect 22704 23480 23980 23508
rect 22704 23468 22710 23480
rect 25590 23468 25596 23520
rect 25648 23508 25654 23520
rect 32766 23508 32772 23520
rect 25648 23480 32772 23508
rect 25648 23468 25654 23480
rect 32766 23468 32772 23480
rect 32824 23468 32830 23520
rect 34238 23468 34244 23520
rect 34296 23468 34302 23520
rect 34606 23468 34612 23520
rect 34664 23468 34670 23520
rect 1104 23418 38272 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38272 23418
rect 1104 23344 38272 23366
rect 1762 23264 1768 23316
rect 1820 23264 1826 23316
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 3789 23307 3847 23313
rect 3789 23304 3801 23307
rect 2924 23276 3801 23304
rect 2924 23264 2930 23276
rect 3789 23273 3801 23276
rect 3835 23273 3847 23307
rect 3789 23267 3847 23273
rect 4356 23276 6132 23304
rect 2961 23171 3019 23177
rect 2961 23137 2973 23171
rect 3007 23168 3019 23171
rect 3142 23168 3148 23180
rect 3007 23140 3148 23168
rect 3007 23137 3019 23140
rect 2961 23131 3019 23137
rect 3142 23128 3148 23140
rect 3200 23128 3206 23180
rect 1949 23103 2007 23109
rect 1949 23069 1961 23103
rect 1995 23100 2007 23103
rect 2685 23103 2743 23109
rect 1995 23072 2360 23100
rect 1995 23069 2007 23072
rect 1949 23063 2007 23069
rect 2332 22973 2360 23072
rect 2685 23069 2697 23103
rect 2731 23100 2743 23103
rect 3326 23100 3332 23112
rect 2731 23072 3332 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 3326 23060 3332 23072
rect 3384 23060 3390 23112
rect 3970 23060 3976 23112
rect 4028 23060 4034 23112
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4356 23100 4384 23276
rect 6104 23236 6132 23276
rect 7650 23264 7656 23316
rect 7708 23304 7714 23316
rect 8021 23307 8079 23313
rect 8021 23304 8033 23307
rect 7708 23276 8033 23304
rect 7708 23264 7714 23276
rect 8021 23273 8033 23276
rect 8067 23273 8079 23307
rect 8021 23267 8079 23273
rect 8110 23264 8116 23316
rect 8168 23304 8174 23316
rect 8168 23276 14136 23304
rect 8168 23264 8174 23276
rect 6362 23236 6368 23248
rect 6104 23208 6368 23236
rect 4798 23128 4804 23180
rect 4856 23168 4862 23180
rect 5442 23168 5448 23180
rect 4856 23140 5448 23168
rect 4856 23128 4862 23140
rect 5442 23128 5448 23140
rect 5500 23128 5506 23180
rect 5626 23128 5632 23180
rect 5684 23168 5690 23180
rect 6104 23168 6132 23208
rect 6362 23196 6368 23208
rect 6420 23236 6426 23248
rect 7282 23236 7288 23248
rect 6420 23208 7288 23236
rect 6420 23196 6426 23208
rect 7282 23196 7288 23208
rect 7340 23236 7346 23248
rect 7340 23208 8432 23236
rect 7340 23196 7346 23208
rect 5684 23140 6132 23168
rect 5684 23128 5690 23140
rect 6914 23128 6920 23180
rect 6972 23168 6978 23180
rect 7193 23171 7251 23177
rect 7193 23168 7205 23171
rect 6972 23140 7205 23168
rect 6972 23128 6978 23140
rect 7193 23137 7205 23140
rect 7239 23137 7251 23171
rect 7193 23131 7251 23137
rect 4212 23072 4384 23100
rect 4433 23103 4491 23109
rect 4212 23060 4218 23072
rect 4433 23069 4445 23103
rect 4479 23100 4491 23103
rect 4614 23100 4620 23112
rect 4479 23072 4620 23100
rect 4479 23069 4491 23072
rect 4433 23063 4491 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 6178 23060 6184 23112
rect 6236 23060 6242 23112
rect 8404 23109 8432 23208
rect 9398 23196 9404 23248
rect 9456 23196 9462 23248
rect 11330 23196 11336 23248
rect 11388 23196 11394 23248
rect 13722 23196 13728 23248
rect 13780 23196 13786 23248
rect 13814 23196 13820 23248
rect 13872 23196 13878 23248
rect 14108 23236 14136 23276
rect 14182 23264 14188 23316
rect 14240 23304 14246 23316
rect 15381 23307 15439 23313
rect 15381 23304 15393 23307
rect 14240 23276 15393 23304
rect 14240 23264 14246 23276
rect 15381 23273 15393 23276
rect 15427 23273 15439 23307
rect 16942 23304 16948 23316
rect 15381 23267 15439 23273
rect 16040 23276 16948 23304
rect 16040 23248 16068 23276
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 17681 23307 17739 23313
rect 17681 23273 17693 23307
rect 17727 23273 17739 23307
rect 17681 23267 17739 23273
rect 17865 23307 17923 23313
rect 17865 23273 17877 23307
rect 17911 23304 17923 23307
rect 18598 23304 18604 23316
rect 17911 23276 18604 23304
rect 17911 23273 17923 23276
rect 17865 23267 17923 23273
rect 14108 23208 15240 23236
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23069 8263 23103
rect 8205 23063 8263 23069
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23069 8447 23103
rect 8389 23063 8447 23069
rect 3602 22992 3608 23044
rect 3660 23032 3666 23044
rect 4338 23041 4344 23044
rect 4065 23035 4123 23041
rect 4065 23032 4077 23035
rect 3660 23004 4077 23032
rect 3660 22992 3666 23004
rect 4065 23001 4077 23004
rect 4111 23001 4123 23035
rect 4065 22995 4123 23001
rect 4295 23035 4344 23041
rect 4295 23001 4307 23035
rect 4341 23001 4344 23035
rect 4295 22995 4344 23001
rect 4338 22992 4344 22995
rect 4396 23032 4402 23044
rect 4982 23032 4988 23044
rect 4396 23004 4988 23032
rect 4396 22992 4402 23004
rect 4982 22992 4988 23004
rect 5040 22992 5046 23044
rect 5074 22992 5080 23044
rect 5132 22992 5138 23044
rect 7006 23032 7012 23044
rect 6564 23004 7012 23032
rect 2317 22967 2375 22973
rect 2317 22933 2329 22967
rect 2363 22933 2375 22967
rect 2317 22927 2375 22933
rect 2774 22924 2780 22976
rect 2832 22924 2838 22976
rect 6564 22973 6592 23004
rect 7006 22992 7012 23004
rect 7064 22992 7070 23044
rect 6549 22967 6607 22973
rect 6549 22933 6561 22967
rect 6595 22933 6607 22967
rect 6549 22927 6607 22933
rect 6638 22924 6644 22976
rect 6696 22924 6702 22976
rect 6730 22924 6736 22976
rect 6788 22964 6794 22976
rect 7101 22967 7159 22973
rect 7101 22964 7113 22967
rect 6788 22936 7113 22964
rect 6788 22924 6794 22936
rect 7101 22933 7113 22936
rect 7147 22933 7159 22967
rect 8226 22964 8254 23063
rect 8478 23060 8484 23112
rect 8536 23109 8542 23112
rect 8536 23103 8565 23109
rect 8553 23069 8565 23103
rect 8536 23063 8565 23069
rect 8536 23060 8542 23063
rect 8662 23060 8668 23112
rect 8720 23060 8726 23112
rect 9416 23100 9444 23196
rect 10137 23171 10195 23177
rect 10137 23137 10149 23171
rect 10183 23168 10195 23171
rect 10226 23168 10232 23180
rect 10183 23140 10232 23168
rect 10183 23137 10195 23140
rect 10137 23131 10195 23137
rect 10226 23128 10232 23140
rect 10284 23128 10290 23180
rect 9585 23103 9643 23109
rect 9585 23100 9597 23103
rect 9416 23072 9597 23100
rect 9585 23069 9597 23072
rect 9631 23069 9643 23103
rect 9585 23063 9643 23069
rect 9677 23103 9735 23109
rect 9677 23069 9689 23103
rect 9723 23100 9735 23103
rect 9861 23103 9919 23109
rect 9861 23100 9873 23103
rect 9723 23072 9873 23100
rect 9723 23069 9735 23072
rect 9677 23063 9735 23069
rect 9861 23069 9873 23072
rect 9907 23069 9919 23103
rect 11348 23100 11376 23196
rect 13446 23168 13452 23180
rect 12912 23140 13452 23168
rect 12912 23112 12940 23140
rect 13446 23128 13452 23140
rect 13504 23168 13510 23180
rect 13740 23168 13768 23196
rect 14829 23171 14887 23177
rect 13504 23140 13584 23168
rect 13740 23140 14228 23168
rect 13504 23128 13510 23140
rect 11270 23072 11376 23100
rect 9861 23063 9919 23069
rect 12894 23060 12900 23112
rect 12952 23060 12958 23112
rect 13556 23109 13584 23140
rect 14200 23112 14228 23140
rect 14829 23137 14841 23171
rect 14875 23168 14887 23171
rect 15102 23168 15108 23180
rect 14875 23140 15108 23168
rect 14875 23137 14887 23140
rect 14829 23131 14887 23137
rect 15102 23128 15108 23140
rect 15160 23128 15166 23180
rect 15212 23168 15240 23208
rect 16022 23196 16028 23248
rect 16080 23196 16086 23248
rect 16298 23196 16304 23248
rect 16356 23196 16362 23248
rect 17586 23236 17592 23248
rect 16500 23208 17592 23236
rect 16500 23168 16528 23208
rect 17586 23196 17592 23208
rect 17644 23196 17650 23248
rect 15212 23140 16528 23168
rect 16666 23128 16672 23180
rect 16724 23168 16730 23180
rect 17034 23168 17040 23180
rect 16724 23140 17040 23168
rect 16724 23128 16730 23140
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 17696 23168 17724 23267
rect 18598 23264 18604 23276
rect 18656 23264 18662 23316
rect 20622 23264 20628 23316
rect 20680 23304 20686 23316
rect 21634 23304 21640 23316
rect 20680 23276 21640 23304
rect 20680 23264 20686 23276
rect 21634 23264 21640 23276
rect 21692 23264 21698 23316
rect 22922 23304 22928 23316
rect 21744 23276 22928 23304
rect 17770 23196 17776 23248
rect 17828 23236 17834 23248
rect 21358 23236 21364 23248
rect 17828 23208 21364 23236
rect 17828 23196 17834 23208
rect 21358 23196 21364 23208
rect 21416 23196 21422 23248
rect 17696 23140 18644 23168
rect 18616 23112 18644 23140
rect 18874 23128 18880 23180
rect 18932 23168 18938 23180
rect 19245 23171 19303 23177
rect 19245 23168 19257 23171
rect 18932 23140 19257 23168
rect 18932 23128 18938 23140
rect 19245 23137 19257 23140
rect 19291 23168 19303 23171
rect 21174 23168 21180 23180
rect 19291 23140 21180 23168
rect 19291 23137 19303 23140
rect 19245 23131 19303 23137
rect 21174 23128 21180 23140
rect 21232 23168 21238 23180
rect 21634 23168 21640 23180
rect 21232 23140 21640 23168
rect 21232 23128 21238 23140
rect 21634 23128 21640 23140
rect 21692 23128 21698 23180
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23069 13599 23103
rect 13541 23063 13599 23069
rect 8294 22992 8300 23044
rect 8352 22992 8358 23044
rect 8938 22992 8944 23044
rect 8996 22992 9002 23044
rect 9122 22992 9128 23044
rect 9180 22992 9186 23044
rect 11882 22992 11888 23044
rect 11940 23032 11946 23044
rect 13372 23032 13400 23063
rect 13722 23060 13728 23112
rect 13780 23100 13786 23112
rect 13909 23103 13967 23109
rect 13909 23100 13921 23103
rect 13780 23072 13921 23100
rect 13780 23060 13786 23072
rect 13909 23069 13921 23072
rect 13955 23100 13967 23103
rect 14093 23103 14151 23109
rect 14093 23100 14105 23103
rect 13955 23072 14105 23100
rect 13955 23069 13967 23072
rect 13909 23063 13967 23069
rect 14093 23069 14105 23072
rect 14139 23069 14151 23103
rect 14093 23063 14151 23069
rect 14182 23060 14188 23112
rect 14240 23060 14246 23112
rect 14921 23103 14979 23109
rect 14921 23069 14933 23103
rect 14967 23100 14979 23103
rect 14967 23072 15148 23100
rect 14967 23069 14979 23072
rect 14921 23063 14979 23069
rect 15120 23032 15148 23072
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 16206 23100 16212 23112
rect 15344 23072 16212 23100
rect 15344 23060 15350 23072
rect 16206 23060 16212 23072
rect 16264 23060 16270 23112
rect 16390 23060 16396 23112
rect 16448 23100 16454 23112
rect 16761 23103 16819 23109
rect 16761 23100 16773 23103
rect 16448 23072 16773 23100
rect 16448 23060 16454 23072
rect 16761 23069 16773 23072
rect 16807 23100 16819 23103
rect 17402 23100 17408 23112
rect 16807 23072 17408 23100
rect 16807 23069 16819 23072
rect 16761 23063 16819 23069
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 17957 23103 18015 23109
rect 17957 23100 17969 23103
rect 17512 23072 17969 23100
rect 17512 23044 17540 23072
rect 17957 23069 17969 23072
rect 18003 23100 18015 23103
rect 18506 23100 18512 23112
rect 18003 23072 18512 23100
rect 18003 23069 18015 23072
rect 17957 23063 18015 23069
rect 18506 23060 18512 23072
rect 18564 23060 18570 23112
rect 18598 23060 18604 23112
rect 18656 23060 18662 23112
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23100 18843 23103
rect 19058 23100 19064 23112
rect 18831 23072 19064 23100
rect 18831 23069 18843 23072
rect 18785 23063 18843 23069
rect 11940 23004 12434 23032
rect 13372 23004 15148 23032
rect 11940 22992 11946 23004
rect 9309 22967 9367 22973
rect 9309 22964 9321 22967
rect 8226 22936 9321 22964
rect 7101 22927 7159 22933
rect 9309 22933 9321 22936
rect 9355 22933 9367 22967
rect 12406 22964 12434 23004
rect 15120 22976 15148 23004
rect 16942 22992 16948 23044
rect 17000 22992 17006 23044
rect 17494 22992 17500 23044
rect 17552 22992 17558 23044
rect 17713 23035 17771 23041
rect 17713 23001 17725 23035
rect 17759 23032 17771 23035
rect 18800 23032 18828 23063
rect 19058 23060 19064 23072
rect 19116 23100 19122 23112
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 19116 23072 19533 23100
rect 19116 23060 19122 23072
rect 19521 23069 19533 23072
rect 19567 23069 19579 23103
rect 20714 23100 20720 23112
rect 19521 23063 19579 23069
rect 19904 23072 20720 23100
rect 19904 23044 19932 23072
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 17759 23004 18828 23032
rect 17759 23001 17771 23004
rect 17713 22995 17771 23001
rect 18966 22992 18972 23044
rect 19024 23032 19030 23044
rect 19613 23035 19671 23041
rect 19024 23004 19564 23032
rect 19024 22992 19030 23004
rect 15010 22964 15016 22976
rect 12406 22936 15016 22964
rect 9309 22927 9367 22933
rect 15010 22924 15016 22936
rect 15068 22924 15074 22976
rect 15102 22924 15108 22976
rect 15160 22924 15166 22976
rect 16960 22964 16988 22992
rect 18049 22967 18107 22973
rect 18049 22964 18061 22967
rect 16960 22936 18061 22964
rect 18049 22933 18061 22936
rect 18095 22933 18107 22967
rect 18049 22927 18107 22933
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 18874 22964 18880 22976
rect 18656 22936 18880 22964
rect 18656 22924 18662 22936
rect 18874 22924 18880 22936
rect 18932 22964 18938 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 18932 22936 19441 22964
rect 18932 22924 18938 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 19536 22964 19564 23004
rect 19613 23001 19625 23035
rect 19659 23032 19671 23035
rect 19886 23032 19892 23044
rect 19659 23004 19892 23032
rect 19659 23001 19671 23004
rect 19613 22995 19671 23001
rect 19886 22992 19892 23004
rect 19944 22992 19950 23044
rect 19981 23035 20039 23041
rect 19981 23001 19993 23035
rect 20027 23032 20039 23035
rect 20070 23032 20076 23044
rect 20027 23004 20076 23032
rect 20027 23001 20039 23004
rect 19981 22995 20039 23001
rect 20070 22992 20076 23004
rect 20128 23032 20134 23044
rect 20254 23032 20260 23044
rect 20128 23004 20260 23032
rect 20128 22992 20134 23004
rect 20254 22992 20260 23004
rect 20312 22992 20318 23044
rect 20530 22992 20536 23044
rect 20588 22992 20594 23044
rect 21652 23032 21680 23128
rect 21744 23109 21772 23276
rect 22922 23264 22928 23276
rect 22980 23264 22986 23316
rect 24578 23264 24584 23316
rect 24636 23304 24642 23316
rect 24673 23307 24731 23313
rect 24673 23304 24685 23307
rect 24636 23276 24685 23304
rect 24636 23264 24642 23276
rect 24673 23273 24685 23276
rect 24719 23273 24731 23307
rect 24673 23267 24731 23273
rect 27341 23307 27399 23313
rect 27341 23273 27353 23307
rect 27387 23304 27399 23307
rect 28810 23304 28816 23316
rect 27387 23276 28816 23304
rect 27387 23273 27399 23276
rect 27341 23267 27399 23273
rect 28810 23264 28816 23276
rect 28868 23264 28874 23316
rect 33870 23264 33876 23316
rect 33928 23304 33934 23316
rect 35618 23304 35624 23316
rect 33928 23276 35624 23304
rect 33928 23264 33934 23276
rect 35618 23264 35624 23276
rect 35676 23304 35682 23316
rect 35676 23276 36492 23304
rect 35676 23264 35682 23276
rect 25777 23239 25835 23245
rect 22388 23208 22876 23236
rect 22388 23180 22416 23208
rect 22186 23128 22192 23180
rect 22244 23168 22250 23180
rect 22244 23140 22325 23168
rect 22244 23128 22250 23140
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23069 21787 23103
rect 21729 23063 21787 23069
rect 21910 23060 21916 23112
rect 21968 23100 21974 23112
rect 21968 23096 22048 23100
rect 22094 23096 22100 23112
rect 21968 23072 22100 23096
rect 21968 23060 21974 23072
rect 22020 23068 22100 23072
rect 22094 23060 22100 23068
rect 22152 23060 22158 23112
rect 22297 23100 22325 23140
rect 22370 23128 22376 23180
rect 22428 23128 22434 23180
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23168 22523 23171
rect 22646 23168 22652 23180
rect 22511 23140 22652 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 22646 23128 22652 23140
rect 22704 23128 22710 23180
rect 22848 23177 22876 23208
rect 25777 23205 25789 23239
rect 25823 23236 25835 23239
rect 34238 23236 34244 23248
rect 25823 23208 34244 23236
rect 25823 23205 25835 23208
rect 25777 23199 25835 23205
rect 34238 23196 34244 23208
rect 34296 23196 34302 23248
rect 35268 23208 36308 23236
rect 22833 23171 22891 23177
rect 22833 23137 22845 23171
rect 22879 23137 22891 23171
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 22833 23131 22891 23137
rect 23124 23140 23489 23168
rect 23124 23112 23152 23140
rect 23477 23137 23489 23140
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 24486 23128 24492 23180
rect 24544 23168 24550 23180
rect 25314 23168 25320 23180
rect 24544 23140 25320 23168
rect 24544 23128 24550 23140
rect 25314 23128 25320 23140
rect 25372 23168 25378 23180
rect 26510 23168 26516 23180
rect 25372 23140 26516 23168
rect 25372 23128 25378 23140
rect 22554 23100 22560 23112
rect 22297 23072 22560 23100
rect 22554 23060 22560 23072
rect 22612 23060 22618 23112
rect 22738 23060 22744 23112
rect 22796 23100 22802 23112
rect 22925 23103 22983 23109
rect 22925 23100 22937 23103
rect 22796 23072 22937 23100
rect 22796 23060 22802 23072
rect 22925 23069 22937 23072
rect 22971 23069 22983 23103
rect 22925 23063 22983 23069
rect 23106 23060 23112 23112
rect 23164 23060 23170 23112
rect 23293 23103 23351 23109
rect 23293 23069 23305 23103
rect 23339 23069 23351 23103
rect 23293 23063 23351 23069
rect 21821 23035 21879 23041
rect 21821 23032 21833 23035
rect 21652 23004 21833 23032
rect 21821 23001 21833 23004
rect 21867 23001 21879 23035
rect 22112 23032 22140 23060
rect 23308 23032 23336 23063
rect 24854 23060 24860 23112
rect 24912 23060 24918 23112
rect 25222 23060 25228 23112
rect 25280 23060 25286 23112
rect 25424 23109 25452 23140
rect 26510 23128 26516 23140
rect 26568 23168 26574 23180
rect 27246 23168 27252 23180
rect 26568 23140 27252 23168
rect 26568 23128 26574 23140
rect 27246 23128 27252 23140
rect 27304 23128 27310 23180
rect 25409 23103 25467 23109
rect 25409 23069 25421 23103
rect 25455 23069 25467 23103
rect 25409 23063 25467 23069
rect 25590 23060 25596 23112
rect 25648 23109 25654 23112
rect 25648 23100 25656 23109
rect 25648 23072 25693 23100
rect 25648 23063 25656 23072
rect 25648 23060 25654 23063
rect 26602 23060 26608 23112
rect 26660 23100 26666 23112
rect 26660 23072 27200 23100
rect 26660 23060 26666 23072
rect 22112 23004 23336 23032
rect 21821 22995 21879 23001
rect 25498 22992 25504 23044
rect 25556 22992 25562 23044
rect 27062 22992 27068 23044
rect 27120 22992 27126 23044
rect 27172 23032 27200 23072
rect 31202 23060 31208 23112
rect 31260 23100 31266 23112
rect 31747 23103 31805 23109
rect 31260 23096 31616 23100
rect 31747 23096 31759 23103
rect 31260 23072 31759 23096
rect 31260 23060 31266 23072
rect 31588 23069 31759 23072
rect 31793 23069 31805 23103
rect 31588 23068 31805 23069
rect 31747 23063 31805 23068
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23100 31999 23103
rect 32122 23100 32128 23112
rect 31987 23072 32128 23100
rect 31987 23069 31999 23072
rect 31941 23063 31999 23069
rect 32122 23060 32128 23072
rect 32180 23060 32186 23112
rect 33962 23060 33968 23112
rect 34020 23100 34026 23112
rect 35268 23109 35296 23208
rect 36081 23171 36139 23177
rect 36081 23168 36093 23171
rect 35452 23140 36093 23168
rect 35452 23109 35480 23140
rect 36081 23137 36093 23140
rect 36127 23137 36139 23171
rect 36081 23131 36139 23137
rect 35253 23103 35311 23109
rect 35253 23100 35265 23103
rect 34020 23072 35265 23100
rect 34020 23060 34026 23072
rect 35253 23069 35265 23072
rect 35299 23069 35311 23103
rect 35253 23063 35311 23069
rect 35437 23103 35495 23109
rect 35437 23069 35449 23103
rect 35483 23069 35495 23103
rect 35437 23063 35495 23069
rect 35268 23032 35296 23063
rect 35618 23060 35624 23112
rect 35676 23100 35682 23112
rect 36280 23109 36308 23208
rect 36464 23109 36492 23276
rect 35713 23103 35771 23109
rect 35713 23100 35725 23103
rect 35676 23072 35725 23100
rect 35676 23060 35682 23072
rect 35713 23069 35725 23072
rect 35759 23100 35771 23103
rect 35989 23103 36047 23109
rect 35989 23100 36001 23103
rect 35759 23072 36001 23100
rect 35759 23069 35771 23072
rect 35713 23063 35771 23069
rect 35989 23069 36001 23072
rect 36035 23069 36047 23103
rect 35989 23063 36047 23069
rect 36265 23103 36323 23109
rect 36265 23069 36277 23103
rect 36311 23069 36323 23103
rect 36265 23063 36323 23069
rect 36449 23103 36507 23109
rect 36449 23069 36461 23103
rect 36495 23069 36507 23103
rect 36449 23063 36507 23069
rect 37274 23060 37280 23112
rect 37332 23100 37338 23112
rect 37553 23103 37611 23109
rect 37553 23100 37565 23103
rect 37332 23072 37565 23100
rect 37332 23060 37338 23072
rect 37553 23069 37565 23072
rect 37599 23069 37611 23103
rect 37553 23063 37611 23069
rect 35529 23035 35587 23041
rect 35529 23032 35541 23035
rect 27172 23004 33640 23032
rect 35268 23004 35541 23032
rect 20548 22964 20576 22992
rect 33612 22976 33640 23004
rect 35529 23001 35541 23004
rect 35575 23001 35587 23035
rect 35529 22995 35587 23001
rect 35802 22992 35808 23044
rect 35860 23032 35866 23044
rect 36357 23035 36415 23041
rect 36357 23032 36369 23035
rect 35860 23004 36369 23032
rect 35860 22992 35866 23004
rect 36357 23001 36369 23004
rect 36403 23001 36415 23035
rect 36357 22995 36415 23001
rect 19536 22936 20576 22964
rect 19429 22927 19487 22933
rect 20990 22924 20996 22976
rect 21048 22964 21054 22976
rect 21453 22967 21511 22973
rect 21453 22964 21465 22967
rect 21048 22936 21465 22964
rect 21048 22924 21054 22936
rect 21453 22933 21465 22936
rect 21499 22933 21511 22967
rect 21453 22927 21511 22933
rect 21913 22967 21971 22973
rect 21913 22933 21925 22967
rect 21959 22964 21971 22967
rect 22094 22964 22100 22976
rect 21959 22936 22100 22964
rect 21959 22933 21971 22936
rect 21913 22927 21971 22933
rect 22094 22924 22100 22936
rect 22152 22964 22158 22976
rect 22370 22964 22376 22976
rect 22152 22936 22376 22964
rect 22152 22924 22158 22936
rect 22370 22924 22376 22936
rect 22428 22924 22434 22976
rect 22554 22924 22560 22976
rect 22612 22964 22618 22976
rect 23658 22964 23664 22976
rect 22612 22936 23664 22964
rect 22612 22924 22618 22936
rect 23658 22924 23664 22936
rect 23716 22924 23722 22976
rect 24394 22924 24400 22976
rect 24452 22964 24458 22976
rect 30926 22964 30932 22976
rect 24452 22936 30932 22964
rect 24452 22924 24458 22936
rect 30926 22924 30932 22936
rect 30984 22924 30990 22976
rect 31941 22967 31999 22973
rect 31941 22933 31953 22967
rect 31987 22964 31999 22967
rect 32306 22964 32312 22976
rect 31987 22936 32312 22964
rect 31987 22933 31999 22936
rect 31941 22927 31999 22933
rect 32306 22924 32312 22936
rect 32364 22924 32370 22976
rect 33594 22924 33600 22976
rect 33652 22924 33658 22976
rect 35342 22924 35348 22976
rect 35400 22924 35406 22976
rect 35894 22924 35900 22976
rect 35952 22924 35958 22976
rect 37366 22924 37372 22976
rect 37424 22924 37430 22976
rect 1104 22874 38272 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38272 22874
rect 1104 22800 38272 22822
rect 1486 22720 1492 22772
rect 1544 22760 1550 22772
rect 2133 22763 2191 22769
rect 2133 22760 2145 22763
rect 1544 22732 2145 22760
rect 1544 22720 1550 22732
rect 2133 22729 2145 22732
rect 2179 22729 2191 22763
rect 2682 22760 2688 22772
rect 2133 22723 2191 22729
rect 2424 22732 2688 22760
rect 2424 22633 2452 22732
rect 2682 22720 2688 22732
rect 2740 22720 2746 22772
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 3329 22763 3387 22769
rect 3329 22760 3341 22763
rect 2832 22732 3341 22760
rect 2832 22720 2838 22732
rect 3329 22729 3341 22732
rect 3375 22729 3387 22763
rect 3329 22723 3387 22729
rect 3602 22720 3608 22772
rect 3660 22720 3666 22772
rect 3970 22720 3976 22772
rect 4028 22760 4034 22772
rect 4433 22763 4491 22769
rect 4433 22760 4445 22763
rect 4028 22732 4445 22760
rect 4028 22720 4034 22732
rect 4433 22729 4445 22732
rect 4479 22729 4491 22763
rect 4433 22723 4491 22729
rect 5074 22720 5080 22772
rect 5132 22760 5138 22772
rect 5353 22763 5411 22769
rect 5353 22760 5365 22763
rect 5132 22732 5365 22760
rect 5132 22720 5138 22732
rect 5353 22729 5365 22732
rect 5399 22729 5411 22763
rect 6638 22760 6644 22772
rect 5353 22723 5411 22729
rect 5552 22732 6644 22760
rect 2700 22692 2728 22720
rect 3145 22695 3203 22701
rect 2700 22664 3004 22692
rect 2409 22627 2467 22633
rect 2409 22593 2421 22627
rect 2455 22593 2467 22627
rect 2409 22587 2467 22593
rect 2498 22584 2504 22636
rect 2556 22584 2562 22636
rect 2590 22584 2596 22636
rect 2648 22584 2654 22636
rect 2774 22584 2780 22636
rect 2832 22584 2838 22636
rect 2976 22556 3004 22664
rect 3145 22661 3157 22695
rect 3191 22692 3203 22695
rect 3620 22692 3648 22720
rect 3191 22664 3648 22692
rect 3191 22661 3203 22664
rect 3145 22655 3203 22661
rect 3694 22652 3700 22704
rect 3752 22692 3758 22704
rect 4154 22692 4160 22704
rect 3752 22664 4160 22692
rect 3752 22652 3758 22664
rect 4154 22652 4160 22664
rect 4212 22652 4218 22704
rect 4246 22652 4252 22704
rect 4304 22692 4310 22704
rect 4525 22695 4583 22701
rect 4525 22692 4537 22695
rect 4304 22664 4537 22692
rect 4304 22652 4310 22664
rect 4525 22661 4537 22664
rect 4571 22661 4583 22695
rect 4525 22655 4583 22661
rect 4755 22661 4813 22667
rect 4755 22658 4767 22661
rect 3050 22584 3056 22636
rect 3108 22584 3114 22636
rect 3237 22627 3295 22633
rect 3237 22593 3249 22627
rect 3283 22593 3295 22627
rect 3237 22587 3295 22593
rect 3252 22556 3280 22587
rect 3510 22584 3516 22636
rect 3568 22584 3574 22636
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22593 3663 22627
rect 3835 22627 3893 22633
rect 3835 22624 3847 22627
rect 3605 22587 3663 22593
rect 3830 22593 3847 22624
rect 3881 22593 3893 22627
rect 3830 22587 3893 22593
rect 2976 22528 3280 22556
rect 3252 22432 3280 22528
rect 3620 22488 3648 22587
rect 3830 22556 3858 22587
rect 3970 22584 3976 22636
rect 4028 22584 4034 22636
rect 4062 22584 4068 22636
rect 4120 22624 4126 22636
rect 4614 22624 4620 22636
rect 4120 22596 4620 22624
rect 4120 22584 4126 22596
rect 4614 22584 4620 22596
rect 4672 22624 4678 22636
rect 4740 22627 4767 22658
rect 4801 22627 4813 22661
rect 5552 22633 5580 22732
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 7190 22720 7196 22772
rect 7248 22720 7254 22772
rect 7650 22760 7656 22772
rect 7300 22732 7656 22760
rect 7009 22695 7067 22701
rect 7009 22661 7021 22695
rect 7055 22692 7067 22695
rect 7208 22692 7236 22720
rect 7055 22664 7236 22692
rect 7055 22661 7067 22664
rect 7009 22655 7067 22661
rect 4740 22624 4813 22627
rect 4672 22621 4813 22624
rect 4985 22627 5043 22633
rect 4672 22596 4768 22621
rect 4672 22584 4678 22596
rect 4985 22593 4997 22627
rect 5031 22624 5043 22627
rect 5537 22627 5595 22633
rect 5031 22596 5212 22624
rect 5031 22593 5043 22596
rect 4985 22587 5043 22593
rect 4338 22556 4344 22568
rect 3830 22528 4344 22556
rect 4338 22516 4344 22528
rect 4396 22516 4402 22568
rect 5077 22491 5135 22497
rect 5077 22488 5089 22491
rect 3620 22460 5089 22488
rect 5077 22457 5089 22460
rect 5123 22457 5135 22491
rect 5077 22451 5135 22457
rect 3234 22380 3240 22432
rect 3292 22420 3298 22432
rect 4246 22420 4252 22432
rect 3292 22392 4252 22420
rect 3292 22380 3298 22392
rect 4246 22380 4252 22392
rect 4304 22380 4310 22432
rect 4709 22423 4767 22429
rect 4709 22389 4721 22423
rect 4755 22420 4767 22423
rect 4798 22420 4804 22432
rect 4755 22392 4804 22420
rect 4755 22389 4767 22392
rect 4709 22383 4767 22389
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 4893 22423 4951 22429
rect 4893 22389 4905 22423
rect 4939 22420 4951 22423
rect 5184 22420 5212 22596
rect 5537 22593 5549 22627
rect 5583 22593 5595 22627
rect 5537 22587 5595 22593
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 6730 22624 6736 22636
rect 6687 22596 6736 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 6825 22627 6883 22633
rect 6825 22593 6837 22627
rect 6871 22593 6883 22627
rect 6825 22587 6883 22593
rect 6840 22556 6868 22587
rect 6914 22584 6920 22636
rect 6972 22584 6978 22636
rect 7098 22584 7104 22636
rect 7156 22633 7162 22636
rect 7156 22627 7185 22633
rect 7173 22593 7185 22627
rect 7156 22587 7185 22593
rect 7156 22584 7162 22587
rect 7300 22565 7328 22732
rect 7650 22720 7656 22732
rect 7708 22760 7714 22772
rect 7708 22732 8156 22760
rect 7708 22720 7714 22732
rect 8128 22704 8156 22732
rect 8294 22720 8300 22772
rect 8352 22720 8358 22772
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10045 22763 10103 22769
rect 10045 22760 10057 22763
rect 9916 22732 10057 22760
rect 9916 22720 9922 22732
rect 10045 22729 10057 22732
rect 10091 22729 10103 22763
rect 10045 22723 10103 22729
rect 11514 22720 11520 22772
rect 11572 22720 11578 22772
rect 11882 22720 11888 22772
rect 11940 22720 11946 22772
rect 11974 22720 11980 22772
rect 12032 22760 12038 22772
rect 15010 22760 15016 22772
rect 12032 22732 12434 22760
rect 12032 22720 12038 22732
rect 7374 22652 7380 22704
rect 7432 22692 7438 22704
rect 7432 22664 7880 22692
rect 7432 22652 7438 22664
rect 7466 22584 7472 22636
rect 7524 22627 7530 22636
rect 7852 22633 7880 22664
rect 8110 22652 8116 22704
rect 8168 22652 8174 22704
rect 8938 22692 8944 22704
rect 8226 22664 8944 22692
rect 8226 22633 8254 22664
rect 8938 22652 8944 22664
rect 8996 22652 9002 22704
rect 10505 22695 10563 22701
rect 10505 22661 10517 22695
rect 10551 22692 10563 22695
rect 10962 22692 10968 22704
rect 10551 22664 10968 22692
rect 10551 22661 10563 22664
rect 10505 22655 10563 22661
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 7580 22627 7638 22633
rect 7524 22599 7592 22627
rect 7524 22584 7530 22599
rect 7576 22596 7592 22599
rect 7580 22593 7592 22596
rect 7626 22593 7638 22627
rect 7745 22627 7803 22633
rect 7745 22624 7757 22627
rect 7580 22587 7638 22593
rect 7668 22596 7757 22624
rect 7285 22559 7343 22565
rect 6840 22528 6960 22556
rect 6932 22488 6960 22528
rect 7285 22525 7297 22559
rect 7331 22525 7343 22559
rect 7285 22519 7343 22525
rect 7377 22491 7435 22497
rect 7377 22488 7389 22491
rect 6932 22460 7389 22488
rect 7377 22457 7389 22460
rect 7423 22457 7435 22491
rect 7377 22451 7435 22457
rect 7190 22420 7196 22432
rect 4939 22392 7196 22420
rect 4939 22389 4951 22392
rect 4893 22383 4951 22389
rect 7190 22380 7196 22392
rect 7248 22380 7254 22432
rect 7282 22380 7288 22432
rect 7340 22420 7346 22432
rect 7558 22420 7564 22432
rect 7340 22392 7564 22420
rect 7340 22380 7346 22392
rect 7558 22380 7564 22392
rect 7616 22420 7622 22432
rect 7668 22420 7696 22596
rect 7745 22593 7757 22596
rect 7791 22593 7803 22627
rect 7745 22587 7803 22593
rect 7837 22627 7895 22633
rect 7837 22593 7849 22627
rect 7883 22624 7895 22627
rect 8205 22627 8263 22633
rect 8205 22624 8217 22627
rect 7883 22596 8217 22624
rect 7883 22593 7895 22596
rect 7837 22587 7895 22593
rect 8205 22593 8217 22596
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22593 8447 22627
rect 8389 22587 8447 22593
rect 10413 22627 10471 22633
rect 10413 22593 10425 22627
rect 10459 22624 10471 22627
rect 11992 22624 12020 22720
rect 10459 22596 12020 22624
rect 12406 22636 12434 22732
rect 14016 22732 15016 22760
rect 14016 22701 14044 22732
rect 15010 22720 15016 22732
rect 15068 22720 15074 22772
rect 21082 22760 21088 22772
rect 15212 22732 21088 22760
rect 14001 22695 14059 22701
rect 14001 22661 14013 22695
rect 14047 22661 14059 22695
rect 15212 22692 15240 22732
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 21269 22763 21327 22769
rect 21269 22729 21281 22763
rect 21315 22760 21327 22763
rect 21450 22760 21456 22772
rect 21315 22732 21456 22760
rect 21315 22729 21327 22732
rect 21269 22723 21327 22729
rect 21450 22720 21456 22732
rect 21508 22760 21514 22772
rect 21910 22760 21916 22772
rect 21508 22732 21916 22760
rect 21508 22720 21514 22732
rect 21910 22720 21916 22732
rect 21968 22760 21974 22772
rect 22189 22763 22247 22769
rect 21968 22732 22140 22760
rect 21968 22720 21974 22732
rect 14001 22655 14059 22661
rect 14936 22664 15240 22692
rect 12406 22596 12440 22636
rect 10459 22593 10471 22596
rect 10413 22587 10471 22593
rect 8404 22432 8432 22587
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 14274 22584 14280 22636
rect 14332 22624 14338 22636
rect 14734 22624 14740 22636
rect 14332 22596 14740 22624
rect 14332 22584 14338 22596
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 10689 22559 10747 22565
rect 10689 22525 10701 22559
rect 10735 22556 10747 22559
rect 10778 22556 10784 22568
rect 10735 22528 10784 22556
rect 10735 22525 10747 22528
rect 10689 22519 10747 22525
rect 10778 22516 10784 22528
rect 10836 22516 10842 22568
rect 11974 22516 11980 22568
rect 12032 22516 12038 22568
rect 12158 22516 12164 22568
rect 12216 22516 12222 22568
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22525 14151 22559
rect 14936 22556 14964 22664
rect 15746 22652 15752 22704
rect 15804 22692 15810 22704
rect 16209 22695 16267 22701
rect 16209 22692 16221 22695
rect 15804 22664 16221 22692
rect 15804 22652 15810 22664
rect 16209 22661 16221 22664
rect 16255 22661 16267 22695
rect 18138 22692 18144 22704
rect 16209 22655 16267 22661
rect 16316 22664 18144 22692
rect 15010 22584 15016 22636
rect 15068 22584 15074 22636
rect 15197 22627 15255 22633
rect 15197 22593 15209 22627
rect 15243 22624 15255 22627
rect 15378 22624 15384 22636
rect 15243 22596 15384 22624
rect 15243 22593 15255 22596
rect 15197 22587 15255 22593
rect 15378 22584 15384 22596
rect 15436 22584 15442 22636
rect 15470 22584 15476 22636
rect 15528 22584 15534 22636
rect 15838 22584 15844 22636
rect 15896 22624 15902 22636
rect 16316 22624 16344 22664
rect 18138 22652 18144 22664
rect 18196 22652 18202 22704
rect 21818 22692 21824 22704
rect 18248 22664 21824 22692
rect 15896 22596 16344 22624
rect 15896 22584 15902 22596
rect 17310 22584 17316 22636
rect 17368 22584 17374 22636
rect 17678 22584 17684 22636
rect 17736 22584 17742 22636
rect 14093 22519 14151 22525
rect 14200 22528 14964 22556
rect 11422 22448 11428 22500
rect 11480 22488 11486 22500
rect 13170 22488 13176 22500
rect 11480 22460 13176 22488
rect 11480 22448 11486 22460
rect 13170 22448 13176 22460
rect 13228 22488 13234 22500
rect 13722 22488 13728 22500
rect 13228 22460 13728 22488
rect 13228 22448 13234 22460
rect 13722 22448 13728 22460
rect 13780 22488 13786 22500
rect 14108 22488 14136 22519
rect 13780 22460 14136 22488
rect 13780 22448 13786 22460
rect 8386 22420 8392 22432
rect 7616 22392 8392 22420
rect 7616 22380 7622 22392
rect 8386 22380 8392 22392
rect 8444 22380 8450 22432
rect 8478 22380 8484 22432
rect 8536 22420 8542 22432
rect 8662 22420 8668 22432
rect 8536 22392 8668 22420
rect 8536 22380 8542 22392
rect 8662 22380 8668 22392
rect 8720 22420 8726 22432
rect 14200 22420 14228 22528
rect 14461 22491 14519 22497
rect 14461 22457 14473 22491
rect 14507 22457 14519 22491
rect 14461 22451 14519 22457
rect 8720 22392 14228 22420
rect 8720 22380 8726 22392
rect 14274 22380 14280 22432
rect 14332 22380 14338 22432
rect 14476 22420 14504 22451
rect 15194 22448 15200 22500
rect 15252 22448 15258 22500
rect 15396 22488 15424 22584
rect 16850 22516 16856 22568
rect 16908 22516 16914 22568
rect 17126 22516 17132 22568
rect 17184 22516 17190 22568
rect 17586 22556 17592 22568
rect 17236 22528 17592 22556
rect 16482 22488 16488 22500
rect 15396 22460 16488 22488
rect 16482 22448 16488 22460
rect 16540 22488 16546 22500
rect 17236 22488 17264 22528
rect 17586 22516 17592 22528
rect 17644 22516 17650 22568
rect 16540 22460 17264 22488
rect 16540 22448 16546 22460
rect 18248 22420 18276 22664
rect 21818 22652 21824 22664
rect 21876 22652 21882 22704
rect 22112 22692 22140 22732
rect 22189 22729 22201 22763
rect 22235 22760 22247 22763
rect 22738 22760 22744 22772
rect 22235 22732 22744 22760
rect 22235 22729 22247 22732
rect 22189 22723 22247 22729
rect 22738 22720 22744 22732
rect 22796 22720 22802 22772
rect 27246 22720 27252 22772
rect 27304 22720 27310 22772
rect 31202 22720 31208 22772
rect 31260 22720 31266 22772
rect 31404 22732 32260 22760
rect 22281 22695 22339 22701
rect 22281 22692 22293 22695
rect 22112 22664 22293 22692
rect 22281 22661 22293 22664
rect 22327 22661 22339 22695
rect 22281 22655 22339 22661
rect 27157 22695 27215 22701
rect 27157 22661 27169 22695
rect 27203 22692 27215 22695
rect 27264 22692 27292 22720
rect 28813 22695 28871 22701
rect 27203 22664 27292 22692
rect 27632 22664 28764 22692
rect 27203 22661 27215 22664
rect 27157 22655 27215 22661
rect 27632 22636 27660 22664
rect 28736 22636 28764 22664
rect 28813 22661 28825 22695
rect 28859 22692 28871 22695
rect 28859 22664 29316 22692
rect 28859 22661 28871 22664
rect 28813 22655 28871 22661
rect 18322 22584 18328 22636
rect 18380 22584 18386 22636
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18417 22587 18475 22593
rect 18340 22497 18368 22584
rect 18432 22556 18460 22587
rect 18966 22584 18972 22636
rect 19024 22584 19030 22636
rect 19058 22584 19064 22636
rect 19116 22584 19122 22636
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 20438 22584 20444 22636
rect 20496 22584 20502 22636
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22624 20591 22627
rect 20622 22624 20628 22636
rect 20579 22596 20628 22624
rect 20579 22593 20591 22596
rect 20533 22587 20591 22593
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22593 20775 22627
rect 20717 22587 20775 22593
rect 18874 22556 18880 22568
rect 18432 22528 18880 22556
rect 18874 22516 18880 22528
rect 18932 22556 18938 22568
rect 19260 22556 19288 22584
rect 18932 22528 19288 22556
rect 18932 22516 18938 22528
rect 18325 22491 18383 22497
rect 18325 22457 18337 22491
rect 18371 22457 18383 22491
rect 18325 22451 18383 22457
rect 20257 22491 20315 22497
rect 20257 22457 20269 22491
rect 20303 22488 20315 22491
rect 20530 22488 20536 22500
rect 20303 22460 20536 22488
rect 20303 22457 20315 22460
rect 20257 22451 20315 22457
rect 20530 22448 20536 22460
rect 20588 22448 20594 22500
rect 20732 22488 20760 22587
rect 20898 22584 20904 22636
rect 20956 22624 20962 22636
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20956 22596 21097 22624
rect 20956 22584 20962 22596
rect 21085 22593 21097 22596
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21100 22556 21128 22587
rect 21174 22584 21180 22636
rect 21232 22584 21238 22636
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22624 22155 22627
rect 22462 22624 22468 22636
rect 22143 22596 22468 22624
rect 22143 22593 22155 22596
rect 22097 22587 22155 22593
rect 22462 22584 22468 22596
rect 22520 22584 22526 22636
rect 25590 22584 25596 22636
rect 25648 22584 25654 22636
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 26970 22624 26976 22636
rect 26384 22596 26976 22624
rect 26384 22584 26390 22596
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 27246 22584 27252 22636
rect 27304 22584 27310 22636
rect 27338 22584 27344 22636
rect 27396 22584 27402 22636
rect 27614 22584 27620 22636
rect 27672 22584 27678 22636
rect 27706 22584 27712 22636
rect 27764 22584 27770 22636
rect 28718 22584 28724 22636
rect 28776 22584 28782 22636
rect 29288 22633 29316 22664
rect 28905 22627 28963 22633
rect 28905 22593 28917 22627
rect 28951 22624 28963 22627
rect 28997 22627 29055 22633
rect 28997 22624 29009 22627
rect 28951 22596 29009 22624
rect 28951 22593 28963 22596
rect 28905 22587 28963 22593
rect 28997 22593 29009 22596
rect 29043 22593 29055 22627
rect 28997 22587 29055 22593
rect 29273 22627 29331 22633
rect 29273 22593 29285 22627
rect 29319 22593 29331 22627
rect 29273 22587 29331 22593
rect 21100 22528 21312 22556
rect 21174 22488 21180 22500
rect 20732 22460 21180 22488
rect 21174 22448 21180 22460
rect 21232 22448 21238 22500
rect 21284 22488 21312 22528
rect 21450 22516 21456 22568
rect 21508 22556 21514 22568
rect 21545 22559 21603 22565
rect 21545 22556 21557 22559
rect 21508 22528 21557 22556
rect 21508 22516 21514 22528
rect 21545 22525 21557 22528
rect 21591 22525 21603 22559
rect 21545 22519 21603 22525
rect 22370 22516 22376 22568
rect 22428 22556 22434 22568
rect 22557 22559 22615 22565
rect 22557 22556 22569 22559
rect 22428 22528 22569 22556
rect 22428 22516 22434 22528
rect 22557 22525 22569 22528
rect 22603 22556 22615 22559
rect 23106 22556 23112 22568
rect 22603 22528 23112 22556
rect 22603 22525 22615 22528
rect 22557 22519 22615 22525
rect 23106 22516 23112 22528
rect 23164 22516 23170 22568
rect 25608 22556 25636 22584
rect 27356 22556 27384 22584
rect 25608 22528 27384 22556
rect 27724 22556 27752 22584
rect 28810 22556 28816 22568
rect 27724 22528 28816 22556
rect 28810 22516 28816 22528
rect 28868 22556 28874 22568
rect 28920 22556 28948 22587
rect 29454 22584 29460 22636
rect 29512 22584 29518 22636
rect 31220 22633 31248 22720
rect 31404 22633 31432 22732
rect 32122 22692 32128 22704
rect 31956 22664 32128 22692
rect 31956 22633 31984 22664
rect 32122 22652 32128 22664
rect 32180 22652 32186 22704
rect 31205 22627 31263 22633
rect 31205 22593 31217 22627
rect 31251 22593 31263 22627
rect 31389 22627 31447 22633
rect 31389 22624 31401 22627
rect 31205 22587 31263 22593
rect 31312 22596 31401 22624
rect 28868 22528 28948 22556
rect 28868 22516 28874 22528
rect 30006 22516 30012 22568
rect 30064 22556 30070 22568
rect 31312 22556 31340 22596
rect 31389 22593 31401 22596
rect 31435 22593 31447 22627
rect 31389 22587 31447 22593
rect 31665 22627 31723 22633
rect 31665 22593 31677 22627
rect 31711 22593 31723 22627
rect 31665 22587 31723 22593
rect 31849 22627 31907 22633
rect 31849 22593 31861 22627
rect 31895 22593 31907 22627
rect 31849 22587 31907 22593
rect 31941 22627 31999 22633
rect 31941 22593 31953 22627
rect 31987 22593 31999 22627
rect 31941 22587 31999 22593
rect 30064 22528 31340 22556
rect 30064 22516 30070 22528
rect 22738 22488 22744 22500
rect 21284 22460 22744 22488
rect 22738 22448 22744 22460
rect 22796 22448 22802 22500
rect 31018 22488 31024 22500
rect 27540 22460 31024 22488
rect 14476 22392 18276 22420
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19981 22423 20039 22429
rect 19981 22420 19993 22423
rect 19392 22392 19993 22420
rect 19392 22380 19398 22392
rect 19981 22389 19993 22392
rect 20027 22389 20039 22423
rect 19981 22383 20039 22389
rect 20346 22380 20352 22432
rect 20404 22380 20410 22432
rect 20806 22380 20812 22432
rect 20864 22380 20870 22432
rect 21358 22380 21364 22432
rect 21416 22420 21422 22432
rect 21453 22423 21511 22429
rect 21453 22420 21465 22423
rect 21416 22392 21465 22420
rect 21416 22380 21422 22392
rect 21453 22389 21465 22392
rect 21499 22420 21511 22423
rect 21726 22420 21732 22432
rect 21499 22392 21732 22420
rect 21499 22389 21511 22392
rect 21453 22383 21511 22389
rect 21726 22380 21732 22392
rect 21784 22380 21790 22432
rect 21818 22380 21824 22432
rect 21876 22380 21882 22432
rect 22278 22380 22284 22432
rect 22336 22420 22342 22432
rect 27540 22429 27568 22460
rect 31018 22448 31024 22460
rect 31076 22448 31082 22500
rect 31297 22491 31355 22497
rect 31297 22457 31309 22491
rect 31343 22488 31355 22491
rect 31680 22488 31708 22587
rect 31754 22516 31760 22568
rect 31812 22556 31818 22568
rect 31864 22556 31892 22587
rect 31812 22528 31892 22556
rect 32232 22556 32260 22732
rect 32306 22720 32312 22772
rect 32364 22720 32370 22772
rect 34609 22763 34667 22769
rect 34609 22760 34621 22763
rect 34348 22732 34621 22760
rect 32324 22692 32352 22720
rect 32324 22664 32444 22692
rect 32416 22636 32444 22664
rect 32600 22664 32996 22692
rect 32306 22584 32312 22636
rect 32364 22584 32370 22636
rect 32398 22584 32404 22636
rect 32456 22584 32462 22636
rect 32600 22633 32628 22664
rect 32968 22636 32996 22664
rect 32585 22627 32643 22633
rect 32585 22593 32597 22627
rect 32631 22593 32643 22627
rect 32585 22587 32643 22593
rect 32677 22627 32735 22633
rect 32677 22593 32689 22627
rect 32723 22593 32735 22627
rect 32677 22587 32735 22593
rect 32692 22556 32720 22587
rect 32950 22584 32956 22636
rect 33008 22584 33014 22636
rect 34146 22584 34152 22636
rect 34204 22584 34210 22636
rect 34348 22633 34376 22732
rect 34609 22729 34621 22732
rect 34655 22760 34667 22763
rect 34698 22760 34704 22772
rect 34655 22732 34704 22760
rect 34655 22729 34667 22732
rect 34609 22723 34667 22729
rect 34698 22720 34704 22732
rect 34756 22720 34762 22772
rect 35894 22720 35900 22772
rect 35952 22720 35958 22772
rect 37366 22720 37372 22772
rect 37424 22720 37430 22772
rect 34425 22695 34483 22701
rect 34425 22661 34437 22695
rect 34471 22692 34483 22695
rect 34790 22692 34796 22704
rect 34471 22664 34796 22692
rect 34471 22661 34483 22664
rect 34425 22655 34483 22661
rect 34790 22652 34796 22664
rect 34848 22652 34854 22704
rect 35802 22692 35808 22704
rect 35636 22664 35808 22692
rect 34333 22627 34391 22633
rect 34333 22593 34345 22627
rect 34379 22593 34391 22627
rect 34333 22587 34391 22593
rect 34698 22584 34704 22636
rect 34756 22584 34762 22636
rect 35636 22633 35664 22664
rect 35802 22652 35808 22664
rect 35860 22652 35866 22704
rect 35621 22627 35679 22633
rect 35621 22593 35633 22627
rect 35667 22593 35679 22627
rect 35621 22587 35679 22593
rect 35713 22627 35771 22633
rect 35713 22593 35725 22627
rect 35759 22624 35771 22627
rect 35912 22624 35940 22720
rect 35759 22596 35940 22624
rect 37384 22624 37412 22720
rect 37645 22627 37703 22633
rect 37645 22624 37657 22627
rect 37384 22596 37657 22624
rect 35759 22593 35771 22596
rect 35713 22587 35771 22593
rect 37645 22593 37657 22596
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 32232 22528 32720 22556
rect 31812 22516 31818 22528
rect 31343 22460 31708 22488
rect 31864 22488 31892 22528
rect 33502 22488 33508 22500
rect 31864 22460 33508 22488
rect 31343 22457 31355 22460
rect 31297 22451 31355 22457
rect 33502 22448 33508 22460
rect 33560 22488 33566 22500
rect 33560 22460 34468 22488
rect 33560 22448 33566 22460
rect 22465 22423 22523 22429
rect 22465 22420 22477 22423
rect 22336 22392 22477 22420
rect 22336 22380 22342 22392
rect 22465 22389 22477 22392
rect 22511 22389 22523 22423
rect 22465 22383 22523 22389
rect 27525 22423 27583 22429
rect 27525 22389 27537 22423
rect 27571 22389 27583 22423
rect 27525 22383 27583 22389
rect 29086 22380 29092 22432
rect 29144 22380 29150 22432
rect 29273 22423 29331 22429
rect 29273 22389 29285 22423
rect 29319 22420 29331 22423
rect 29730 22420 29736 22432
rect 29319 22392 29736 22420
rect 29319 22389 29331 22392
rect 29273 22383 29331 22389
rect 29730 22380 29736 22392
rect 29788 22380 29794 22432
rect 31478 22380 31484 22432
rect 31536 22380 31542 22432
rect 32122 22380 32128 22432
rect 32180 22380 32186 22432
rect 34238 22380 34244 22432
rect 34296 22380 34302 22432
rect 34440 22429 34468 22460
rect 37826 22448 37832 22500
rect 37884 22448 37890 22500
rect 34425 22423 34483 22429
rect 34425 22389 34437 22423
rect 34471 22389 34483 22423
rect 34425 22383 34483 22389
rect 35894 22380 35900 22432
rect 35952 22380 35958 22432
rect 1104 22330 38272 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38272 22330
rect 1104 22256 38272 22278
rect 3510 22176 3516 22228
rect 3568 22216 3574 22228
rect 3789 22219 3847 22225
rect 3789 22216 3801 22219
rect 3568 22188 3801 22216
rect 3568 22176 3574 22188
rect 3789 22185 3801 22188
rect 3835 22185 3847 22219
rect 3789 22179 3847 22185
rect 6914 22176 6920 22228
rect 6972 22176 6978 22228
rect 7006 22176 7012 22228
rect 7064 22216 7070 22228
rect 7193 22219 7251 22225
rect 7193 22216 7205 22219
rect 7064 22188 7205 22216
rect 7064 22176 7070 22188
rect 7193 22185 7205 22188
rect 7239 22216 7251 22219
rect 7466 22216 7472 22228
rect 7239 22188 7472 22216
rect 7239 22185 7251 22188
rect 7193 22179 7251 22185
rect 7466 22176 7472 22188
rect 7524 22216 7530 22228
rect 10873 22219 10931 22225
rect 7524 22188 7880 22216
rect 7524 22176 7530 22188
rect 3326 22108 3332 22160
rect 3384 22148 3390 22160
rect 3384 22120 4292 22148
rect 3384 22108 3390 22120
rect 3234 22040 3240 22092
rect 3292 22080 3298 22092
rect 4065 22083 4123 22089
rect 4065 22080 4077 22083
rect 3292 22052 4077 22080
rect 3292 22040 3298 22052
rect 4065 22049 4077 22052
rect 4111 22049 4123 22083
rect 4065 22043 4123 22049
rect 4264 22021 4292 22120
rect 4982 22108 4988 22160
rect 5040 22148 5046 22160
rect 6638 22148 6644 22160
rect 5040 22120 6644 22148
rect 5040 22108 5046 22120
rect 4890 22040 4896 22092
rect 4948 22080 4954 22092
rect 5261 22083 5319 22089
rect 5261 22080 5273 22083
rect 4948 22052 5273 22080
rect 4948 22040 4954 22052
rect 5261 22049 5273 22052
rect 5307 22049 5319 22083
rect 5261 22043 5319 22049
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3804 21984 3985 22012
rect 3804 21876 3832 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4157 22015 4215 22021
rect 4157 21981 4169 22015
rect 4203 21981 4215 22015
rect 4157 21975 4215 21981
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4798 22012 4804 22024
rect 4295 21984 4804 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 3878 21904 3884 21956
rect 3936 21944 3942 21956
rect 4172 21944 4200 21975
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 5445 22015 5503 22021
rect 5445 21981 5457 22015
rect 5491 21981 5503 22015
rect 5445 21975 5503 21981
rect 4617 21947 4675 21953
rect 4617 21944 4629 21947
rect 3936 21916 4200 21944
rect 4540 21916 4629 21944
rect 3936 21904 3942 21916
rect 4540 21888 4568 21916
rect 4617 21913 4629 21916
rect 4663 21913 4675 21947
rect 4617 21907 4675 21913
rect 4154 21876 4160 21888
rect 3804 21848 4160 21876
rect 4154 21836 4160 21848
rect 4212 21836 4218 21888
rect 4522 21836 4528 21888
rect 4580 21836 4586 21888
rect 4982 21836 4988 21888
rect 5040 21836 5046 21888
rect 5460 21876 5488 21975
rect 5626 21972 5632 22024
rect 5684 21972 5690 22024
rect 5762 22021 5790 22120
rect 6638 22108 6644 22120
rect 6696 22108 6702 22160
rect 6932 22148 6960 22176
rect 7561 22151 7619 22157
rect 7561 22148 7573 22151
rect 6932 22120 7573 22148
rect 7561 22117 7573 22120
rect 7607 22117 7619 22151
rect 7561 22111 7619 22117
rect 5902 22040 5908 22092
rect 5960 22040 5966 22092
rect 6178 22040 6184 22092
rect 6236 22080 6242 22092
rect 6236 22052 6316 22080
rect 6236 22040 6242 22052
rect 5747 22015 5805 22021
rect 5747 21981 5759 22015
rect 5793 21981 5805 22015
rect 5747 21975 5805 21981
rect 5534 21904 5540 21956
rect 5592 21904 5598 21956
rect 5994 21904 6000 21956
rect 6052 21904 6058 21956
rect 6181 21947 6239 21953
rect 6181 21913 6193 21947
rect 6227 21944 6239 21947
rect 6288 21944 6316 22052
rect 7190 21972 7196 22024
rect 7248 21987 7254 22024
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 7248 21981 7297 21987
rect 7248 21972 7251 21981
rect 6227 21916 6316 21944
rect 7009 21947 7067 21953
rect 6227 21913 6239 21916
rect 6181 21907 6239 21913
rect 7009 21913 7021 21947
rect 7055 21944 7067 21947
rect 7098 21944 7104 21956
rect 7055 21916 7104 21944
rect 7055 21913 7067 21916
rect 7009 21907 7067 21913
rect 7098 21904 7104 21916
rect 7156 21904 7162 21956
rect 7224 21950 7251 21972
rect 7239 21947 7251 21950
rect 7285 21947 7297 21981
rect 7239 21941 7297 21947
rect 7392 21984 7481 22012
rect 6365 21879 6423 21885
rect 6365 21876 6377 21879
rect 5460 21848 6377 21876
rect 6365 21845 6377 21848
rect 6411 21845 6423 21879
rect 6365 21839 6423 21845
rect 6638 21836 6644 21888
rect 6696 21876 6702 21888
rect 7392 21885 7420 21984
rect 7469 21981 7481 21984
rect 7515 21981 7527 22015
rect 7852 22012 7880 22188
rect 10873 22185 10885 22219
rect 10919 22216 10931 22219
rect 11974 22216 11980 22228
rect 10919 22188 11980 22216
rect 10919 22185 10931 22188
rect 10873 22179 10931 22185
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12406 22188 18828 22216
rect 8294 22108 8300 22160
rect 8352 22148 8358 22160
rect 8570 22148 8576 22160
rect 8352 22120 8576 22148
rect 8352 22108 8358 22120
rect 8570 22108 8576 22120
rect 8628 22148 8634 22160
rect 12406 22148 12434 22188
rect 8628 22120 12434 22148
rect 8628 22108 8634 22120
rect 15378 22108 15384 22160
rect 15436 22148 15442 22160
rect 16577 22151 16635 22157
rect 15436 22120 16160 22148
rect 15436 22108 15442 22120
rect 8113 22083 8171 22089
rect 8113 22049 8125 22083
rect 8159 22080 8171 22083
rect 8159 22052 9260 22080
rect 8159 22049 8171 22052
rect 8113 22043 8171 22049
rect 7929 22015 7987 22021
rect 7929 22012 7941 22015
rect 7852 21984 7941 22012
rect 7469 21975 7527 21981
rect 7929 21981 7941 21984
rect 7975 21981 7987 22015
rect 7929 21975 7987 21981
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 9122 22012 9128 22024
rect 8444 21984 9128 22012
rect 8444 21972 8450 21984
rect 9122 21972 9128 21984
rect 9180 21972 9186 22024
rect 9232 22012 9260 22052
rect 9306 22040 9312 22092
rect 9364 22040 9370 22092
rect 11514 22040 11520 22092
rect 11572 22040 11578 22092
rect 11624 22052 12756 22080
rect 11624 22012 11652 22052
rect 9232 21984 11652 22012
rect 12250 21972 12256 22024
rect 12308 21972 12314 22024
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 7742 21904 7748 21956
rect 7800 21944 7806 21956
rect 8941 21947 8999 21953
rect 8941 21944 8953 21947
rect 7800 21916 8953 21944
rect 7800 21904 7806 21916
rect 8941 21913 8953 21916
rect 8987 21913 8999 21947
rect 8941 21907 8999 21913
rect 10318 21904 10324 21956
rect 10376 21944 10382 21956
rect 10870 21944 10876 21956
rect 10376 21916 10876 21944
rect 10376 21904 10382 21916
rect 10870 21904 10876 21916
rect 10928 21944 10934 21956
rect 11241 21947 11299 21953
rect 11241 21944 11253 21947
rect 10928 21916 11253 21944
rect 10928 21904 10934 21916
rect 11241 21913 11253 21916
rect 11287 21913 11299 21947
rect 11241 21907 11299 21913
rect 7377 21879 7435 21885
rect 7377 21876 7389 21879
rect 6696 21848 7389 21876
rect 6696 21836 6702 21848
rect 7377 21845 7389 21848
rect 7423 21845 7435 21879
rect 7377 21839 7435 21845
rect 11330 21836 11336 21888
rect 11388 21836 11394 21888
rect 12268 21885 12296 21972
rect 12544 21944 12572 21975
rect 12618 21972 12624 22024
rect 12676 21972 12682 22024
rect 12728 22021 12756 22052
rect 15028 22052 15792 22080
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 12894 21972 12900 22024
rect 12952 21972 12958 22024
rect 15028 21944 15056 22052
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 15194 22012 15200 22024
rect 15151 21984 15200 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 21981 15347 22015
rect 15289 21975 15347 21981
rect 12544 21916 15056 21944
rect 12253 21879 12311 21885
rect 12253 21845 12265 21879
rect 12299 21845 12311 21879
rect 12253 21839 12311 21845
rect 14918 21836 14924 21888
rect 14976 21876 14982 21888
rect 15304 21876 15332 21975
rect 15764 21944 15792 22052
rect 15838 22040 15844 22092
rect 15896 22040 15902 22092
rect 16132 22089 16160 22120
rect 16577 22117 16589 22151
rect 16623 22148 16635 22151
rect 16758 22148 16764 22160
rect 16623 22120 16764 22148
rect 16623 22117 16635 22120
rect 16577 22111 16635 22117
rect 16758 22108 16764 22120
rect 16816 22108 16822 22160
rect 18141 22151 18199 22157
rect 18141 22117 18153 22151
rect 18187 22148 18199 22151
rect 18690 22148 18696 22160
rect 18187 22120 18696 22148
rect 18187 22117 18199 22120
rect 18141 22111 18199 22117
rect 18690 22108 18696 22120
rect 18748 22108 18754 22160
rect 18800 22148 18828 22188
rect 20346 22176 20352 22228
rect 20404 22216 20410 22228
rect 20625 22219 20683 22225
rect 20625 22216 20637 22219
rect 20404 22188 20637 22216
rect 20404 22176 20410 22188
rect 20625 22185 20637 22188
rect 20671 22185 20683 22219
rect 20625 22179 20683 22185
rect 20806 22176 20812 22228
rect 20864 22216 20870 22228
rect 20901 22219 20959 22225
rect 20901 22216 20913 22219
rect 20864 22188 20913 22216
rect 20864 22176 20870 22188
rect 20901 22185 20913 22188
rect 20947 22185 20959 22219
rect 20901 22179 20959 22185
rect 20990 22176 20996 22228
rect 21048 22176 21054 22228
rect 21085 22219 21143 22225
rect 21085 22185 21097 22219
rect 21131 22216 21143 22219
rect 21818 22216 21824 22228
rect 21131 22188 21824 22216
rect 21131 22185 21143 22188
rect 21085 22179 21143 22185
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 25498 22216 25504 22228
rect 22066 22188 25504 22216
rect 22066 22148 22094 22188
rect 25498 22176 25504 22188
rect 25556 22176 25562 22228
rect 28350 22216 28356 22228
rect 25608 22188 28356 22216
rect 18800 22120 22094 22148
rect 22186 22108 22192 22160
rect 22244 22148 22250 22160
rect 22370 22148 22376 22160
rect 22244 22120 22376 22148
rect 22244 22108 22250 22120
rect 22370 22108 22376 22120
rect 22428 22108 22434 22160
rect 24394 22108 24400 22160
rect 24452 22108 24458 22160
rect 24946 22108 24952 22160
rect 25004 22148 25010 22160
rect 25608 22148 25636 22188
rect 28350 22176 28356 22188
rect 28408 22176 28414 22228
rect 29181 22219 29239 22225
rect 29181 22185 29193 22219
rect 29227 22216 29239 22219
rect 29454 22216 29460 22228
rect 29227 22188 29460 22216
rect 29227 22185 29239 22188
rect 29181 22179 29239 22185
rect 29454 22176 29460 22188
rect 29512 22176 29518 22228
rect 30374 22176 30380 22228
rect 30432 22216 30438 22228
rect 31389 22219 31447 22225
rect 31389 22216 31401 22219
rect 30432 22188 31401 22216
rect 30432 22176 30438 22188
rect 31389 22185 31401 22188
rect 31435 22185 31447 22219
rect 31389 22179 31447 22185
rect 31478 22176 31484 22228
rect 31536 22216 31542 22228
rect 31536 22188 32260 22216
rect 31536 22176 31542 22188
rect 25004 22120 25636 22148
rect 25685 22151 25743 22157
rect 25004 22108 25010 22120
rect 25685 22117 25697 22151
rect 25731 22148 25743 22151
rect 27614 22148 27620 22160
rect 25731 22120 27620 22148
rect 25731 22117 25743 22120
rect 25685 22111 25743 22117
rect 27614 22108 27620 22120
rect 27672 22108 27678 22160
rect 28077 22151 28135 22157
rect 28077 22117 28089 22151
rect 28123 22148 28135 22151
rect 28166 22148 28172 22160
rect 28123 22120 28172 22148
rect 28123 22117 28135 22120
rect 28077 22111 28135 22117
rect 28166 22108 28172 22120
rect 28224 22108 28230 22160
rect 16117 22083 16175 22089
rect 16117 22049 16129 22083
rect 16163 22049 16175 22083
rect 16117 22043 16175 22049
rect 16500 22052 16804 22080
rect 16500 22021 16528 22052
rect 16776 22024 16804 22052
rect 17586 22040 17592 22092
rect 17644 22080 17650 22092
rect 18785 22083 18843 22089
rect 17644 22052 18368 22080
rect 17644 22040 17650 22052
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 16758 21972 16764 22024
rect 16816 21972 16822 22024
rect 16850 21972 16856 22024
rect 16908 21972 16914 22024
rect 17126 21972 17132 22024
rect 17184 21972 17190 22024
rect 18049 22015 18107 22021
rect 18049 21981 18061 22015
rect 18095 22012 18107 22015
rect 18138 22012 18144 22024
rect 18095 21984 18144 22012
rect 18095 21981 18107 21984
rect 18049 21975 18107 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 18340 22021 18368 22052
rect 18785 22049 18797 22083
rect 18831 22080 18843 22083
rect 19058 22080 19064 22092
rect 18831 22052 19064 22080
rect 18831 22049 18843 22052
rect 18785 22043 18843 22049
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 22649 22083 22707 22089
rect 20312 22052 21404 22080
rect 20312 22040 20318 22052
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 21981 18383 22015
rect 18325 21975 18383 21981
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 22012 21235 22015
rect 21266 22012 21272 22024
rect 21223 21984 21272 22012
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 21266 21972 21272 21984
rect 21324 21972 21330 22024
rect 21376 22021 21404 22052
rect 22649 22049 22661 22083
rect 22695 22080 22707 22083
rect 23198 22080 23204 22092
rect 22695 22052 23204 22080
rect 22695 22049 22707 22052
rect 22649 22043 22707 22049
rect 23198 22040 23204 22052
rect 23256 22040 23262 22092
rect 26881 22083 26939 22089
rect 24688 22052 25636 22080
rect 21361 22015 21419 22021
rect 21361 21981 21373 22015
rect 21407 21981 21419 22015
rect 21361 21975 21419 21981
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 21545 22015 21603 22021
rect 21545 22012 21557 22015
rect 21508 21984 21557 22012
rect 21508 21972 21514 21984
rect 21545 21981 21557 21984
rect 21591 21981 21603 22015
rect 21545 21975 21603 21981
rect 21634 21972 21640 22024
rect 21692 22012 21698 22024
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 21692 21984 22017 22012
rect 21692 21972 21698 21984
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22189 22015 22247 22021
rect 22189 22012 22201 22015
rect 22152 21984 22201 22012
rect 22152 21972 22158 21984
rect 22189 21981 22201 21984
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 22278 21972 22284 22024
rect 22336 21972 22342 22024
rect 24688 22021 24716 22052
rect 24673 22015 24731 22021
rect 22374 21993 22432 21999
rect 22374 21959 22386 21993
rect 22420 21959 22432 21993
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 22374 21956 22432 21959
rect 15764 21916 22325 21944
rect 14976 21848 15332 21876
rect 14976 21836 14982 21848
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 21450 21876 21456 21888
rect 19484 21848 21456 21876
rect 19484 21836 19490 21848
rect 21450 21836 21456 21848
rect 21508 21836 21514 21888
rect 21729 21879 21787 21885
rect 21729 21845 21741 21879
rect 21775 21876 21787 21879
rect 22186 21876 22192 21888
rect 21775 21848 22192 21876
rect 21775 21845 21787 21848
rect 21729 21839 21787 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22297 21876 22325 21916
rect 22370 21904 22376 21956
rect 22428 21904 22434 21956
rect 22830 21904 22836 21956
rect 22888 21944 22894 21956
rect 24780 21944 24808 21975
rect 24854 21972 24860 22024
rect 24912 21972 24918 22024
rect 24946 21972 24952 22024
rect 25004 22012 25010 22024
rect 25041 22015 25099 22021
rect 25041 22012 25053 22015
rect 25004 21984 25053 22012
rect 25004 21972 25010 21984
rect 25041 21981 25053 21984
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 25130 21972 25136 22024
rect 25188 21972 25194 22024
rect 25406 21972 25412 22024
rect 25464 21972 25470 22024
rect 25498 21972 25504 22024
rect 25556 21972 25562 22024
rect 25608 22012 25636 22052
rect 26881 22049 26893 22083
rect 26927 22080 26939 22083
rect 26970 22080 26976 22092
rect 26927 22052 26976 22080
rect 26927 22049 26939 22052
rect 26881 22043 26939 22049
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 27540 22052 28212 22080
rect 25608 21984 25912 22012
rect 22888 21916 24808 21944
rect 22888 21904 22894 21916
rect 25314 21904 25320 21956
rect 25372 21944 25378 21956
rect 25682 21944 25688 21956
rect 25372 21916 25688 21944
rect 25372 21904 25378 21916
rect 25682 21904 25688 21916
rect 25740 21904 25746 21956
rect 25884 21944 25912 21984
rect 25958 21972 25964 22024
rect 26016 22012 26022 22024
rect 27065 22015 27123 22021
rect 27065 22012 27077 22015
rect 26016 21984 27077 22012
rect 26016 21972 26022 21984
rect 27065 21981 27077 21984
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 27338 21972 27344 22024
rect 27396 22012 27402 22024
rect 27540 22021 27568 22052
rect 27525 22015 27583 22021
rect 27525 22012 27537 22015
rect 27396 21984 27537 22012
rect 27396 21972 27402 21984
rect 27525 21981 27537 21984
rect 27571 21981 27583 22015
rect 27525 21975 27583 21981
rect 27893 22015 27951 22021
rect 27893 21981 27905 22015
rect 27939 22009 27951 22015
rect 27982 22009 27988 22024
rect 27939 21981 27988 22009
rect 27893 21975 27951 21981
rect 27982 21972 27988 21981
rect 28040 21972 28046 22024
rect 28184 22021 28212 22052
rect 28810 22040 28816 22092
rect 28868 22040 28874 22092
rect 28169 22015 28227 22021
rect 28169 21981 28181 22015
rect 28215 21981 28227 22015
rect 28169 21975 28227 21981
rect 28534 21972 28540 22024
rect 28592 21972 28598 22024
rect 28718 21972 28724 22024
rect 28776 22012 28782 22024
rect 28997 22015 29055 22021
rect 28997 22012 29009 22015
rect 28776 21984 29009 22012
rect 28776 21972 28782 21984
rect 28997 21981 29009 21984
rect 29043 21981 29055 22015
rect 29472 22012 29500 22176
rect 30650 22148 30656 22160
rect 30576 22120 30656 22148
rect 30576 22089 30604 22120
rect 30650 22108 30656 22120
rect 30708 22148 30714 22160
rect 31570 22148 31576 22160
rect 30708 22120 31576 22148
rect 30708 22108 30714 22120
rect 31570 22108 31576 22120
rect 31628 22108 31634 22160
rect 31665 22151 31723 22157
rect 31665 22117 31677 22151
rect 31711 22148 31723 22151
rect 31938 22148 31944 22160
rect 31711 22120 31944 22148
rect 31711 22117 31723 22120
rect 31665 22111 31723 22117
rect 31938 22108 31944 22120
rect 31996 22108 32002 22160
rect 32033 22151 32091 22157
rect 32033 22117 32045 22151
rect 32079 22148 32091 22151
rect 32079 22120 32113 22148
rect 32079 22117 32091 22120
rect 32033 22111 32091 22117
rect 30561 22083 30619 22089
rect 29662 22052 30512 22080
rect 29549 22015 29607 22021
rect 29549 22012 29561 22015
rect 29472 21984 29561 22012
rect 28997 21975 29055 21981
rect 29549 21981 29561 21984
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 26878 21944 26884 21956
rect 25884 21916 26884 21944
rect 26878 21904 26884 21916
rect 26936 21904 26942 21956
rect 27709 21947 27767 21953
rect 27709 21944 27721 21947
rect 26988 21916 27721 21944
rect 23750 21876 23756 21888
rect 22297 21848 23756 21876
rect 23750 21836 23756 21848
rect 23808 21876 23814 21888
rect 26988 21876 27016 21916
rect 27709 21913 27721 21916
rect 27755 21913 27767 21947
rect 27709 21907 27767 21913
rect 23808 21848 27016 21876
rect 27249 21879 27307 21885
rect 23808 21836 23814 21848
rect 27249 21845 27261 21879
rect 27295 21876 27307 21879
rect 27614 21876 27620 21888
rect 27295 21848 27620 21876
rect 27295 21845 27307 21848
rect 27249 21839 27307 21845
rect 27614 21836 27620 21848
rect 27672 21836 27678 21888
rect 27724 21876 27752 21907
rect 27798 21904 27804 21956
rect 27856 21904 27862 21956
rect 27908 21916 28304 21944
rect 27908 21876 27936 21916
rect 27724 21848 27936 21876
rect 28276 21876 28304 21916
rect 28350 21904 28356 21956
rect 28408 21904 28414 21956
rect 28442 21904 28448 21956
rect 28500 21904 28506 21956
rect 29662 21944 29690 22052
rect 29730 21972 29736 22024
rect 29788 21972 29794 22024
rect 29825 22015 29883 22021
rect 29825 21981 29837 22015
rect 29871 22012 29883 22015
rect 29871 21984 30328 22012
rect 29871 21981 29883 21984
rect 29825 21975 29883 21981
rect 28552 21916 29690 21944
rect 28552 21876 28580 21916
rect 28276 21848 28580 21876
rect 28721 21879 28779 21885
rect 28721 21845 28733 21879
rect 28767 21876 28779 21879
rect 28994 21876 29000 21888
rect 28767 21848 29000 21876
rect 28767 21845 28779 21848
rect 28721 21839 28779 21845
rect 28994 21836 29000 21848
rect 29052 21836 29058 21888
rect 29086 21836 29092 21888
rect 29144 21876 29150 21888
rect 29647 21879 29705 21885
rect 29647 21876 29659 21879
rect 29144 21848 29659 21876
rect 29144 21836 29150 21848
rect 29647 21845 29659 21848
rect 29693 21845 29705 21879
rect 29647 21839 29705 21845
rect 29914 21836 29920 21888
rect 29972 21876 29978 21888
rect 30009 21879 30067 21885
rect 30009 21876 30021 21879
rect 29972 21848 30021 21876
rect 29972 21836 29978 21848
rect 30009 21845 30021 21848
rect 30055 21845 30067 21879
rect 30300 21876 30328 21984
rect 30374 21972 30380 22024
rect 30432 21972 30438 22024
rect 30484 21944 30512 22052
rect 30561 22049 30573 22083
rect 30607 22080 30619 22083
rect 32048 22080 32076 22111
rect 30607 22052 30641 22080
rect 31036 22052 32076 22080
rect 32232 22080 32260 22188
rect 33704 22188 35204 22216
rect 32306 22108 32312 22160
rect 32364 22148 32370 22160
rect 32364 22120 32628 22148
rect 32364 22108 32370 22120
rect 32600 22080 32628 22120
rect 32674 22108 32680 22160
rect 32732 22148 32738 22160
rect 33704 22148 33732 22188
rect 35176 22148 35204 22188
rect 35434 22148 35440 22160
rect 32732 22120 33732 22148
rect 32732 22108 32738 22120
rect 32232 22052 32352 22080
rect 32600 22052 33456 22080
rect 30607 22049 30619 22052
rect 30561 22043 30619 22049
rect 31036 22021 31064 22052
rect 31021 22015 31079 22021
rect 31021 21981 31033 22015
rect 31067 21981 31079 22015
rect 31021 21975 31079 21981
rect 31202 21972 31208 22024
rect 31260 21972 31266 22024
rect 31570 21972 31576 22024
rect 31628 21972 31634 22024
rect 31757 22015 31815 22021
rect 31757 21981 31769 22015
rect 31803 21981 31815 22015
rect 31757 21975 31815 21981
rect 31772 21944 31800 21975
rect 31846 21972 31852 22024
rect 31904 21972 31910 22024
rect 32030 21972 32036 22024
rect 32088 21972 32094 22024
rect 32122 21972 32128 22024
rect 32180 22012 32186 22024
rect 32324 22021 32352 22052
rect 32217 22015 32275 22021
rect 32217 22012 32229 22015
rect 32180 21984 32229 22012
rect 32180 21972 32186 21984
rect 32217 21981 32229 21984
rect 32263 21981 32275 22015
rect 32217 21975 32275 21981
rect 32309 22015 32367 22021
rect 32309 21981 32321 22015
rect 32355 21981 32367 22015
rect 32309 21975 32367 21981
rect 32398 21972 32404 22024
rect 32456 22012 32462 22024
rect 32677 22015 32735 22021
rect 32677 22012 32689 22015
rect 32456 21984 32689 22012
rect 32456 21972 32462 21984
rect 32677 21981 32689 21984
rect 32723 21981 32735 22015
rect 32677 21975 32735 21981
rect 32769 22015 32827 22021
rect 32769 21981 32781 22015
rect 32815 21981 32827 22015
rect 32769 21975 32827 21981
rect 32416 21944 32444 21972
rect 30484 21916 31248 21944
rect 31772 21916 31892 21944
rect 30466 21876 30472 21888
rect 30300 21848 30472 21876
rect 30009 21839 30067 21845
rect 30466 21836 30472 21848
rect 30524 21836 30530 21888
rect 31220 21885 31248 21916
rect 31205 21879 31263 21885
rect 31205 21845 31217 21879
rect 31251 21876 31263 21879
rect 31294 21876 31300 21888
rect 31251 21848 31300 21876
rect 31251 21845 31263 21848
rect 31205 21839 31263 21845
rect 31294 21836 31300 21848
rect 31352 21836 31358 21888
rect 31864 21876 31892 21916
rect 32324 21916 32444 21944
rect 32324 21876 32352 21916
rect 32784 21888 32812 21975
rect 32858 21972 32864 22024
rect 32916 21972 32922 22024
rect 33045 22015 33103 22021
rect 33045 21981 33057 22015
rect 33091 22012 33103 22015
rect 33134 22012 33140 22024
rect 33091 21984 33140 22012
rect 33091 21981 33103 21984
rect 33045 21975 33103 21981
rect 33134 21972 33140 21984
rect 33192 21972 33198 22024
rect 31864 21848 32352 21876
rect 32401 21879 32459 21885
rect 32401 21845 32413 21879
rect 32447 21876 32459 21879
rect 32490 21876 32496 21888
rect 32447 21848 32496 21876
rect 32447 21845 32459 21848
rect 32401 21839 32459 21845
rect 32490 21836 32496 21848
rect 32548 21836 32554 21888
rect 32766 21836 32772 21888
rect 32824 21876 32830 21888
rect 33137 21879 33195 21885
rect 33137 21876 33149 21879
rect 32824 21848 33149 21876
rect 32824 21836 32830 21848
rect 33137 21845 33149 21848
rect 33183 21845 33195 21879
rect 33428 21876 33456 22052
rect 33502 22040 33508 22092
rect 33560 22040 33566 22092
rect 33704 22089 33732 22120
rect 34348 22120 34744 22148
rect 35176 22120 35440 22148
rect 33689 22083 33747 22089
rect 33689 22049 33701 22083
rect 33735 22080 33747 22083
rect 34348 22080 34376 22120
rect 33735 22052 33769 22080
rect 34164 22052 34376 22080
rect 34425 22083 34483 22089
rect 33735 22049 33747 22052
rect 33689 22043 33747 22049
rect 33520 21953 33548 22040
rect 34164 22021 34192 22052
rect 34425 22049 34437 22083
rect 34471 22080 34483 22083
rect 34606 22080 34612 22092
rect 34471 22052 34612 22080
rect 34471 22049 34483 22052
rect 34425 22043 34483 22049
rect 34606 22040 34612 22052
rect 34664 22040 34670 22092
rect 34149 22015 34207 22021
rect 34149 22012 34161 22015
rect 33888 21984 34161 22012
rect 33888 21956 33916 21984
rect 34149 21981 34161 21984
rect 34195 21981 34207 22015
rect 34149 21975 34207 21981
rect 34241 22015 34299 22021
rect 34241 21981 34253 22015
rect 34287 21981 34299 22015
rect 34241 21975 34299 21981
rect 33505 21947 33563 21953
rect 33505 21913 33517 21947
rect 33551 21913 33563 21947
rect 33505 21907 33563 21913
rect 33870 21904 33876 21956
rect 33928 21904 33934 21956
rect 34256 21944 34284 21975
rect 34330 21972 34336 22024
rect 34388 21972 34394 22024
rect 34716 22012 34744 22120
rect 35268 22089 35296 22120
rect 35434 22108 35440 22120
rect 35492 22108 35498 22160
rect 35253 22083 35311 22089
rect 35253 22049 35265 22083
rect 35299 22049 35311 22083
rect 35253 22043 35311 22049
rect 35529 22083 35587 22089
rect 35529 22049 35541 22083
rect 35575 22080 35587 22083
rect 35802 22080 35808 22092
rect 35575 22052 35808 22080
rect 35575 22049 35587 22052
rect 35529 22043 35587 22049
rect 35802 22040 35808 22052
rect 35860 22040 35866 22092
rect 35989 22015 36047 22021
rect 35989 22012 36001 22015
rect 34716 21984 36001 22012
rect 35989 21981 36001 21984
rect 36035 21981 36047 22015
rect 35989 21975 36047 21981
rect 35894 21944 35900 21956
rect 34256 21916 35900 21944
rect 35894 21904 35900 21916
rect 35952 21904 35958 21956
rect 33597 21879 33655 21885
rect 33597 21876 33609 21879
rect 33428 21848 33609 21876
rect 33137 21839 33195 21845
rect 33597 21845 33609 21848
rect 33643 21876 33655 21879
rect 33965 21879 34023 21885
rect 33965 21876 33977 21879
rect 33643 21848 33977 21876
rect 33643 21845 33655 21848
rect 33597 21839 33655 21845
rect 33965 21845 33977 21848
rect 34011 21845 34023 21879
rect 33965 21839 34023 21845
rect 34146 21836 34152 21888
rect 34204 21876 34210 21888
rect 34701 21879 34759 21885
rect 34701 21876 34713 21879
rect 34204 21848 34713 21876
rect 34204 21836 34210 21848
rect 34701 21845 34713 21848
rect 34747 21845 34759 21879
rect 34701 21839 34759 21845
rect 34790 21836 34796 21888
rect 34848 21876 34854 21888
rect 35069 21879 35127 21885
rect 35069 21876 35081 21879
rect 34848 21848 35081 21876
rect 34848 21836 34854 21848
rect 35069 21845 35081 21848
rect 35115 21845 35127 21879
rect 35069 21839 35127 21845
rect 35161 21879 35219 21885
rect 35161 21845 35173 21879
rect 35207 21876 35219 21879
rect 35805 21879 35863 21885
rect 35805 21876 35817 21879
rect 35207 21848 35817 21876
rect 35207 21845 35219 21848
rect 35161 21839 35219 21845
rect 35805 21845 35817 21848
rect 35851 21845 35863 21879
rect 35805 21839 35863 21845
rect 1104 21786 38272 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38272 21786
rect 1104 21712 38272 21734
rect 2409 21675 2467 21681
rect 2409 21641 2421 21675
rect 2455 21672 2467 21675
rect 2590 21672 2596 21684
rect 2455 21644 2596 21672
rect 2455 21641 2467 21644
rect 2409 21635 2467 21641
rect 2590 21632 2596 21644
rect 2648 21632 2654 21684
rect 5902 21632 5908 21684
rect 5960 21672 5966 21684
rect 7006 21672 7012 21684
rect 5960 21644 7012 21672
rect 5960 21632 5966 21644
rect 7006 21632 7012 21644
rect 7064 21632 7070 21684
rect 8202 21632 8208 21684
rect 8260 21672 8266 21684
rect 9585 21675 9643 21681
rect 9585 21672 9597 21675
rect 8260 21644 9597 21672
rect 8260 21632 8266 21644
rect 9585 21641 9597 21644
rect 9631 21641 9643 21675
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 9585 21635 9643 21641
rect 9692 21644 10241 21672
rect 2498 21604 2504 21616
rect 2240 21576 2504 21604
rect 2240 21545 2268 21576
rect 2498 21564 2504 21576
rect 2556 21604 2562 21616
rect 2556 21576 4016 21604
rect 2556 21564 2562 21576
rect 3988 21548 4016 21576
rect 5258 21564 5264 21616
rect 5316 21604 5322 21616
rect 5353 21607 5411 21613
rect 5353 21604 5365 21607
rect 5316 21576 5365 21604
rect 5316 21564 5322 21576
rect 5353 21573 5365 21576
rect 5399 21573 5411 21607
rect 5994 21604 6000 21616
rect 5353 21567 5411 21573
rect 5644 21576 6000 21604
rect 2225 21539 2283 21545
rect 2225 21505 2237 21539
rect 2271 21505 2283 21539
rect 2225 21499 2283 21505
rect 2406 21496 2412 21548
rect 2464 21496 2470 21548
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 3878 21536 3884 21548
rect 2915 21508 3884 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 3878 21496 3884 21508
rect 3936 21496 3942 21548
rect 3970 21496 3976 21548
rect 4028 21536 4034 21548
rect 4522 21536 4528 21548
rect 4028 21508 4528 21536
rect 4028 21496 4034 21508
rect 4522 21496 4528 21508
rect 4580 21536 4586 21548
rect 5169 21539 5227 21545
rect 5169 21536 5181 21539
rect 4580 21508 5181 21536
rect 4580 21496 4586 21508
rect 5169 21505 5181 21508
rect 5215 21505 5227 21539
rect 5169 21499 5227 21505
rect 2958 21428 2964 21480
rect 3016 21428 3022 21480
rect 3050 21428 3056 21480
rect 3108 21428 3114 21480
rect 5184 21400 5212 21499
rect 5368 21468 5396 21567
rect 5644 21545 5672 21576
rect 5994 21564 6000 21576
rect 6052 21604 6058 21616
rect 6638 21604 6644 21616
rect 6052 21576 6644 21604
rect 6052 21564 6058 21576
rect 6638 21564 6644 21576
rect 6696 21564 6702 21616
rect 8846 21564 8852 21616
rect 8904 21604 8910 21616
rect 9692 21604 9720 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 10229 21635 10287 21641
rect 13354 21632 13360 21684
rect 13412 21632 13418 21684
rect 15013 21675 15071 21681
rect 15013 21641 15025 21675
rect 15059 21672 15071 21675
rect 15470 21672 15476 21684
rect 15059 21644 15476 21672
rect 15059 21641 15071 21644
rect 15013 21635 15071 21641
rect 15470 21632 15476 21644
rect 15528 21632 15534 21684
rect 16758 21632 16764 21684
rect 16816 21672 16822 21684
rect 16853 21675 16911 21681
rect 16853 21672 16865 21675
rect 16816 21644 16865 21672
rect 16816 21632 16822 21644
rect 16853 21641 16865 21644
rect 16899 21672 16911 21675
rect 17678 21672 17684 21684
rect 16899 21644 17684 21672
rect 16899 21641 16911 21644
rect 16853 21635 16911 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 18969 21675 19027 21681
rect 18969 21641 18981 21675
rect 19015 21672 19027 21675
rect 19978 21672 19984 21684
rect 19015 21644 19984 21672
rect 19015 21641 19027 21644
rect 18969 21635 19027 21641
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 20809 21675 20867 21681
rect 20809 21641 20821 21675
rect 20855 21672 20867 21675
rect 22094 21672 22100 21684
rect 20855 21644 22100 21672
rect 20855 21641 20867 21644
rect 20809 21635 20867 21641
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 25130 21632 25136 21684
rect 25188 21672 25194 21684
rect 25958 21672 25964 21684
rect 25188 21644 25964 21672
rect 25188 21632 25194 21644
rect 25958 21632 25964 21644
rect 26016 21672 26022 21684
rect 26145 21675 26203 21681
rect 26145 21672 26157 21675
rect 26016 21644 26157 21672
rect 26016 21632 26022 21644
rect 26145 21641 26157 21644
rect 26191 21641 26203 21675
rect 26145 21635 26203 21641
rect 27890 21632 27896 21684
rect 27948 21632 27954 21684
rect 29730 21632 29736 21684
rect 29788 21632 29794 21684
rect 30098 21632 30104 21684
rect 30156 21672 30162 21684
rect 30193 21675 30251 21681
rect 30193 21672 30205 21675
rect 30156 21644 30205 21672
rect 30156 21632 30162 21644
rect 30193 21641 30205 21644
rect 30239 21641 30251 21675
rect 30193 21635 30251 21641
rect 31202 21632 31208 21684
rect 31260 21672 31266 21684
rect 31389 21675 31447 21681
rect 31389 21672 31401 21675
rect 31260 21644 31401 21672
rect 31260 21632 31266 21644
rect 31389 21641 31401 21644
rect 31435 21641 31447 21675
rect 31389 21635 31447 21641
rect 32122 21632 32128 21684
rect 32180 21632 32186 21684
rect 32398 21632 32404 21684
rect 32456 21632 32462 21684
rect 32858 21632 32864 21684
rect 32916 21632 32922 21684
rect 34146 21632 34152 21684
rect 34204 21632 34210 21684
rect 34330 21632 34336 21684
rect 34388 21672 34394 21684
rect 34793 21675 34851 21681
rect 34793 21672 34805 21675
rect 34388 21644 34805 21672
rect 34388 21632 34394 21644
rect 34793 21641 34805 21644
rect 34839 21641 34851 21675
rect 34793 21635 34851 21641
rect 8904 21576 9720 21604
rect 12805 21607 12863 21613
rect 8904 21564 8910 21576
rect 12805 21573 12817 21607
rect 12851 21604 12863 21607
rect 12894 21604 12900 21616
rect 12851 21576 12900 21604
rect 12851 21573 12863 21576
rect 12805 21567 12863 21573
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21505 5687 21539
rect 5629 21499 5687 21505
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 6178 21536 6184 21548
rect 5859 21508 6184 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 5828 21468 5856 21499
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 5368 21440 5856 21468
rect 7742 21400 7748 21412
rect 5184 21372 7748 21400
rect 7742 21360 7748 21372
rect 7800 21360 7806 21412
rect 2498 21292 2504 21344
rect 2556 21292 2562 21344
rect 5534 21292 5540 21344
rect 5592 21292 5598 21344
rect 5718 21292 5724 21344
rect 5776 21292 5782 21344
rect 9232 21332 9260 21499
rect 9306 21496 9312 21548
rect 9364 21496 9370 21548
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21505 9459 21539
rect 9401 21499 9459 21505
rect 9677 21539 9735 21545
rect 9677 21505 9689 21539
rect 9723 21534 9735 21539
rect 9766 21534 9772 21548
rect 9723 21506 9772 21534
rect 9723 21505 9735 21506
rect 9677 21499 9735 21505
rect 9416 21468 9444 21499
rect 9766 21496 9772 21506
rect 9824 21496 9830 21548
rect 9858 21496 9864 21548
rect 9916 21496 9922 21548
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 10045 21539 10103 21545
rect 10045 21505 10057 21539
rect 10091 21536 10103 21539
rect 10686 21536 10692 21548
rect 10091 21508 10692 21536
rect 10091 21505 10103 21508
rect 10045 21499 10103 21505
rect 10060 21468 10088 21499
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 9416 21440 10088 21468
rect 10318 21428 10324 21480
rect 10376 21468 10382 21480
rect 12820 21468 12848 21567
rect 12894 21564 12900 21576
rect 12952 21604 12958 21616
rect 14829 21607 14887 21613
rect 12952 21576 14596 21604
rect 12952 21564 12958 21576
rect 13354 21496 13360 21548
rect 13412 21496 13418 21548
rect 10376 21440 12848 21468
rect 10376 21428 10382 21440
rect 12894 21428 12900 21480
rect 12952 21468 12958 21480
rect 13449 21471 13507 21477
rect 13449 21468 13461 21471
rect 12952 21440 13461 21468
rect 12952 21428 12958 21440
rect 13449 21437 13461 21440
rect 13495 21437 13507 21471
rect 14568 21468 14596 21576
rect 14829 21573 14841 21607
rect 14875 21604 14887 21607
rect 15194 21604 15200 21616
rect 14875 21576 15200 21604
rect 14875 21573 14887 21576
rect 14829 21567 14887 21573
rect 15194 21564 15200 21576
rect 15252 21564 15258 21616
rect 16390 21564 16396 21616
rect 16448 21564 16454 21616
rect 18509 21607 18567 21613
rect 16500 21576 18092 21604
rect 14645 21539 14703 21545
rect 14645 21505 14657 21539
rect 14691 21536 14703 21539
rect 14918 21536 14924 21548
rect 14691 21508 14924 21536
rect 14691 21505 14703 21508
rect 14645 21499 14703 21505
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 15010 21496 15016 21548
rect 15068 21536 15074 21548
rect 16022 21536 16028 21548
rect 15068 21508 16028 21536
rect 15068 21496 15074 21508
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 16206 21496 16212 21548
rect 16264 21496 16270 21548
rect 16500 21468 16528 21576
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16853 21539 16911 21545
rect 16715 21508 16804 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 14568 21440 16528 21468
rect 13449 21431 13507 21437
rect 16776 21412 16804 21508
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 17405 21539 17463 21545
rect 16899 21508 17264 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 17236 21412 17264 21508
rect 17405 21505 17417 21539
rect 17451 21505 17463 21539
rect 17405 21499 17463 21505
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 9398 21360 9404 21412
rect 9456 21400 9462 21412
rect 9456 21372 9904 21400
rect 9456 21360 9462 21372
rect 9766 21332 9772 21344
rect 9232 21304 9772 21332
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 9876 21332 9904 21372
rect 16758 21360 16764 21412
rect 16816 21360 16822 21412
rect 17218 21360 17224 21412
rect 17276 21360 17282 21412
rect 17420 21400 17448 21499
rect 17586 21496 17592 21548
rect 17644 21536 17650 21548
rect 17770 21536 17776 21548
rect 17644 21508 17776 21536
rect 17644 21496 17650 21508
rect 17770 21496 17776 21508
rect 17828 21536 17834 21548
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 17828 21508 17877 21536
rect 17828 21496 17834 21508
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 17954 21496 17960 21548
rect 18012 21496 18018 21548
rect 18064 21536 18092 21576
rect 18509 21573 18521 21607
rect 18555 21604 18567 21607
rect 18874 21604 18880 21616
rect 18555 21576 18880 21604
rect 18555 21573 18567 21576
rect 18509 21567 18567 21573
rect 18874 21564 18880 21576
rect 18932 21564 18938 21616
rect 18984 21576 20208 21604
rect 18984 21536 19012 21576
rect 18064 21508 19012 21536
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 19337 21539 19395 21545
rect 19337 21536 19349 21539
rect 19116 21508 19349 21536
rect 19116 21496 19122 21508
rect 19337 21505 19349 21508
rect 19383 21505 19395 21539
rect 19337 21499 19395 21505
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21505 19763 21539
rect 19705 21499 19763 21505
rect 19153 21471 19211 21477
rect 19153 21468 19165 21471
rect 18340 21440 19165 21468
rect 17420 21372 17724 21400
rect 17696 21344 17724 21372
rect 17954 21360 17960 21412
rect 18012 21400 18018 21412
rect 18340 21400 18368 21440
rect 19153 21437 19165 21440
rect 19199 21468 19211 21471
rect 19426 21468 19432 21480
rect 19199 21440 19432 21468
rect 19199 21437 19211 21440
rect 19153 21431 19211 21437
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 19613 21471 19671 21477
rect 19613 21437 19625 21471
rect 19659 21437 19671 21471
rect 19613 21431 19671 21437
rect 18012 21372 18368 21400
rect 18012 21360 18018 21372
rect 18874 21360 18880 21412
rect 18932 21400 18938 21412
rect 19628 21400 19656 21431
rect 19720 21412 19748 21499
rect 20180 21412 20208 21576
rect 20714 21564 20720 21616
rect 20772 21604 20778 21616
rect 21266 21604 21272 21616
rect 20772 21576 21272 21604
rect 20772 21564 20778 21576
rect 21266 21564 21272 21576
rect 21324 21604 21330 21616
rect 21913 21607 21971 21613
rect 21913 21604 21925 21607
rect 21324 21576 21925 21604
rect 21324 21564 21330 21576
rect 21913 21573 21925 21576
rect 21959 21573 21971 21607
rect 21913 21567 21971 21573
rect 22281 21607 22339 21613
rect 22281 21573 22293 21607
rect 22327 21604 22339 21607
rect 22646 21604 22652 21616
rect 22327 21576 22652 21604
rect 22327 21573 22339 21576
rect 22281 21567 22339 21573
rect 22646 21564 22652 21576
rect 22704 21564 22710 21616
rect 24670 21604 24676 21616
rect 22940 21576 24676 21604
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20732 21508 21097 21536
rect 20732 21480 20760 21508
rect 21085 21505 21097 21508
rect 21131 21505 21143 21539
rect 21085 21499 21143 21505
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22370 21536 22376 21548
rect 22244 21508 22376 21536
rect 22244 21496 22250 21508
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 22830 21496 22836 21548
rect 22888 21496 22894 21548
rect 22940 21545 22968 21576
rect 24670 21564 24676 21576
rect 24728 21604 24734 21616
rect 27525 21607 27583 21613
rect 27525 21604 27537 21607
rect 24728 21576 27537 21604
rect 24728 21564 24734 21576
rect 27525 21573 27537 21576
rect 27571 21604 27583 21607
rect 27571 21576 28580 21604
rect 27571 21573 27583 21576
rect 27525 21567 27583 21573
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21505 22983 21539
rect 22925 21499 22983 21505
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21505 23075 21539
rect 23017 21499 23075 21505
rect 20714 21428 20720 21480
rect 20772 21428 20778 21480
rect 20806 21428 20812 21480
rect 20864 21468 20870 21480
rect 20993 21471 21051 21477
rect 20993 21468 21005 21471
rect 20864 21440 21005 21468
rect 20864 21428 20870 21440
rect 20993 21437 21005 21440
rect 21039 21437 21051 21471
rect 21177 21471 21235 21477
rect 21177 21468 21189 21471
rect 20993 21431 21051 21437
rect 21100 21440 21189 21468
rect 21100 21412 21128 21440
rect 21177 21437 21189 21440
rect 21223 21437 21235 21471
rect 21177 21431 21235 21437
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21468 21327 21471
rect 21358 21468 21364 21480
rect 21315 21440 21364 21468
rect 21315 21437 21327 21440
rect 21269 21431 21327 21437
rect 21358 21428 21364 21440
rect 21416 21468 21422 21480
rect 22097 21471 22155 21477
rect 22097 21468 22109 21471
rect 21416 21440 22109 21468
rect 21416 21428 21422 21440
rect 22097 21437 22109 21440
rect 22143 21468 22155 21471
rect 22278 21468 22284 21480
rect 22143 21440 22284 21468
rect 22143 21437 22155 21440
rect 22097 21431 22155 21437
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 22848 21468 22876 21496
rect 23032 21468 23060 21499
rect 23106 21496 23112 21548
rect 23164 21496 23170 21548
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 25041 21539 25099 21545
rect 25041 21505 25053 21539
rect 25087 21536 25099 21539
rect 25130 21536 25136 21548
rect 25087 21508 25136 21536
rect 25087 21505 25099 21508
rect 25041 21499 25099 21505
rect 22848 21440 23060 21468
rect 18932 21372 19656 21400
rect 18932 21360 18938 21372
rect 19702 21360 19708 21412
rect 19760 21360 19766 21412
rect 20162 21360 20168 21412
rect 20220 21360 20226 21412
rect 21082 21360 21088 21412
rect 21140 21360 21146 21412
rect 21913 21403 21971 21409
rect 21913 21369 21925 21403
rect 21959 21400 21971 21403
rect 22002 21400 22008 21412
rect 21959 21372 22008 21400
rect 21959 21369 21971 21372
rect 21913 21363 21971 21369
rect 22002 21360 22008 21372
rect 22060 21360 22066 21412
rect 23308 21400 23336 21499
rect 25130 21496 25136 21508
rect 25188 21496 25194 21548
rect 25222 21496 25228 21548
rect 25280 21496 25286 21548
rect 25314 21496 25320 21548
rect 25372 21536 25378 21548
rect 25685 21539 25743 21545
rect 25685 21536 25697 21539
rect 25372 21508 25697 21536
rect 25372 21496 25378 21508
rect 25685 21505 25697 21508
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 25774 21496 25780 21548
rect 25832 21536 25838 21548
rect 25869 21539 25927 21545
rect 25869 21536 25881 21539
rect 25832 21508 25881 21536
rect 25832 21496 25838 21508
rect 25869 21505 25881 21508
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 25958 21496 25964 21548
rect 26016 21496 26022 21548
rect 26053 21539 26111 21545
rect 26053 21505 26065 21539
rect 26099 21505 26111 21539
rect 26053 21499 26111 21505
rect 24857 21471 24915 21477
rect 24857 21437 24869 21471
rect 24903 21468 24915 21471
rect 25240 21468 25268 21496
rect 26068 21468 26096 21499
rect 26786 21496 26792 21548
rect 26844 21536 26850 21548
rect 27338 21536 27344 21548
rect 26844 21508 27344 21536
rect 26844 21496 26850 21508
rect 27338 21496 27344 21508
rect 27396 21496 27402 21548
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21505 27675 21539
rect 27617 21499 27675 21505
rect 24903 21440 25268 21468
rect 25792 21440 26096 21468
rect 24903 21437 24915 21440
rect 24857 21431 24915 21437
rect 25792 21409 25820 21440
rect 26970 21428 26976 21480
rect 27028 21468 27034 21480
rect 27632 21468 27660 21499
rect 27706 21496 27712 21548
rect 27764 21496 27770 21548
rect 27798 21468 27804 21480
rect 27028 21440 27804 21468
rect 27028 21428 27034 21440
rect 27798 21428 27804 21440
rect 27856 21468 27862 21480
rect 28442 21468 28448 21480
rect 27856 21440 28448 21468
rect 27856 21428 27862 21440
rect 28442 21428 28448 21440
rect 28500 21428 28506 21480
rect 22388 21372 23336 21400
rect 22388 21344 22416 21372
rect 17586 21332 17592 21344
rect 9876 21304 17592 21332
rect 17586 21292 17592 21304
rect 17644 21292 17650 21344
rect 17678 21292 17684 21344
rect 17736 21292 17742 21344
rect 17862 21292 17868 21344
rect 17920 21332 17926 21344
rect 22278 21332 22284 21344
rect 17920 21304 22284 21332
rect 17920 21292 17926 21304
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 22370 21292 22376 21344
rect 22428 21292 22434 21344
rect 22649 21335 22707 21341
rect 22649 21301 22661 21335
rect 22695 21332 22707 21335
rect 23014 21332 23020 21344
rect 22695 21304 23020 21332
rect 22695 21301 22707 21304
rect 22649 21295 22707 21301
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 23308 21332 23336 21372
rect 25777 21403 25835 21409
rect 25777 21369 25789 21403
rect 25823 21369 25835 21403
rect 28552 21400 28580 21576
rect 28718 21496 28724 21548
rect 28776 21536 28782 21548
rect 28997 21539 29055 21545
rect 28997 21536 29009 21539
rect 28776 21508 29009 21536
rect 28776 21496 28782 21508
rect 28997 21505 29009 21508
rect 29043 21505 29055 21539
rect 28997 21499 29055 21505
rect 29178 21496 29184 21548
rect 29236 21496 29242 21548
rect 29641 21539 29699 21545
rect 29641 21505 29653 21539
rect 29687 21536 29699 21539
rect 29748 21536 29776 21632
rect 32140 21604 32168 21632
rect 31680 21576 32168 21604
rect 32416 21604 32444 21632
rect 32416 21576 32996 21604
rect 30101 21542 30159 21545
rect 30190 21542 30196 21548
rect 30101 21539 30196 21542
rect 29687 21508 30052 21536
rect 29687 21505 29699 21508
rect 29641 21499 29699 21505
rect 29733 21471 29791 21477
rect 29733 21437 29745 21471
rect 29779 21468 29791 21471
rect 29914 21468 29920 21480
rect 29779 21440 29920 21468
rect 29779 21437 29791 21440
rect 29733 21431 29791 21437
rect 29914 21428 29920 21440
rect 29972 21428 29978 21480
rect 30024 21468 30052 21508
rect 30101 21505 30113 21539
rect 30147 21514 30196 21539
rect 30147 21505 30159 21514
rect 30101 21499 30159 21505
rect 30190 21496 30196 21514
rect 30248 21496 30254 21548
rect 30285 21539 30343 21545
rect 30285 21505 30297 21539
rect 30331 21505 30343 21539
rect 30285 21499 30343 21505
rect 30300 21468 30328 21499
rect 31478 21496 31484 21548
rect 31536 21536 31542 21548
rect 31680 21545 31708 21576
rect 31573 21539 31631 21545
rect 31573 21536 31585 21539
rect 31536 21508 31585 21536
rect 31536 21496 31542 21508
rect 31573 21505 31585 21508
rect 31619 21505 31631 21539
rect 31573 21499 31631 21505
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21505 31723 21539
rect 31665 21499 31723 21505
rect 31846 21496 31852 21548
rect 31904 21496 31910 21548
rect 32030 21496 32036 21548
rect 32088 21496 32094 21548
rect 32306 21496 32312 21548
rect 32364 21496 32370 21548
rect 32416 21545 32444 21576
rect 32401 21539 32459 21545
rect 32401 21505 32413 21539
rect 32447 21505 32459 21539
rect 32401 21499 32459 21505
rect 32582 21496 32588 21548
rect 32640 21496 32646 21548
rect 32766 21496 32772 21548
rect 32824 21496 32830 21548
rect 32968 21545 32996 21576
rect 32953 21539 33011 21545
rect 32953 21505 32965 21539
rect 32999 21505 33011 21539
rect 32953 21499 33011 21505
rect 33134 21496 33140 21548
rect 33192 21536 33198 21548
rect 33873 21539 33931 21545
rect 33873 21536 33885 21539
rect 33192 21508 33885 21536
rect 33192 21496 33198 21508
rect 30024 21440 30328 21468
rect 31757 21471 31815 21477
rect 31757 21437 31769 21471
rect 31803 21468 31815 21471
rect 32048 21468 32076 21496
rect 33336 21480 33364 21508
rect 33873 21505 33885 21508
rect 33919 21505 33931 21539
rect 33873 21499 33931 21505
rect 34054 21496 34060 21548
rect 34112 21496 34118 21548
rect 34164 21545 34192 21632
rect 34149 21539 34207 21545
rect 34149 21505 34161 21539
rect 34195 21505 34207 21539
rect 34149 21499 34207 21505
rect 34275 21539 34333 21545
rect 34275 21505 34287 21539
rect 34321 21536 34333 21539
rect 34698 21536 34704 21548
rect 34321 21508 34704 21536
rect 34321 21505 34333 21508
rect 34275 21499 34333 21505
rect 34698 21496 34704 21508
rect 34756 21496 34762 21548
rect 32493 21471 32551 21477
rect 32493 21468 32505 21471
rect 31803 21440 32505 21468
rect 31803 21437 31815 21440
rect 31757 21431 31815 21437
rect 32493 21437 32505 21440
rect 32539 21437 32551 21471
rect 32493 21431 32551 21437
rect 33318 21428 33324 21480
rect 33376 21428 33382 21480
rect 28552 21372 30328 21400
rect 25777 21363 25835 21369
rect 24946 21332 24952 21344
rect 23308 21304 24952 21332
rect 24946 21292 24952 21304
rect 25004 21292 25010 21344
rect 25222 21292 25228 21344
rect 25280 21292 25286 21344
rect 28997 21335 29055 21341
rect 28997 21301 29009 21335
rect 29043 21332 29055 21335
rect 29454 21332 29460 21344
rect 29043 21304 29460 21332
rect 29043 21301 29055 21304
rect 28997 21295 29055 21301
rect 29454 21292 29460 21304
rect 29512 21292 29518 21344
rect 29914 21292 29920 21344
rect 29972 21332 29978 21344
rect 30009 21335 30067 21341
rect 30009 21332 30021 21335
rect 29972 21304 30021 21332
rect 29972 21292 29978 21304
rect 30009 21301 30021 21304
rect 30055 21301 30067 21335
rect 30300 21332 30328 21372
rect 30466 21360 30472 21412
rect 30524 21400 30530 21412
rect 32125 21403 32183 21409
rect 32125 21400 32137 21403
rect 30524 21372 32137 21400
rect 30524 21360 30530 21372
rect 32125 21369 32137 21372
rect 32171 21369 32183 21403
rect 34517 21403 34575 21409
rect 34517 21400 34529 21403
rect 32125 21363 32183 21369
rect 33152 21372 34529 21400
rect 30926 21332 30932 21344
rect 30300 21304 30932 21332
rect 30009 21295 30067 21301
rect 30926 21292 30932 21304
rect 30984 21332 30990 21344
rect 33152 21332 33180 21372
rect 34517 21369 34529 21372
rect 34563 21369 34575 21403
rect 34517 21363 34575 21369
rect 30984 21304 33180 21332
rect 30984 21292 30990 21304
rect 1104 21242 38272 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38272 21242
rect 1104 21168 38272 21190
rect 1670 21128 1676 21140
rect 1412 21100 1676 21128
rect 1412 21001 1440 21100
rect 1670 21088 1676 21100
rect 1728 21088 1734 21140
rect 4157 21131 4215 21137
rect 4157 21097 4169 21131
rect 4203 21128 4215 21131
rect 4614 21128 4620 21140
rect 4203 21100 4620 21128
rect 4203 21097 4215 21100
rect 4157 21091 4215 21097
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20961 1455 20995
rect 1397 20955 1455 20961
rect 3142 20952 3148 21004
rect 3200 20992 3206 21004
rect 3789 20995 3847 21001
rect 3789 20992 3801 20995
rect 3200 20964 3801 20992
rect 3200 20952 3206 20964
rect 3789 20961 3801 20964
rect 3835 20992 3847 20995
rect 3878 20992 3884 21004
rect 3835 20964 3884 20992
rect 3835 20961 3847 20964
rect 3789 20955 3847 20961
rect 3878 20952 3884 20964
rect 3936 20992 3942 21004
rect 4062 20992 4068 21004
rect 3936 20964 4068 20992
rect 3936 20952 3942 20964
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 4264 20933 4292 21100
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 5534 21088 5540 21140
rect 5592 21088 5598 21140
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 9272 21100 10149 21128
rect 9272 21088 9278 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 10778 21088 10784 21140
rect 10836 21088 10842 21140
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 12805 21131 12863 21137
rect 12805 21128 12817 21131
rect 12492 21100 12817 21128
rect 12492 21088 12498 21100
rect 12805 21097 12817 21100
rect 12851 21097 12863 21131
rect 12805 21091 12863 21097
rect 14734 21088 14740 21140
rect 14792 21088 14798 21140
rect 16485 21131 16543 21137
rect 16485 21097 16497 21131
rect 16531 21128 16543 21131
rect 16574 21128 16580 21140
rect 16531 21100 16580 21128
rect 16531 21097 16543 21100
rect 16485 21091 16543 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 17310 21088 17316 21140
rect 17368 21088 17374 21140
rect 17494 21088 17500 21140
rect 17552 21128 17558 21140
rect 17589 21131 17647 21137
rect 17589 21128 17601 21131
rect 17552 21100 17601 21128
rect 17552 21088 17558 21100
rect 17589 21097 17601 21100
rect 17635 21097 17647 21131
rect 17589 21091 17647 21097
rect 17770 21088 17776 21140
rect 17828 21128 17834 21140
rect 18141 21131 18199 21137
rect 18141 21128 18153 21131
rect 17828 21100 18153 21128
rect 17828 21088 17834 21100
rect 18141 21097 18153 21100
rect 18187 21097 18199 21131
rect 18141 21091 18199 21097
rect 18248 21100 22692 21128
rect 5552 20992 5580 21088
rect 10318 21060 10324 21072
rect 5920 21032 10324 21060
rect 5552 20964 5764 20992
rect 3973 20927 4031 20933
rect 3973 20893 3985 20927
rect 4019 20893 4031 20927
rect 3973 20887 4031 20893
rect 4249 20927 4307 20933
rect 4249 20893 4261 20927
rect 4295 20893 4307 20927
rect 4249 20887 4307 20893
rect 5537 20927 5595 20933
rect 5537 20893 5549 20927
rect 5583 20893 5595 20927
rect 5537 20887 5595 20893
rect 1670 20816 1676 20868
rect 1728 20816 1734 20868
rect 3234 20856 3240 20868
rect 2898 20828 3240 20856
rect 3234 20816 3240 20828
rect 3292 20816 3298 20868
rect 3988 20856 4016 20887
rect 4154 20856 4160 20868
rect 3988 20828 4160 20856
rect 4154 20816 4160 20828
rect 4212 20856 4218 20868
rect 5552 20856 5580 20887
rect 5626 20884 5632 20936
rect 5684 20884 5690 20936
rect 5736 20933 5764 20964
rect 5920 20933 5948 21032
rect 10318 21020 10324 21032
rect 10376 21020 10382 21072
rect 17862 21060 17868 21072
rect 12544 21032 17868 21060
rect 9968 20964 10640 20992
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20893 5779 20927
rect 5721 20887 5779 20893
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20893 5963 20927
rect 5905 20887 5963 20893
rect 9122 20884 9128 20936
rect 9180 20924 9186 20936
rect 9585 20927 9643 20933
rect 9585 20924 9597 20927
rect 9180 20896 9597 20924
rect 9180 20884 9186 20896
rect 9585 20893 9597 20896
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 9968 20933 9996 20964
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20893 10011 20927
rect 9953 20887 10011 20893
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20924 10287 20927
rect 10318 20924 10324 20936
rect 10275 20896 10324 20924
rect 10275 20893 10287 20896
rect 10229 20887 10287 20893
rect 10318 20884 10324 20896
rect 10376 20884 10382 20936
rect 10410 20884 10416 20936
rect 10468 20884 10474 20936
rect 10612 20933 10640 20964
rect 10597 20927 10655 20933
rect 10597 20893 10609 20927
rect 10643 20924 10655 20927
rect 10686 20924 10692 20936
rect 10643 20896 10692 20924
rect 10643 20893 10655 20896
rect 10597 20887 10655 20893
rect 10686 20884 10692 20896
rect 10744 20884 10750 20936
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 12250 20924 12256 20936
rect 11204 20896 12256 20924
rect 11204 20884 11210 20896
rect 12250 20884 12256 20896
rect 12308 20884 12314 20936
rect 12544 20933 12572 21032
rect 17862 21020 17868 21032
rect 17920 21020 17926 21072
rect 14458 20992 14464 21004
rect 14108 20964 14464 20992
rect 12710 20933 12716 20936
rect 12529 20927 12587 20933
rect 12529 20893 12541 20927
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 12673 20927 12716 20933
rect 12673 20893 12685 20927
rect 12768 20924 12774 20936
rect 13354 20924 13360 20936
rect 12768 20896 13360 20924
rect 12673 20887 12716 20893
rect 12710 20884 12716 20887
rect 12768 20884 12774 20896
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 14108 20933 14136 20964
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 15304 20964 17448 20992
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14241 20927 14299 20933
rect 14241 20893 14253 20927
rect 14287 20924 14299 20927
rect 14369 20927 14427 20933
rect 14287 20893 14320 20924
rect 14241 20887 14320 20893
rect 14369 20893 14381 20927
rect 14415 20893 14427 20927
rect 14369 20887 14427 20893
rect 14599 20927 14657 20933
rect 14599 20893 14611 20927
rect 14645 20924 14657 20927
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 14645 20896 14933 20924
rect 14645 20893 14657 20896
rect 14599 20887 14657 20893
rect 14921 20893 14933 20896
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 9398 20856 9404 20868
rect 4212 20828 4476 20856
rect 5552 20828 9404 20856
rect 4212 20816 4218 20828
rect 4448 20800 4476 20828
rect 9398 20816 9404 20828
rect 9456 20816 9462 20868
rect 9858 20816 9864 20868
rect 9916 20816 9922 20868
rect 10134 20816 10140 20868
rect 10192 20856 10198 20868
rect 10505 20859 10563 20865
rect 10505 20856 10517 20859
rect 10192 20828 10517 20856
rect 10192 20816 10198 20828
rect 10505 20825 10517 20828
rect 10551 20825 10563 20859
rect 10505 20819 10563 20825
rect 12158 20816 12164 20868
rect 12216 20856 12222 20868
rect 12437 20859 12495 20865
rect 12437 20856 12449 20859
rect 12216 20828 12449 20856
rect 12216 20816 12222 20828
rect 12437 20825 12449 20828
rect 12483 20825 12495 20859
rect 12437 20819 12495 20825
rect 3694 20748 3700 20800
rect 3752 20788 3758 20800
rect 4341 20791 4399 20797
rect 4341 20788 4353 20791
rect 3752 20760 4353 20788
rect 3752 20748 3758 20760
rect 4341 20757 4353 20760
rect 4387 20757 4399 20791
rect 4341 20751 4399 20757
rect 4430 20748 4436 20800
rect 4488 20748 4494 20800
rect 5258 20748 5264 20800
rect 5316 20748 5322 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 9950 20788 9956 20800
rect 9732 20760 9956 20788
rect 9732 20748 9738 20760
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 10410 20748 10416 20800
rect 10468 20788 10474 20800
rect 12176 20788 12204 20816
rect 10468 20760 12204 20788
rect 10468 20748 10474 20760
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14292 20788 14320 20887
rect 14384 20800 14412 20887
rect 15010 20884 15016 20936
rect 15068 20924 15074 20936
rect 15105 20927 15163 20933
rect 15105 20924 15117 20927
rect 15068 20896 15117 20924
rect 15068 20884 15074 20896
rect 15105 20893 15117 20896
rect 15151 20893 15163 20927
rect 15105 20887 15163 20893
rect 14461 20859 14519 20865
rect 14461 20825 14473 20859
rect 14507 20856 14519 20859
rect 14734 20856 14740 20868
rect 14507 20828 14740 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 14734 20816 14740 20828
rect 14792 20816 14798 20868
rect 13872 20760 14320 20788
rect 13872 20748 13878 20760
rect 14366 20748 14372 20800
rect 14424 20748 14430 20800
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15304 20797 15332 20964
rect 15381 20927 15439 20933
rect 15381 20893 15393 20927
rect 15427 20924 15439 20927
rect 15427 20896 15700 20924
rect 15427 20893 15439 20896
rect 15381 20887 15439 20893
rect 15672 20800 15700 20896
rect 16298 20884 16304 20936
rect 16356 20884 16362 20936
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 17420 20933 17448 20964
rect 17586 20952 17592 21004
rect 17644 20992 17650 21004
rect 18248 20992 18276 21100
rect 18874 21020 18880 21072
rect 18932 21060 18938 21072
rect 18932 21032 19656 21060
rect 18932 21020 18938 21032
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 17644 20964 18276 20992
rect 18340 20964 19257 20992
rect 17644 20952 17650 20964
rect 18340 20936 18368 20964
rect 19245 20961 19257 20964
rect 19291 20961 19303 20995
rect 19245 20955 19303 20961
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 19521 20995 19579 21001
rect 19521 20992 19533 20995
rect 19484 20964 19533 20992
rect 19484 20952 19490 20964
rect 19521 20961 19533 20964
rect 19567 20961 19579 20995
rect 19628 20992 19656 21032
rect 21910 21020 21916 21072
rect 21968 21060 21974 21072
rect 22005 21063 22063 21069
rect 22005 21060 22017 21063
rect 21968 21032 22017 21060
rect 21968 21020 21974 21032
rect 22005 21029 22017 21032
rect 22051 21029 22063 21063
rect 22005 21023 22063 21029
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19628 20964 19993 20992
rect 19521 20955 19579 20961
rect 19981 20961 19993 20964
rect 20027 20961 20039 20995
rect 19981 20955 20039 20961
rect 20162 20952 20168 21004
rect 20220 20992 20226 21004
rect 22370 20992 22376 21004
rect 20220 20964 22376 20992
rect 20220 20952 20226 20964
rect 22370 20952 22376 20964
rect 22428 20952 22434 21004
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 16540 20896 16773 20924
rect 16540 20884 16546 20896
rect 16761 20893 16773 20896
rect 16807 20893 16819 20927
rect 16761 20887 16819 20893
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20893 17279 20927
rect 17221 20887 17279 20893
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20893 17463 20927
rect 17770 20924 17776 20936
rect 17731 20896 17776 20924
rect 17405 20887 17463 20893
rect 15746 20816 15752 20868
rect 15804 20856 15810 20868
rect 16500 20856 16528 20884
rect 15804 20828 16528 20856
rect 15804 20816 15810 20828
rect 16574 20816 16580 20868
rect 16632 20856 16638 20868
rect 17236 20856 17264 20887
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 18012 20896 18245 20924
rect 18012 20884 18018 20896
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 18248 20856 18276 20887
rect 18322 20884 18328 20936
rect 18380 20884 18386 20936
rect 18874 20933 18880 20936
rect 18418 20927 18476 20933
rect 18418 20893 18430 20927
rect 18464 20893 18476 20927
rect 18418 20887 18476 20893
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 18831 20927 18880 20933
rect 18831 20893 18843 20927
rect 18877 20893 18880 20927
rect 18831 20887 18880 20893
rect 18432 20856 18460 20887
rect 16632 20828 17264 20856
rect 17328 20828 18184 20856
rect 18248 20828 18460 20856
rect 16632 20816 16638 20828
rect 15289 20791 15347 20797
rect 15289 20788 15301 20791
rect 15252 20760 15301 20788
rect 15252 20748 15258 20760
rect 15289 20757 15301 20760
rect 15335 20757 15347 20791
rect 15289 20751 15347 20757
rect 15654 20748 15660 20800
rect 15712 20748 15718 20800
rect 16022 20748 16028 20800
rect 16080 20788 16086 20800
rect 16669 20791 16727 20797
rect 16669 20788 16681 20791
rect 16080 20760 16681 20788
rect 16080 20748 16086 20760
rect 16669 20757 16681 20760
rect 16715 20788 16727 20791
rect 17328 20788 17356 20828
rect 16715 20760 17356 20788
rect 16715 20757 16727 20760
rect 16669 20751 16727 20757
rect 17678 20748 17684 20800
rect 17736 20788 17742 20800
rect 17773 20791 17831 20797
rect 17773 20788 17785 20791
rect 17736 20760 17785 20788
rect 17736 20748 17742 20760
rect 17773 20757 17785 20760
rect 17819 20757 17831 20791
rect 18156 20788 18184 20828
rect 18598 20816 18604 20868
rect 18656 20816 18662 20868
rect 18708 20856 18736 20887
rect 18874 20884 18880 20887
rect 18932 20884 18938 20936
rect 19058 20884 19064 20936
rect 19116 20924 19122 20936
rect 19705 20927 19763 20933
rect 19705 20926 19717 20927
rect 19536 20924 19717 20926
rect 19116 20898 19717 20924
rect 19116 20896 19564 20898
rect 19116 20884 19122 20896
rect 19705 20893 19717 20898
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 20073 20927 20131 20933
rect 20073 20893 20085 20927
rect 20119 20893 20131 20927
rect 20073 20887 20131 20893
rect 18708 20828 19380 20856
rect 18708 20788 18736 20828
rect 18156 20760 18736 20788
rect 17773 20751 17831 20757
rect 18966 20748 18972 20800
rect 19024 20748 19030 20800
rect 19352 20788 19380 20828
rect 19426 20816 19432 20868
rect 19484 20816 19490 20868
rect 19702 20788 19708 20800
rect 19352 20760 19708 20788
rect 19702 20748 19708 20760
rect 19760 20788 19766 20800
rect 20088 20788 20116 20887
rect 20714 20884 20720 20936
rect 20772 20884 20778 20936
rect 20806 20884 20812 20936
rect 20864 20884 20870 20936
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20893 21051 20927
rect 20993 20887 21051 20893
rect 20732 20856 20760 20884
rect 21008 20856 21036 20887
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 21361 20927 21419 20933
rect 21361 20924 21373 20927
rect 21140 20896 21373 20924
rect 21140 20884 21146 20896
rect 21361 20893 21373 20896
rect 21407 20893 21419 20927
rect 21361 20887 21419 20893
rect 21450 20884 21456 20936
rect 21508 20924 21514 20936
rect 21729 20927 21787 20933
rect 21729 20924 21741 20927
rect 21508 20896 21741 20924
rect 21508 20884 21514 20896
rect 21729 20893 21741 20896
rect 21775 20893 21787 20927
rect 22664 20924 22692 21100
rect 23750 21088 23756 21140
rect 23808 21088 23814 21140
rect 26878 21128 26884 21140
rect 23952 21100 26884 21128
rect 23952 21001 23980 21100
rect 26878 21088 26884 21100
rect 26936 21128 26942 21140
rect 26936 21100 27016 21128
rect 26936 21088 26942 21100
rect 26988 21060 27016 21100
rect 27154 21088 27160 21140
rect 27212 21128 27218 21140
rect 27249 21131 27307 21137
rect 27249 21128 27261 21131
rect 27212 21100 27261 21128
rect 27212 21088 27218 21100
rect 27249 21097 27261 21100
rect 27295 21097 27307 21131
rect 27249 21091 27307 21097
rect 27614 21088 27620 21140
rect 27672 21128 27678 21140
rect 34701 21131 34759 21137
rect 27672 21100 31754 21128
rect 27672 21088 27678 21100
rect 28350 21060 28356 21072
rect 24044 21032 26924 21060
rect 26988 21032 28356 21060
rect 23937 20995 23995 21001
rect 23937 20961 23949 20995
rect 23983 20961 23995 20995
rect 23937 20955 23995 20961
rect 24044 20933 24072 21032
rect 24118 20952 24124 21004
rect 24176 20952 24182 21004
rect 24412 20964 24992 20992
rect 24029 20927 24087 20933
rect 24029 20924 24041 20927
rect 22664 20896 24041 20924
rect 21729 20887 21787 20893
rect 24029 20893 24041 20896
rect 24075 20893 24087 20927
rect 24136 20924 24164 20952
rect 24412 20933 24440 20964
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 24136 20896 24409 20924
rect 24029 20887 24087 20893
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 24486 20884 24492 20936
rect 24544 20924 24550 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24544 20896 24777 20924
rect 24544 20884 24550 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 20732 20828 21036 20856
rect 23753 20859 23811 20865
rect 23753 20825 23765 20859
rect 23799 20856 23811 20859
rect 24118 20856 24124 20868
rect 23799 20828 24124 20856
rect 23799 20825 23811 20828
rect 23753 20819 23811 20825
rect 24118 20816 24124 20828
rect 24176 20856 24182 20868
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 24176 20828 24593 20856
rect 24176 20816 24182 20828
rect 24581 20825 24593 20828
rect 24627 20825 24639 20859
rect 24581 20819 24639 20825
rect 24673 20859 24731 20865
rect 24673 20825 24685 20859
rect 24719 20856 24731 20859
rect 24854 20856 24860 20868
rect 24719 20828 24860 20856
rect 24719 20825 24731 20828
rect 24673 20819 24731 20825
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 24964 20856 24992 20964
rect 25038 20952 25044 21004
rect 25096 20952 25102 21004
rect 25130 20952 25136 21004
rect 25188 20952 25194 21004
rect 25406 20952 25412 21004
rect 25464 20952 25470 21004
rect 26896 20992 26924 21032
rect 28350 21020 28356 21032
rect 28408 21060 28414 21072
rect 31726 21060 31754 21100
rect 34701 21097 34713 21131
rect 34747 21128 34759 21131
rect 34790 21128 34796 21140
rect 34747 21100 34796 21128
rect 34747 21097 34759 21100
rect 34701 21091 34759 21097
rect 34790 21088 34796 21100
rect 34848 21088 34854 21140
rect 28408 21032 30696 21060
rect 31726 21032 37412 21060
rect 28408 21020 28414 21032
rect 30193 20995 30251 21001
rect 30193 20992 30205 20995
rect 26896 20964 30205 20992
rect 25148 20924 25176 20952
rect 25225 20927 25283 20933
rect 25225 20924 25237 20927
rect 25148 20896 25237 20924
rect 25225 20893 25237 20896
rect 25271 20893 25283 20927
rect 26697 20927 26755 20933
rect 26697 20924 26709 20927
rect 25225 20887 25283 20893
rect 26068 20896 26709 20924
rect 26068 20868 26096 20896
rect 26697 20893 26709 20896
rect 26743 20924 26755 20927
rect 26786 20924 26792 20936
rect 26743 20896 26792 20924
rect 26743 20893 26755 20896
rect 26697 20887 26755 20893
rect 26786 20884 26792 20896
rect 26844 20884 26850 20936
rect 26896 20933 26924 20964
rect 30193 20961 30205 20964
rect 30239 20961 30251 20995
rect 30193 20955 30251 20961
rect 26881 20927 26939 20933
rect 26881 20893 26893 20927
rect 26927 20893 26939 20927
rect 26881 20887 26939 20893
rect 27065 20927 27123 20933
rect 27065 20893 27077 20927
rect 27111 20924 27123 20927
rect 27154 20924 27160 20936
rect 27111 20896 27160 20924
rect 27111 20893 27123 20896
rect 27065 20887 27123 20893
rect 27154 20884 27160 20896
rect 27212 20884 27218 20936
rect 27246 20884 27252 20936
rect 27304 20884 27310 20936
rect 29822 20884 29828 20936
rect 29880 20884 29886 20936
rect 29914 20884 29920 20936
rect 29972 20924 29978 20936
rect 30009 20927 30067 20933
rect 30009 20924 30021 20927
rect 29972 20896 30021 20924
rect 29972 20884 29978 20896
rect 30009 20893 30021 20896
rect 30055 20893 30067 20927
rect 30009 20887 30067 20893
rect 26050 20856 26056 20868
rect 24964 20828 26056 20856
rect 26050 20816 26056 20828
rect 26108 20816 26114 20868
rect 26326 20816 26332 20868
rect 26384 20856 26390 20868
rect 26970 20856 26976 20868
rect 26384 20828 26976 20856
rect 26384 20816 26390 20828
rect 26970 20816 26976 20828
rect 27028 20816 27034 20868
rect 20162 20788 20168 20800
rect 19760 20760 20168 20788
rect 19760 20748 19766 20760
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 24210 20748 24216 20800
rect 24268 20748 24274 20800
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 27264 20788 27292 20884
rect 24995 20760 27292 20788
rect 30024 20788 30052 20887
rect 30668 20856 30696 21032
rect 32401 20995 32459 21001
rect 32401 20961 32413 20995
rect 32447 20992 32459 20995
rect 32490 20992 32496 21004
rect 32447 20964 32496 20992
rect 32447 20961 32459 20964
rect 32401 20955 32459 20961
rect 31294 20884 31300 20936
rect 31352 20924 31358 20936
rect 32309 20927 32367 20933
rect 32309 20924 32321 20927
rect 31352 20896 32321 20924
rect 31352 20884 31358 20896
rect 32309 20893 32321 20896
rect 32355 20893 32367 20927
rect 32309 20887 32367 20893
rect 32416 20856 32444 20955
rect 32490 20952 32496 20964
rect 32548 20952 32554 21004
rect 34698 20952 34704 21004
rect 34756 20992 34762 21004
rect 34977 20995 35035 21001
rect 34977 20992 34989 20995
rect 34756 20964 34989 20992
rect 34756 20952 34762 20964
rect 34977 20961 34989 20964
rect 35023 20961 35035 20995
rect 34977 20955 35035 20961
rect 35069 20995 35127 21001
rect 35069 20961 35081 20995
rect 35115 20992 35127 20995
rect 35621 20995 35679 21001
rect 35621 20992 35633 20995
rect 35115 20964 35633 20992
rect 35115 20961 35127 20964
rect 35069 20955 35127 20961
rect 35621 20961 35633 20964
rect 35667 20961 35679 20995
rect 35621 20955 35679 20961
rect 35894 20952 35900 21004
rect 35952 20952 35958 21004
rect 34514 20884 34520 20936
rect 34572 20924 34578 20936
rect 34885 20927 34943 20933
rect 34885 20924 34897 20927
rect 34572 20896 34897 20924
rect 34572 20884 34578 20896
rect 34885 20893 34897 20896
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 35158 20884 35164 20936
rect 35216 20884 35222 20936
rect 35529 20927 35587 20933
rect 35529 20893 35541 20927
rect 35575 20924 35587 20927
rect 35912 20924 35940 20952
rect 37384 20933 37412 21032
rect 35575 20896 35940 20924
rect 37369 20927 37427 20933
rect 35575 20893 35587 20896
rect 35529 20887 35587 20893
rect 37369 20893 37381 20927
rect 37415 20893 37427 20927
rect 37369 20887 37427 20893
rect 37553 20859 37611 20865
rect 37553 20856 37565 20859
rect 30668 20828 32444 20856
rect 37200 20828 37565 20856
rect 31110 20788 31116 20800
rect 30024 20760 31116 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 31110 20748 31116 20760
rect 31168 20748 31174 20800
rect 32677 20791 32735 20797
rect 32677 20757 32689 20791
rect 32723 20788 32735 20791
rect 33042 20788 33048 20800
rect 32723 20760 33048 20788
rect 32723 20757 32735 20760
rect 32677 20751 32735 20757
rect 33042 20748 33048 20760
rect 33100 20748 33106 20800
rect 37200 20797 37228 20828
rect 37553 20825 37565 20828
rect 37599 20825 37611 20859
rect 37553 20819 37611 20825
rect 37185 20791 37243 20797
rect 37185 20757 37197 20791
rect 37231 20757 37243 20791
rect 37185 20751 37243 20757
rect 37829 20791 37887 20797
rect 37829 20757 37841 20791
rect 37875 20788 37887 20791
rect 37875 20760 38424 20788
rect 37875 20757 37887 20760
rect 37829 20751 37887 20757
rect 38396 20732 38424 20760
rect 1104 20698 38272 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38272 20698
rect 38378 20680 38384 20732
rect 38436 20680 38442 20732
rect 1104 20624 38272 20646
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 992 20556 1593 20584
rect 992 20544 998 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 1670 20544 1676 20596
rect 1728 20584 1734 20596
rect 2317 20587 2375 20593
rect 2317 20584 2329 20587
rect 1728 20556 2329 20584
rect 1728 20544 1734 20556
rect 2317 20553 2329 20556
rect 2363 20553 2375 20587
rect 2317 20547 2375 20553
rect 2498 20544 2504 20596
rect 2556 20544 2562 20596
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 3421 20587 3479 20593
rect 3421 20584 3433 20587
rect 3016 20556 3433 20584
rect 3016 20544 3022 20556
rect 3421 20553 3433 20556
rect 3467 20553 3479 20587
rect 3421 20547 3479 20553
rect 3602 20544 3608 20596
rect 3660 20544 3666 20596
rect 4890 20584 4896 20596
rect 4080 20556 4896 20584
rect 1489 20519 1547 20525
rect 1489 20485 1501 20519
rect 1535 20516 1547 20519
rect 1762 20516 1768 20528
rect 1535 20488 1768 20516
rect 1535 20485 1547 20488
rect 1489 20479 1547 20485
rect 1762 20476 1768 20488
rect 1820 20476 1826 20528
rect 2222 20408 2228 20460
rect 2280 20408 2286 20460
rect 2516 20457 2544 20544
rect 3620 20516 3648 20544
rect 3789 20519 3847 20525
rect 3789 20516 3801 20519
rect 3620 20488 3801 20516
rect 3789 20485 3801 20488
rect 3835 20485 3847 20519
rect 3789 20479 3847 20485
rect 3927 20519 3985 20525
rect 3927 20485 3939 20519
rect 3973 20516 3985 20519
rect 4080 20516 4108 20556
rect 4890 20544 4896 20556
rect 4948 20544 4954 20596
rect 8570 20544 8576 20596
rect 8628 20544 8634 20596
rect 9490 20544 9496 20596
rect 9548 20584 9554 20596
rect 9585 20587 9643 20593
rect 9585 20584 9597 20587
rect 9548 20556 9597 20584
rect 9548 20544 9554 20556
rect 9585 20553 9597 20556
rect 9631 20553 9643 20587
rect 10502 20584 10508 20596
rect 9585 20547 9643 20553
rect 9692 20556 10508 20584
rect 4430 20516 4436 20528
rect 3973 20488 4108 20516
rect 4172 20488 4436 20516
rect 3973 20485 3985 20488
rect 3927 20479 3985 20485
rect 2501 20451 2559 20457
rect 2501 20417 2513 20451
rect 2547 20417 2559 20451
rect 2501 20411 2559 20417
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 1486 20204 1492 20256
rect 1544 20244 1550 20256
rect 2041 20247 2099 20253
rect 2041 20244 2053 20247
rect 1544 20216 2053 20244
rect 1544 20204 1550 20216
rect 2041 20213 2053 20216
rect 2087 20213 2099 20247
rect 2700 20244 2728 20411
rect 3234 20340 3240 20392
rect 3292 20340 3298 20392
rect 3620 20312 3648 20411
rect 3694 20408 3700 20460
rect 3752 20408 3758 20460
rect 4062 20408 4068 20460
rect 4120 20408 4126 20460
rect 4172 20457 4200 20488
rect 4430 20476 4436 20488
rect 4488 20516 4494 20528
rect 4488 20488 4936 20516
rect 4488 20476 4494 20488
rect 4908 20460 4936 20488
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20417 4215 20451
rect 4157 20411 4215 20417
rect 4246 20408 4252 20460
rect 4304 20448 4310 20460
rect 4341 20451 4399 20457
rect 4341 20448 4353 20451
rect 4304 20420 4353 20448
rect 4304 20408 4310 20420
rect 4341 20417 4353 20420
rect 4387 20417 4399 20451
rect 4341 20411 4399 20417
rect 4890 20408 4896 20460
rect 4948 20408 4954 20460
rect 8234 20420 8340 20448
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 6871 20352 6960 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 4525 20315 4583 20321
rect 4525 20312 4537 20315
rect 3620 20284 4537 20312
rect 4525 20281 4537 20284
rect 4571 20281 4583 20315
rect 4525 20275 4583 20281
rect 6932 20256 6960 20352
rect 7098 20340 7104 20392
rect 7156 20340 7162 20392
rect 8312 20256 8340 20420
rect 9030 20408 9036 20460
rect 9088 20408 9094 20460
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 9232 20312 9260 20411
rect 9306 20408 9312 20460
rect 9364 20408 9370 20460
rect 9692 20457 9720 20556
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 10870 20544 10876 20596
rect 10928 20544 10934 20596
rect 11882 20544 11888 20596
rect 11940 20544 11946 20596
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 14182 20584 14188 20596
rect 12023 20556 14188 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 9766 20476 9772 20528
rect 9824 20516 9830 20528
rect 9861 20519 9919 20525
rect 9861 20516 9873 20519
rect 9824 20488 9873 20516
rect 9824 20476 9830 20488
rect 9861 20485 9873 20488
rect 9907 20485 9919 20519
rect 9861 20479 9919 20485
rect 10226 20476 10232 20528
rect 10284 20516 10290 20528
rect 10284 20488 10640 20516
rect 10284 20476 10290 20488
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20417 9459 20451
rect 9401 20411 9459 20417
rect 9677 20451 9735 20457
rect 9677 20417 9689 20451
rect 9723 20417 9735 20451
rect 9677 20411 9735 20417
rect 9416 20380 9444 20411
rect 9950 20408 9956 20460
rect 10008 20408 10014 20460
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10060 20380 10088 20411
rect 10318 20408 10324 20460
rect 10376 20408 10382 20460
rect 10410 20408 10416 20460
rect 10468 20448 10474 20460
rect 10612 20457 10640 20488
rect 10888 20488 12756 20516
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10468 20420 10517 20448
rect 10468 20408 10474 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 10597 20451 10655 20457
rect 10597 20417 10609 20451
rect 10643 20417 10655 20451
rect 10597 20411 10655 20417
rect 10686 20408 10692 20460
rect 10744 20448 10750 20460
rect 10888 20448 10916 20488
rect 12728 20460 12756 20488
rect 10744 20420 10916 20448
rect 10744 20408 10750 20420
rect 11790 20408 11796 20460
rect 11848 20408 11854 20460
rect 12158 20408 12164 20460
rect 12216 20408 12222 20460
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 10704 20380 10732 20408
rect 9416 20352 10732 20380
rect 12636 20380 12664 20411
rect 12710 20408 12716 20460
rect 12768 20408 12774 20460
rect 12820 20380 12848 20556
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 14274 20544 14280 20596
rect 14332 20584 14338 20596
rect 14461 20587 14519 20593
rect 14461 20584 14473 20587
rect 14332 20556 14473 20584
rect 14332 20544 14338 20556
rect 14461 20553 14473 20556
rect 14507 20553 14519 20587
rect 14461 20547 14519 20553
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 14792 20556 15056 20584
rect 14792 20544 14798 20556
rect 15028 20525 15056 20556
rect 15102 20544 15108 20596
rect 15160 20584 15166 20596
rect 15289 20587 15347 20593
rect 15289 20584 15301 20587
rect 15160 20556 15301 20584
rect 15160 20544 15166 20556
rect 15289 20553 15301 20556
rect 15335 20553 15347 20587
rect 16758 20584 16764 20596
rect 15289 20547 15347 20553
rect 15488 20556 16764 20584
rect 14921 20519 14979 20525
rect 14921 20516 14933 20519
rect 14384 20488 14933 20516
rect 14384 20460 14412 20488
rect 14921 20485 14933 20488
rect 14967 20485 14979 20519
rect 14921 20479 14979 20485
rect 15013 20519 15071 20525
rect 15013 20485 15025 20519
rect 15059 20516 15071 20519
rect 15488 20516 15516 20556
rect 16758 20544 16764 20556
rect 16816 20584 16822 20596
rect 16816 20556 20300 20584
rect 16816 20544 16822 20556
rect 15059 20488 15516 20516
rect 15059 20485 15071 20488
rect 15013 20479 15071 20485
rect 16574 20476 16580 20528
rect 16632 20516 16638 20528
rect 16853 20519 16911 20525
rect 16853 20516 16865 20519
rect 16632 20488 16865 20516
rect 16632 20476 16638 20488
rect 16853 20485 16865 20488
rect 16899 20485 16911 20519
rect 16853 20479 16911 20485
rect 17310 20476 17316 20528
rect 17368 20516 17374 20528
rect 17678 20516 17684 20528
rect 17368 20488 17684 20516
rect 17368 20476 17374 20488
rect 17678 20476 17684 20488
rect 17736 20476 17742 20528
rect 18322 20476 18328 20528
rect 18380 20476 18386 20528
rect 18598 20476 18604 20528
rect 18656 20516 18662 20528
rect 19058 20516 19064 20528
rect 18656 20488 19064 20516
rect 18656 20476 18662 20488
rect 19058 20476 19064 20488
rect 19116 20476 19122 20528
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 13722 20448 13728 20460
rect 12943 20420 13728 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 12636 20352 12848 20380
rect 10229 20315 10287 20321
rect 9232 20284 9674 20312
rect 5810 20244 5816 20256
rect 2700 20216 5816 20244
rect 2041 20207 2099 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 6914 20204 6920 20256
rect 6972 20204 6978 20256
rect 8294 20204 8300 20256
rect 8352 20204 8358 20256
rect 9646 20244 9674 20284
rect 10229 20281 10241 20315
rect 10275 20312 10287 20315
rect 11238 20312 11244 20324
rect 10275 20284 11244 20312
rect 10275 20281 10287 20284
rect 10229 20275 10287 20281
rect 11238 20272 11244 20284
rect 11296 20272 11302 20324
rect 11609 20315 11667 20321
rect 11609 20281 11621 20315
rect 11655 20312 11667 20315
rect 12912 20312 12940 20411
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 13965 20451 14023 20457
rect 13965 20417 13977 20451
rect 14011 20448 14023 20451
rect 14011 20417 14044 20448
rect 13965 20411 14044 20417
rect 13832 20380 13860 20411
rect 13832 20352 13946 20380
rect 11655 20284 12940 20312
rect 11655 20281 11667 20284
rect 11609 20275 11667 20281
rect 9766 20244 9772 20256
rect 9646 20216 9772 20244
rect 9766 20204 9772 20216
rect 9824 20244 9830 20256
rect 10410 20244 10416 20256
rect 9824 20216 10416 20244
rect 9824 20204 9830 20216
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 12360 20244 12388 20284
rect 12434 20244 12440 20256
rect 12360 20216 12440 20244
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 13918 20244 13946 20352
rect 14016 20312 14044 20411
rect 14090 20408 14096 20460
rect 14148 20408 14154 20460
rect 14366 20457 14372 20460
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 14323 20451 14372 20457
rect 14323 20417 14335 20451
rect 14369 20417 14372 20451
rect 14323 20411 14372 20417
rect 14200 20380 14228 20411
rect 14366 20408 14372 20411
rect 14424 20448 14430 20460
rect 14424 20420 14471 20448
rect 14424 20408 14430 20420
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 14645 20451 14703 20457
rect 14645 20448 14657 20451
rect 14608 20420 14657 20448
rect 14608 20408 14614 20420
rect 14645 20417 14657 20420
rect 14691 20417 14703 20451
rect 14645 20411 14703 20417
rect 14793 20451 14851 20457
rect 14793 20417 14805 20451
rect 14839 20448 14851 20451
rect 14839 20420 15056 20448
rect 14839 20417 14851 20420
rect 14793 20411 14851 20417
rect 14458 20380 14464 20392
rect 14200 20352 14464 20380
rect 14458 20340 14464 20352
rect 14516 20380 14522 20392
rect 15028 20380 15056 20420
rect 15102 20408 15108 20460
rect 15160 20457 15166 20460
rect 15160 20448 15168 20457
rect 15160 20420 15205 20448
rect 15160 20411 15168 20420
rect 15160 20408 15166 20411
rect 15470 20408 15476 20460
rect 15528 20408 15534 20460
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 15712 20420 16681 20448
rect 15712 20408 15718 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 17218 20448 17224 20460
rect 16669 20411 16727 20417
rect 16776 20420 17224 20448
rect 15488 20380 15516 20408
rect 16776 20380 16804 20420
rect 17218 20408 17224 20420
rect 17276 20448 17282 20460
rect 18340 20448 18368 20476
rect 20272 20460 20300 20556
rect 24118 20544 24124 20596
rect 24176 20584 24182 20596
rect 24213 20587 24271 20593
rect 24213 20584 24225 20587
rect 24176 20556 24225 20584
rect 24176 20544 24182 20556
rect 24213 20553 24225 20556
rect 24259 20553 24271 20587
rect 33962 20584 33968 20596
rect 24213 20547 24271 20553
rect 24964 20556 33968 20584
rect 22925 20519 22983 20525
rect 22925 20485 22937 20519
rect 22971 20516 22983 20519
rect 23658 20516 23664 20528
rect 22971 20488 23664 20516
rect 22971 20485 22983 20488
rect 22925 20479 22983 20485
rect 23658 20476 23664 20488
rect 23716 20476 23722 20528
rect 17276 20420 18368 20448
rect 17276 20408 17282 20420
rect 17696 20392 17724 20420
rect 20070 20408 20076 20460
rect 20128 20408 20134 20460
rect 20254 20408 20260 20460
rect 20312 20408 20318 20460
rect 20346 20408 20352 20460
rect 20404 20408 20410 20460
rect 20714 20408 20720 20460
rect 20772 20408 20778 20460
rect 20806 20408 20812 20460
rect 20864 20408 20870 20460
rect 21266 20408 21272 20460
rect 21324 20408 21330 20460
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 23014 20448 23020 20460
rect 22336 20420 23020 20448
rect 22336 20408 22342 20420
rect 23014 20408 23020 20420
rect 23072 20448 23078 20460
rect 23201 20451 23259 20457
rect 23201 20448 23213 20451
rect 23072 20420 23213 20448
rect 23072 20408 23078 20420
rect 23201 20417 23213 20420
rect 23247 20417 23259 20451
rect 23201 20411 23259 20417
rect 23934 20408 23940 20460
rect 23992 20448 23998 20460
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 23992 20420 24133 20448
rect 23992 20408 23998 20420
rect 24121 20417 24133 20420
rect 24167 20448 24179 20451
rect 24964 20448 24992 20556
rect 33962 20544 33968 20556
rect 34020 20584 34026 20596
rect 35713 20587 35771 20593
rect 35713 20584 35725 20587
rect 34020 20556 35725 20584
rect 34020 20544 34026 20556
rect 35713 20553 35725 20556
rect 35759 20553 35771 20587
rect 35713 20547 35771 20553
rect 35894 20544 35900 20596
rect 35952 20544 35958 20596
rect 25317 20519 25375 20525
rect 25317 20485 25329 20519
rect 25363 20516 25375 20519
rect 28994 20516 29000 20528
rect 25363 20488 25728 20516
rect 25363 20485 25375 20488
rect 25317 20479 25375 20485
rect 25700 20460 25728 20488
rect 28828 20488 29000 20516
rect 24167 20420 24992 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 25038 20408 25044 20460
rect 25096 20448 25102 20460
rect 25133 20451 25191 20457
rect 25133 20448 25145 20451
rect 25096 20420 25145 20448
rect 25096 20408 25102 20420
rect 25133 20417 25145 20420
rect 25179 20417 25191 20451
rect 25133 20411 25191 20417
rect 25406 20408 25412 20460
rect 25464 20408 25470 20460
rect 25498 20408 25504 20460
rect 25556 20408 25562 20460
rect 25682 20408 25688 20460
rect 25740 20408 25746 20460
rect 25774 20408 25780 20460
rect 25832 20408 25838 20460
rect 28828 20457 28856 20488
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 35912 20516 35940 20544
rect 35912 20488 36032 20516
rect 28813 20451 28871 20457
rect 28813 20417 28825 20451
rect 28859 20417 28871 20451
rect 28813 20411 28871 20417
rect 28902 20408 28908 20460
rect 28960 20408 28966 20460
rect 29089 20451 29147 20457
rect 29089 20417 29101 20451
rect 29135 20417 29147 20451
rect 29089 20411 29147 20417
rect 29181 20451 29239 20457
rect 29181 20417 29193 20451
rect 29227 20448 29239 20451
rect 29362 20448 29368 20460
rect 29227 20420 29368 20448
rect 29227 20417 29239 20420
rect 29181 20411 29239 20417
rect 14516 20352 14964 20380
rect 15028 20352 15516 20380
rect 15580 20352 16804 20380
rect 14516 20340 14522 20352
rect 14734 20312 14740 20324
rect 14016 20284 14740 20312
rect 14734 20272 14740 20284
rect 14792 20272 14798 20324
rect 14936 20312 14964 20352
rect 15194 20312 15200 20324
rect 14936 20284 15200 20312
rect 15194 20272 15200 20284
rect 15252 20272 15258 20324
rect 14550 20244 14556 20256
rect 13918 20216 14556 20244
rect 14550 20204 14556 20216
rect 14608 20244 14614 20256
rect 15580 20244 15608 20352
rect 17034 20340 17040 20392
rect 17092 20340 17098 20392
rect 17678 20340 17684 20392
rect 17736 20340 17742 20392
rect 18046 20340 18052 20392
rect 18104 20380 18110 20392
rect 18690 20380 18696 20392
rect 18104 20352 18696 20380
rect 18104 20340 18110 20352
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 19889 20383 19947 20389
rect 19889 20349 19901 20383
rect 19935 20380 19947 20383
rect 20824 20380 20852 20408
rect 19935 20352 20852 20380
rect 23109 20383 23167 20389
rect 19935 20349 19947 20352
rect 19889 20343 19947 20349
rect 23109 20349 23121 20383
rect 23155 20380 23167 20383
rect 23750 20380 23756 20392
rect 23155 20352 23756 20380
rect 23155 20349 23167 20352
rect 23109 20343 23167 20349
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 25516 20380 25544 20408
rect 25792 20380 25820 20408
rect 25516 20352 25820 20380
rect 29104 20380 29132 20411
rect 29362 20408 29368 20420
rect 29420 20408 29426 20460
rect 29454 20408 29460 20460
rect 29512 20408 29518 20460
rect 29546 20408 29552 20460
rect 29604 20448 29610 20460
rect 29641 20451 29699 20457
rect 29641 20448 29653 20451
rect 29604 20420 29653 20448
rect 29604 20408 29610 20420
rect 29641 20417 29653 20420
rect 29687 20417 29699 20451
rect 29641 20411 29699 20417
rect 29825 20451 29883 20457
rect 29825 20417 29837 20451
rect 29871 20448 29883 20451
rect 30098 20448 30104 20460
rect 29871 20420 30104 20448
rect 29871 20417 29883 20420
rect 29825 20411 29883 20417
rect 30098 20408 30104 20420
rect 30156 20408 30162 20460
rect 34790 20408 34796 20460
rect 34848 20448 34854 20460
rect 36004 20457 36032 20488
rect 35161 20451 35219 20457
rect 35161 20448 35173 20451
rect 34848 20420 35173 20448
rect 34848 20408 34854 20420
rect 35161 20417 35173 20420
rect 35207 20417 35219 20451
rect 35161 20411 35219 20417
rect 35897 20451 35955 20457
rect 35897 20417 35909 20451
rect 35943 20417 35955 20451
rect 35897 20411 35955 20417
rect 35989 20451 36047 20457
rect 35989 20417 36001 20451
rect 36035 20417 36047 20451
rect 35989 20411 36047 20417
rect 29472 20380 29500 20408
rect 29914 20380 29920 20392
rect 29104 20352 29316 20380
rect 29472 20352 29920 20380
rect 15838 20272 15844 20324
rect 15896 20312 15902 20324
rect 19978 20312 19984 20324
rect 15896 20284 19984 20312
rect 15896 20272 15902 20284
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 23382 20272 23388 20324
rect 23440 20272 23446 20324
rect 24946 20272 24952 20324
rect 25004 20312 25010 20324
rect 27522 20312 27528 20324
rect 25004 20284 27528 20312
rect 25004 20272 25010 20284
rect 27522 20272 27528 20284
rect 27580 20312 27586 20324
rect 27580 20284 29132 20312
rect 27580 20272 27586 20284
rect 29104 20256 29132 20284
rect 29288 20256 29316 20352
rect 29914 20340 29920 20352
rect 29972 20340 29978 20392
rect 33870 20340 33876 20392
rect 33928 20380 33934 20392
rect 34422 20380 34428 20392
rect 33928 20352 34428 20380
rect 33928 20340 33934 20352
rect 34422 20340 34428 20352
rect 34480 20380 34486 20392
rect 35253 20383 35311 20389
rect 35253 20380 35265 20383
rect 34480 20352 35265 20380
rect 34480 20340 34486 20352
rect 35253 20349 35265 20352
rect 35299 20349 35311 20383
rect 35253 20343 35311 20349
rect 35434 20340 35440 20392
rect 35492 20340 35498 20392
rect 34793 20315 34851 20321
rect 34793 20281 34805 20315
rect 34839 20312 34851 20315
rect 35342 20312 35348 20324
rect 34839 20284 35348 20312
rect 34839 20281 34851 20284
rect 34793 20275 34851 20281
rect 35342 20272 35348 20284
rect 35400 20312 35406 20324
rect 35912 20312 35940 20411
rect 36170 20408 36176 20460
rect 36228 20408 36234 20460
rect 36262 20408 36268 20460
rect 36320 20408 36326 20460
rect 35400 20284 35940 20312
rect 35400 20272 35406 20284
rect 14608 20216 15608 20244
rect 14608 20204 14614 20216
rect 16206 20204 16212 20256
rect 16264 20244 16270 20256
rect 18966 20244 18972 20256
rect 16264 20216 18972 20244
rect 16264 20204 16270 20216
rect 18966 20204 18972 20216
rect 19024 20244 19030 20256
rect 20533 20247 20591 20253
rect 20533 20244 20545 20247
rect 19024 20216 20545 20244
rect 19024 20204 19030 20216
rect 20533 20213 20545 20216
rect 20579 20244 20591 20247
rect 21082 20244 21088 20256
rect 20579 20216 21088 20244
rect 20579 20213 20591 20216
rect 20533 20207 20591 20213
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 23198 20204 23204 20256
rect 23256 20204 23262 20256
rect 25685 20247 25743 20253
rect 25685 20213 25697 20247
rect 25731 20244 25743 20247
rect 28442 20244 28448 20256
rect 25731 20216 28448 20244
rect 25731 20213 25743 20216
rect 25685 20207 25743 20213
rect 28442 20204 28448 20216
rect 28500 20204 28506 20256
rect 28626 20204 28632 20256
rect 28684 20204 28690 20256
rect 29086 20204 29092 20256
rect 29144 20204 29150 20256
rect 29270 20204 29276 20256
rect 29328 20204 29334 20256
rect 29454 20204 29460 20256
rect 29512 20204 29518 20256
rect 1104 20154 38272 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38272 20154
rect 1104 20080 38272 20102
rect 7098 20000 7104 20052
rect 7156 20040 7162 20052
rect 7377 20043 7435 20049
rect 7377 20040 7389 20043
rect 7156 20012 7389 20040
rect 7156 20000 7162 20012
rect 7377 20009 7389 20012
rect 7423 20009 7435 20043
rect 7377 20003 7435 20009
rect 9306 20000 9312 20052
rect 9364 20040 9370 20052
rect 13998 20040 14004 20052
rect 9364 20012 14004 20040
rect 9364 20000 9370 20012
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 14090 20000 14096 20052
rect 14148 20040 14154 20052
rect 14645 20043 14703 20049
rect 14645 20040 14657 20043
rect 14148 20012 14657 20040
rect 14148 20000 14154 20012
rect 14645 20009 14657 20012
rect 14691 20009 14703 20043
rect 14645 20003 14703 20009
rect 15102 20000 15108 20052
rect 15160 20040 15166 20052
rect 16117 20043 16175 20049
rect 16117 20040 16129 20043
rect 15160 20012 16129 20040
rect 15160 20000 15166 20012
rect 16117 20009 16129 20012
rect 16163 20009 16175 20043
rect 16117 20003 16175 20009
rect 17402 20000 17408 20052
rect 17460 20040 17466 20052
rect 17865 20043 17923 20049
rect 17865 20040 17877 20043
rect 17460 20012 17877 20040
rect 17460 20000 17466 20012
rect 17865 20009 17877 20012
rect 17911 20009 17923 20043
rect 17865 20003 17923 20009
rect 18414 20000 18420 20052
rect 18472 20000 18478 20052
rect 18966 20000 18972 20052
rect 19024 20000 19030 20052
rect 20346 20000 20352 20052
rect 20404 20040 20410 20052
rect 20809 20043 20867 20049
rect 20809 20040 20821 20043
rect 20404 20012 20821 20040
rect 20404 20000 20410 20012
rect 20809 20009 20821 20012
rect 20855 20009 20867 20043
rect 20809 20003 20867 20009
rect 21450 20000 21456 20052
rect 21508 20000 21514 20052
rect 23198 20000 23204 20052
rect 23256 20040 23262 20052
rect 24397 20043 24455 20049
rect 24397 20040 24409 20043
rect 23256 20012 24409 20040
rect 23256 20000 23262 20012
rect 24397 20009 24409 20012
rect 24443 20009 24455 20043
rect 24397 20003 24455 20009
rect 26602 20000 26608 20052
rect 26660 20040 26666 20052
rect 26697 20043 26755 20049
rect 26697 20040 26709 20043
rect 26660 20012 26709 20040
rect 26660 20000 26666 20012
rect 26697 20009 26709 20012
rect 26743 20009 26755 20043
rect 28258 20040 28264 20052
rect 26697 20003 26755 20009
rect 26804 20012 28264 20040
rect 11606 19932 11612 19984
rect 11664 19972 11670 19984
rect 11790 19972 11796 19984
rect 11664 19944 11796 19972
rect 11664 19932 11670 19944
rect 11790 19932 11796 19944
rect 11848 19972 11854 19984
rect 11977 19975 12035 19981
rect 11977 19972 11989 19975
rect 11848 19944 11989 19972
rect 11848 19932 11854 19944
rect 11977 19941 11989 19944
rect 12023 19941 12035 19975
rect 11977 19935 12035 19941
rect 14366 19932 14372 19984
rect 14424 19932 14430 19984
rect 15381 19975 15439 19981
rect 15381 19972 15393 19975
rect 15304 19944 15393 19972
rect 3329 19907 3387 19913
rect 3329 19873 3341 19907
rect 3375 19904 3387 19907
rect 3878 19904 3884 19916
rect 3375 19876 3884 19904
rect 3375 19873 3387 19876
rect 3329 19867 3387 19873
rect 3878 19864 3884 19876
rect 3936 19864 3942 19916
rect 5718 19864 5724 19916
rect 5776 19864 5782 19916
rect 8018 19864 8024 19916
rect 8076 19904 8082 19916
rect 8297 19907 8355 19913
rect 8297 19904 8309 19907
rect 8076 19876 8309 19904
rect 8076 19864 8082 19876
rect 8297 19873 8309 19876
rect 8343 19873 8355 19907
rect 8297 19867 8355 19873
rect 8570 19864 8576 19916
rect 8628 19864 8634 19916
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19904 11759 19907
rect 11882 19904 11888 19916
rect 11747 19876 11888 19904
rect 11747 19873 11759 19876
rect 11701 19867 11759 19873
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 12308 19876 12357 19904
rect 12308 19864 12314 19876
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 12345 19867 12403 19873
rect 14734 19864 14740 19916
rect 14792 19864 14798 19916
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19904 14887 19907
rect 15194 19904 15200 19916
rect 14875 19876 15200 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15194 19864 15200 19876
rect 15252 19864 15258 19916
rect 15304 19913 15332 19944
rect 15381 19941 15393 19944
rect 15427 19972 15439 19975
rect 15654 19972 15660 19984
rect 15427 19944 15660 19972
rect 15427 19941 15439 19944
rect 15381 19935 15439 19941
rect 15654 19932 15660 19944
rect 15712 19932 15718 19984
rect 15838 19972 15844 19984
rect 15764 19944 15844 19972
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19873 15347 19907
rect 15289 19867 15347 19873
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19836 3111 19839
rect 3142 19836 3148 19848
rect 3099 19808 3148 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19836 4123 19839
rect 4154 19836 4160 19848
rect 4111 19808 4160 19836
rect 4111 19805 4123 19808
rect 4065 19799 4123 19805
rect 4154 19796 4160 19808
rect 4212 19836 4218 19848
rect 5442 19836 5448 19848
rect 4212 19808 5448 19836
rect 4212 19796 4218 19808
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 5629 19839 5687 19845
rect 5629 19805 5641 19839
rect 5675 19836 5687 19839
rect 5810 19836 5816 19848
rect 5675 19808 5816 19836
rect 5675 19805 5687 19808
rect 5629 19799 5687 19805
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 8205 19839 8263 19845
rect 7607 19808 7788 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 3234 19728 3240 19780
rect 3292 19768 3298 19780
rect 3292 19740 5948 19768
rect 3292 19728 3298 19740
rect 5920 19712 5948 19740
rect 2682 19660 2688 19712
rect 2740 19660 2746 19712
rect 3142 19660 3148 19712
rect 3200 19660 3206 19712
rect 3878 19660 3884 19712
rect 3936 19660 3942 19712
rect 5902 19660 5908 19712
rect 5960 19660 5966 19712
rect 5994 19660 6000 19712
rect 6052 19660 6058 19712
rect 7760 19709 7788 19808
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8588 19836 8616 19864
rect 12529 19839 12587 19845
rect 12529 19836 12541 19839
rect 8251 19808 8616 19836
rect 12406 19808 12541 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 11146 19768 11152 19780
rect 9916 19740 11152 19768
rect 9916 19728 9922 19740
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 7745 19703 7803 19709
rect 7745 19669 7757 19703
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 8113 19703 8171 19709
rect 8113 19669 8125 19703
rect 8159 19700 8171 19703
rect 9306 19700 9312 19712
rect 8159 19672 9312 19700
rect 8159 19669 8171 19672
rect 8113 19663 8171 19669
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 9582 19660 9588 19712
rect 9640 19700 9646 19712
rect 12161 19703 12219 19709
rect 12161 19700 12173 19703
rect 9640 19672 12173 19700
rect 9640 19660 9646 19672
rect 12161 19669 12173 19672
rect 12207 19700 12219 19703
rect 12406 19700 12434 19808
rect 12529 19805 12541 19808
rect 12575 19805 12587 19839
rect 12529 19799 12587 19805
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19836 14519 19839
rect 14752 19836 14780 19864
rect 14507 19808 14780 19836
rect 14921 19839 14979 19845
rect 14507 19805 14519 19808
rect 14461 19799 14519 19805
rect 14921 19805 14933 19839
rect 14967 19836 14979 19839
rect 14967 19808 15608 19836
rect 14967 19805 14979 19808
rect 14921 19799 14979 19805
rect 12802 19728 12808 19780
rect 12860 19768 12866 19780
rect 13446 19768 13452 19780
rect 12860 19740 13452 19768
rect 12860 19728 12866 19740
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 15197 19771 15255 19777
rect 15197 19737 15209 19771
rect 15243 19768 15255 19771
rect 15470 19768 15476 19780
rect 15243 19740 15476 19768
rect 15243 19737 15255 19740
rect 15197 19731 15255 19737
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 15580 19768 15608 19808
rect 15654 19796 15660 19848
rect 15712 19796 15718 19848
rect 15764 19845 15792 19944
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 20070 19972 20076 19984
rect 15948 19944 20076 19972
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19836 15899 19839
rect 15948 19836 15976 19944
rect 17034 19904 17040 19916
rect 16132 19876 17040 19904
rect 15887 19808 15976 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 16022 19796 16028 19848
rect 16080 19796 16086 19848
rect 16132 19845 16160 19876
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19836 16359 19839
rect 16482 19836 16488 19848
rect 16347 19808 16488 19836
rect 16347 19805 16359 19808
rect 16301 19799 16359 19805
rect 16132 19768 16160 19799
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 16850 19796 16856 19848
rect 16908 19836 16914 19848
rect 17313 19839 17371 19845
rect 17313 19836 17325 19839
rect 16908 19808 17325 19836
rect 16908 19796 16914 19808
rect 17313 19805 17325 19808
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 17586 19796 17592 19848
rect 17644 19796 17650 19848
rect 17728 19845 17756 19944
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 24210 19932 24216 19984
rect 24268 19972 24274 19984
rect 24765 19975 24823 19981
rect 24765 19972 24777 19975
rect 24268 19944 24777 19972
rect 24268 19932 24274 19944
rect 24765 19941 24777 19944
rect 24811 19941 24823 19975
rect 24765 19935 24823 19941
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 19426 19904 19432 19916
rect 17920 19876 19432 19904
rect 17920 19864 17926 19876
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 20220 19876 20545 19904
rect 20220 19864 20226 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 26804 19904 26832 20012
rect 27264 19913 27292 20012
rect 28258 20000 28264 20012
rect 28316 20000 28322 20052
rect 28445 20043 28503 20049
rect 28445 20009 28457 20043
rect 28491 20040 28503 20043
rect 28902 20040 28908 20052
rect 28491 20012 28908 20040
rect 28491 20009 28503 20012
rect 28445 20003 28503 20009
rect 28902 20000 28908 20012
rect 28960 20000 28966 20052
rect 34790 20000 34796 20052
rect 34848 20000 34854 20052
rect 35161 20043 35219 20049
rect 35161 20009 35173 20043
rect 35207 20040 35219 20043
rect 36170 20040 36176 20052
rect 35207 20012 36176 20040
rect 35207 20009 35219 20012
rect 35161 20003 35219 20009
rect 36170 20000 36176 20012
rect 36228 20000 36234 20052
rect 27801 19975 27859 19981
rect 27801 19941 27813 19975
rect 27847 19972 27859 19975
rect 29270 19972 29276 19984
rect 27847 19944 29276 19972
rect 27847 19941 27859 19944
rect 27801 19935 27859 19941
rect 29270 19932 29276 19944
rect 29328 19932 29334 19984
rect 34057 19975 34115 19981
rect 34057 19972 34069 19975
rect 33152 19944 34069 19972
rect 20533 19867 20591 19873
rect 23860 19876 26832 19904
rect 27249 19907 27307 19913
rect 17709 19839 17767 19845
rect 17709 19805 17721 19839
rect 17755 19805 17767 19839
rect 18542 19839 18600 19845
rect 18542 19836 18554 19839
rect 17709 19799 17767 19805
rect 17880 19808 18554 19836
rect 15580 19740 16160 19768
rect 12207 19672 12434 19700
rect 12207 19669 12219 19672
rect 12161 19663 12219 19669
rect 12618 19660 12624 19712
rect 12676 19700 12682 19712
rect 12713 19703 12771 19709
rect 12713 19700 12725 19703
rect 12676 19672 12725 19700
rect 12676 19660 12682 19672
rect 12713 19669 12725 19672
rect 12759 19669 12771 19703
rect 16500 19700 16528 19796
rect 17880 19780 17908 19808
rect 18542 19805 18554 19808
rect 18588 19805 18600 19839
rect 18542 19799 18600 19805
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19061 19839 19119 19845
rect 19061 19836 19073 19839
rect 18748 19808 19073 19836
rect 18748 19796 18754 19808
rect 19061 19805 19073 19808
rect 19107 19836 19119 19839
rect 19242 19836 19248 19848
rect 19107 19808 19248 19836
rect 19107 19805 19119 19808
rect 19061 19799 19119 19805
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 20625 19839 20683 19845
rect 20625 19836 20637 19839
rect 20548 19808 20637 19836
rect 17497 19771 17555 19777
rect 17497 19737 17509 19771
rect 17543 19737 17555 19771
rect 17497 19731 17555 19737
rect 17512 19700 17540 19731
rect 17862 19728 17868 19780
rect 17920 19728 17926 19780
rect 18414 19728 18420 19780
rect 18472 19768 18478 19780
rect 18472 19740 20208 19768
rect 18472 19728 18478 19740
rect 18601 19703 18659 19709
rect 18601 19700 18613 19703
rect 16500 19672 18613 19700
rect 12713 19663 12771 19669
rect 18601 19669 18613 19672
rect 18647 19700 18659 19703
rect 19058 19700 19064 19712
rect 18647 19672 19064 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 19058 19660 19064 19672
rect 19116 19660 19122 19712
rect 20180 19709 20208 19740
rect 20548 19712 20576 19808
rect 20625 19805 20637 19808
rect 20671 19805 20683 19839
rect 20625 19799 20683 19805
rect 22554 19796 22560 19848
rect 22612 19836 22618 19848
rect 23860 19845 23888 19876
rect 22741 19839 22799 19845
rect 22741 19836 22753 19839
rect 22612 19808 22753 19836
rect 22612 19796 22618 19808
rect 22741 19805 22753 19808
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19805 23903 19839
rect 24026 19836 24032 19848
rect 23845 19799 23903 19805
rect 23952 19808 24032 19836
rect 21177 19771 21235 19777
rect 21177 19768 21189 19771
rect 20732 19740 21189 19768
rect 20165 19703 20223 19709
rect 20165 19669 20177 19703
rect 20211 19669 20223 19703
rect 20165 19663 20223 19669
rect 20530 19660 20536 19712
rect 20588 19660 20594 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 20732 19700 20760 19740
rect 21177 19737 21189 19740
rect 21223 19737 21235 19771
rect 21177 19731 21235 19737
rect 22922 19728 22928 19780
rect 22980 19768 22986 19780
rect 23569 19771 23627 19777
rect 23569 19768 23581 19771
rect 22980 19740 23581 19768
rect 22980 19728 22986 19740
rect 23569 19737 23581 19740
rect 23615 19768 23627 19771
rect 23952 19768 23980 19808
rect 24026 19796 24032 19808
rect 24084 19836 24090 19848
rect 24596 19845 24624 19876
rect 27249 19873 27261 19907
rect 27295 19873 27307 19907
rect 27890 19904 27896 19916
rect 27249 19867 27307 19873
rect 27816 19876 27896 19904
rect 24581 19839 24639 19845
rect 24084 19808 24262 19836
rect 24084 19796 24090 19808
rect 23615 19740 23980 19768
rect 24234 19768 24262 19808
rect 24581 19805 24593 19839
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 24670 19796 24676 19848
rect 24728 19796 24734 19848
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19836 24915 19839
rect 24946 19836 24952 19848
rect 24903 19808 24952 19836
rect 24903 19805 24915 19808
rect 24857 19799 24915 19805
rect 24872 19768 24900 19799
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 25590 19836 25596 19848
rect 25547 19808 25596 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 25866 19796 25872 19848
rect 25924 19796 25930 19848
rect 25958 19796 25964 19848
rect 26016 19836 26022 19848
rect 26790 19839 26848 19845
rect 26790 19836 26802 19839
rect 26016 19808 26802 19836
rect 26016 19796 26022 19808
rect 26790 19805 26802 19808
rect 26836 19805 26848 19839
rect 26790 19799 26848 19805
rect 26878 19796 26884 19848
rect 26936 19836 26942 19848
rect 27816 19845 27844 19876
rect 27890 19864 27896 19876
rect 27948 19904 27954 19916
rect 27948 19876 28396 19904
rect 27948 19864 27954 19876
rect 27157 19839 27215 19845
rect 27157 19836 27169 19839
rect 26936 19808 27169 19836
rect 26936 19796 26942 19808
rect 27157 19805 27169 19808
rect 27203 19805 27215 19839
rect 27801 19839 27859 19845
rect 27801 19836 27813 19839
rect 27157 19799 27215 19805
rect 27586 19808 27813 19836
rect 24234 19740 24900 19768
rect 23615 19737 23627 19740
rect 23569 19731 23627 19737
rect 25682 19728 25688 19780
rect 25740 19728 25746 19780
rect 25774 19728 25780 19780
rect 25832 19728 25838 19780
rect 27586 19768 27614 19808
rect 27801 19805 27813 19808
rect 27847 19805 27859 19839
rect 27801 19799 27859 19805
rect 27985 19839 28043 19845
rect 27985 19805 27997 19839
rect 28031 19836 28043 19839
rect 28074 19836 28080 19848
rect 28031 19808 28080 19836
rect 28031 19805 28043 19808
rect 27985 19799 28043 19805
rect 28074 19796 28080 19808
rect 28132 19796 28138 19848
rect 28368 19845 28396 19876
rect 28442 19864 28448 19916
rect 28500 19904 28506 19916
rect 28813 19907 28871 19913
rect 28500 19876 28672 19904
rect 28500 19864 28506 19876
rect 28353 19839 28411 19845
rect 28353 19805 28365 19839
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 28537 19839 28595 19845
rect 28537 19805 28549 19839
rect 28583 19805 28595 19839
rect 28537 19799 28595 19805
rect 26068 19740 27614 19768
rect 28092 19768 28120 19796
rect 28552 19768 28580 19799
rect 28092 19740 28580 19768
rect 28644 19768 28672 19876
rect 28813 19873 28825 19907
rect 28859 19904 28871 19907
rect 28994 19904 29000 19916
rect 28859 19876 29000 19904
rect 28859 19873 28871 19876
rect 28813 19867 28871 19873
rect 28994 19864 29000 19876
rect 29052 19864 29058 19916
rect 28718 19796 28724 19848
rect 28776 19836 28782 19848
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 28776 19808 28917 19836
rect 28776 19796 28782 19808
rect 28905 19805 28917 19808
rect 28951 19836 28963 19839
rect 29546 19836 29552 19848
rect 28951 19808 29552 19836
rect 28951 19805 28963 19808
rect 28905 19799 28963 19805
rect 29546 19796 29552 19808
rect 29604 19796 29610 19848
rect 29914 19796 29920 19848
rect 29972 19796 29978 19848
rect 30098 19796 30104 19848
rect 30156 19796 30162 19848
rect 33152 19845 33180 19944
rect 34057 19941 34069 19944
rect 34103 19941 34115 19975
rect 34057 19935 34115 19941
rect 34425 19975 34483 19981
rect 34425 19941 34437 19975
rect 34471 19972 34483 19975
rect 34698 19972 34704 19984
rect 34471 19944 34704 19972
rect 34471 19941 34483 19944
rect 34425 19935 34483 19941
rect 33137 19839 33195 19845
rect 33137 19836 33149 19839
rect 30208 19808 33149 19836
rect 30208 19768 30236 19808
rect 33137 19805 33149 19808
rect 33183 19805 33195 19839
rect 33137 19799 33195 19805
rect 33226 19796 33232 19848
rect 33284 19836 33290 19848
rect 33321 19839 33379 19845
rect 33321 19836 33333 19839
rect 33284 19808 33333 19836
rect 33284 19796 33290 19808
rect 33321 19805 33333 19808
rect 33367 19836 33379 19839
rect 33781 19839 33839 19845
rect 33781 19836 33793 19839
rect 33367 19808 33793 19836
rect 33367 19805 33379 19808
rect 33321 19799 33379 19805
rect 33781 19805 33793 19808
rect 33827 19805 33839 19839
rect 34072 19836 34100 19935
rect 34698 19932 34704 19944
rect 34756 19932 34762 19984
rect 34808 19972 34836 20000
rect 34977 19975 35035 19981
rect 34977 19972 34989 19975
rect 34808 19944 34989 19972
rect 34977 19941 34989 19944
rect 35023 19941 35035 19975
rect 34977 19935 35035 19941
rect 35342 19932 35348 19984
rect 35400 19932 35406 19984
rect 34716 19904 34744 19932
rect 35360 19904 35388 19932
rect 34716 19876 35112 19904
rect 35084 19848 35112 19876
rect 35176 19876 35388 19904
rect 34333 19839 34391 19845
rect 34333 19836 34345 19839
rect 34072 19808 34345 19836
rect 33781 19799 33839 19805
rect 34333 19805 34345 19808
rect 34379 19805 34391 19839
rect 34333 19799 34391 19805
rect 34517 19839 34575 19845
rect 34517 19805 34529 19839
rect 34563 19805 34575 19839
rect 34517 19799 34575 19805
rect 34885 19839 34943 19845
rect 34885 19805 34897 19839
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 28644 19740 30236 19768
rect 20680 19672 20760 19700
rect 20680 19660 20686 19672
rect 23934 19660 23940 19712
rect 23992 19700 23998 19712
rect 24394 19700 24400 19712
rect 23992 19672 24400 19700
rect 23992 19660 23998 19672
rect 24394 19660 24400 19672
rect 24452 19660 24458 19712
rect 25590 19660 25596 19712
rect 25648 19700 25654 19712
rect 25700 19700 25728 19728
rect 26068 19709 26096 19740
rect 30282 19728 30288 19780
rect 30340 19728 30346 19780
rect 30377 19771 30435 19777
rect 30377 19737 30389 19771
rect 30423 19768 30435 19771
rect 30834 19768 30840 19780
rect 30423 19740 30840 19768
rect 30423 19737 30435 19740
rect 30377 19731 30435 19737
rect 30834 19728 30840 19740
rect 30892 19728 30898 19780
rect 33796 19768 33824 19799
rect 34532 19768 34560 19799
rect 33796 19740 34560 19768
rect 25648 19672 25728 19700
rect 26053 19703 26111 19709
rect 25648 19660 25654 19672
rect 26053 19669 26065 19703
rect 26099 19669 26111 19703
rect 26053 19663 26111 19669
rect 28166 19660 28172 19712
rect 28224 19660 28230 19712
rect 28258 19660 28264 19712
rect 28316 19700 28322 19712
rect 29178 19700 29184 19712
rect 28316 19672 29184 19700
rect 28316 19660 28322 19672
rect 29178 19660 29184 19672
rect 29236 19660 29242 19712
rect 29273 19703 29331 19709
rect 29273 19669 29285 19703
rect 29319 19700 29331 19703
rect 30466 19700 30472 19712
rect 29319 19672 30472 19700
rect 29319 19669 29331 19672
rect 29273 19663 29331 19669
rect 30466 19660 30472 19672
rect 30524 19660 30530 19712
rect 33226 19660 33232 19712
rect 33284 19660 33290 19712
rect 34238 19660 34244 19712
rect 34296 19660 34302 19712
rect 34514 19660 34520 19712
rect 34572 19700 34578 19712
rect 34900 19700 34928 19799
rect 35066 19796 35072 19848
rect 35124 19796 35130 19848
rect 35176 19845 35204 19876
rect 35161 19839 35219 19845
rect 35161 19805 35173 19839
rect 35207 19805 35219 19839
rect 35161 19799 35219 19805
rect 35345 19839 35403 19845
rect 35345 19805 35357 19839
rect 35391 19836 35403 19839
rect 35894 19836 35900 19848
rect 35391 19808 35900 19836
rect 35391 19805 35403 19808
rect 35345 19799 35403 19805
rect 35894 19796 35900 19808
rect 35952 19796 35958 19848
rect 34572 19672 34928 19700
rect 34572 19660 34578 19672
rect 1104 19610 38272 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38272 19610
rect 1104 19536 38272 19558
rect 2682 19456 2688 19508
rect 2740 19456 2746 19508
rect 4706 19496 4712 19508
rect 4264 19468 4712 19496
rect 1946 19320 1952 19372
rect 2004 19320 2010 19372
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 2700 19360 2728 19456
rect 4264 19369 4292 19468
rect 4706 19456 4712 19468
rect 4764 19496 4770 19508
rect 6914 19496 6920 19508
rect 4764 19468 6920 19496
rect 4764 19456 4770 19468
rect 6914 19456 6920 19468
rect 6972 19456 6978 19508
rect 9306 19456 9312 19508
rect 9364 19456 9370 19508
rect 10781 19499 10839 19505
rect 10781 19465 10793 19499
rect 10827 19496 10839 19499
rect 10827 19468 11008 19496
rect 10827 19465 10839 19468
rect 10781 19459 10839 19465
rect 5994 19388 6000 19440
rect 6052 19428 6058 19440
rect 6549 19431 6607 19437
rect 6549 19428 6561 19431
rect 6052 19400 6561 19428
rect 6052 19388 6058 19400
rect 6549 19397 6561 19400
rect 6595 19397 6607 19431
rect 6549 19391 6607 19397
rect 6641 19431 6699 19437
rect 6641 19397 6653 19431
rect 6687 19428 6699 19431
rect 9324 19428 9352 19456
rect 10870 19428 10876 19440
rect 6687 19400 8708 19428
rect 9324 19400 10876 19428
rect 6687 19397 6699 19400
rect 6641 19391 6699 19397
rect 8680 19372 8708 19400
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 10980 19428 11008 19468
rect 11146 19456 11152 19508
rect 11204 19496 11210 19508
rect 15102 19496 15108 19508
rect 11204 19468 15108 19496
rect 11204 19456 11210 19468
rect 15102 19456 15108 19468
rect 15160 19456 15166 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15562 19496 15568 19508
rect 15252 19468 15568 19496
rect 15252 19456 15258 19468
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 24305 19499 24363 19505
rect 16632 19468 20760 19496
rect 16632 19456 16638 19468
rect 11054 19428 11060 19440
rect 10980 19400 11060 19428
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 12360 19400 15056 19428
rect 2271 19332 2728 19360
rect 4249 19363 4307 19369
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 4249 19329 4261 19363
rect 4295 19329 4307 19363
rect 5902 19360 5908 19372
rect 5658 19332 5908 19360
rect 4249 19323 4307 19329
rect 5902 19320 5908 19332
rect 5960 19320 5966 19372
rect 6362 19320 6368 19372
rect 6420 19360 6426 19372
rect 6420 19332 6684 19360
rect 6420 19320 6426 19332
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19261 2099 19295
rect 2041 19255 2099 19261
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 4614 19292 4620 19304
rect 4571 19264 4620 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 2056 19168 2084 19255
rect 4614 19252 4620 19264
rect 4672 19252 4678 19304
rect 6656 19292 6684 19332
rect 6730 19320 6736 19372
rect 6788 19320 6794 19372
rect 7190 19320 7196 19372
rect 7248 19320 7254 19372
rect 7558 19320 7564 19372
rect 7616 19360 7622 19372
rect 7653 19363 7711 19369
rect 7653 19360 7665 19363
rect 7616 19332 7665 19360
rect 7616 19320 7622 19332
rect 7653 19329 7665 19332
rect 7699 19329 7711 19363
rect 7653 19323 7711 19329
rect 8662 19320 8668 19372
rect 8720 19320 8726 19372
rect 9125 19363 9183 19369
rect 9125 19329 9137 19363
rect 9171 19360 9183 19363
rect 9582 19360 9588 19372
rect 9171 19332 9588 19360
rect 9171 19329 9183 19332
rect 9125 19323 9183 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 10413 19363 10471 19369
rect 10413 19329 10425 19363
rect 10459 19360 10471 19363
rect 10962 19360 10968 19372
rect 10459 19332 10968 19360
rect 10459 19329 10471 19332
rect 10413 19323 10471 19329
rect 10962 19320 10968 19332
rect 11020 19360 11026 19372
rect 12360 19364 12388 19400
rect 12176 19360 12388 19364
rect 11020 19336 12388 19360
rect 11020 19332 12204 19336
rect 11020 19320 11026 19332
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 13044 19332 13369 19360
rect 13044 19320 13050 19332
rect 13357 19329 13369 19332
rect 13403 19360 13415 19363
rect 13541 19363 13599 19369
rect 13403 19332 13492 19360
rect 13403 19329 13415 19332
rect 13357 19323 13415 19329
rect 7208 19292 7236 19320
rect 6656 19264 7236 19292
rect 8938 19252 8944 19304
rect 8996 19252 9002 19304
rect 10505 19295 10563 19301
rect 10505 19261 10517 19295
rect 10551 19292 10563 19295
rect 10778 19292 10784 19304
rect 10551 19264 10784 19292
rect 10551 19261 10563 19264
rect 10505 19255 10563 19261
rect 10778 19252 10784 19264
rect 10836 19292 10842 19304
rect 11514 19292 11520 19304
rect 10836 19264 11520 19292
rect 10836 19252 10842 19264
rect 11514 19252 11520 19264
rect 11572 19292 11578 19304
rect 12526 19292 12532 19304
rect 11572 19264 12532 19292
rect 11572 19252 11578 19264
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 6822 19184 6828 19236
rect 6880 19224 6886 19236
rect 11882 19224 11888 19236
rect 6880 19196 11888 19224
rect 6880 19184 6886 19196
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 12710 19184 12716 19236
rect 12768 19224 12774 19236
rect 13464 19224 13492 19332
rect 13541 19329 13553 19363
rect 13587 19360 13599 19363
rect 13814 19360 13820 19372
rect 13587 19332 13820 19360
rect 13587 19329 13599 19332
rect 13541 19323 13599 19329
rect 13814 19320 13820 19332
rect 13872 19320 13878 19372
rect 14918 19360 14924 19372
rect 13924 19332 14924 19360
rect 13630 19252 13636 19304
rect 13688 19252 13694 19304
rect 13924 19224 13952 19332
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 15028 19360 15056 19400
rect 15212 19400 17264 19428
rect 15212 19360 15240 19400
rect 15028 19332 15240 19360
rect 15470 19320 15476 19372
rect 15528 19360 15534 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 15528 19332 16865 19360
rect 15528 19320 15534 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 17236 19360 17264 19400
rect 17586 19388 17592 19440
rect 17644 19388 17650 19440
rect 20162 19428 20168 19440
rect 17696 19400 20168 19428
rect 17696 19360 17724 19400
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 20732 19428 20760 19468
rect 24305 19465 24317 19499
rect 24351 19496 24363 19499
rect 24762 19496 24768 19508
rect 24351 19468 24768 19496
rect 24351 19465 24363 19468
rect 24305 19459 24363 19465
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 25869 19499 25927 19505
rect 25869 19465 25881 19499
rect 25915 19496 25927 19499
rect 25958 19496 25964 19508
rect 25915 19468 25964 19496
rect 25915 19465 25927 19468
rect 25869 19459 25927 19465
rect 20272 19400 20673 19428
rect 17236 19332 17724 19360
rect 16853 19323 16911 19329
rect 18690 19320 18696 19372
rect 18748 19320 18754 19372
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 15160 19264 17908 19292
rect 15160 19252 15166 19264
rect 12768 19196 13308 19224
rect 13464 19196 13952 19224
rect 12768 19184 12774 19196
rect 1762 19116 1768 19168
rect 1820 19116 1826 19168
rect 2038 19116 2044 19168
rect 2096 19116 2102 19168
rect 2406 19116 2412 19168
rect 2464 19116 2470 19168
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 5994 19156 6000 19168
rect 5868 19128 6000 19156
rect 5868 19116 5874 19128
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 6917 19159 6975 19165
rect 6917 19125 6929 19159
rect 6963 19156 6975 19159
rect 7006 19156 7012 19168
rect 6963 19128 7012 19156
rect 6963 19125 6975 19128
rect 6917 19119 6975 19125
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7466 19116 7472 19168
rect 7524 19116 7530 19168
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 13078 19156 13084 19168
rect 9364 19128 13084 19156
rect 9364 19116 9370 19128
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 13170 19116 13176 19168
rect 13228 19116 13234 19168
rect 13280 19156 13308 19196
rect 17126 19184 17132 19236
rect 17184 19224 17190 19236
rect 17221 19227 17279 19233
rect 17221 19224 17233 19227
rect 17184 19196 17233 19224
rect 17184 19184 17190 19196
rect 17221 19193 17233 19196
rect 17267 19193 17279 19227
rect 17221 19187 17279 19193
rect 17770 19184 17776 19236
rect 17828 19184 17834 19236
rect 17880 19224 17908 19264
rect 18598 19252 18604 19304
rect 18656 19252 18662 19304
rect 18892 19292 18920 19323
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19337 19363 19395 19369
rect 19337 19360 19349 19363
rect 19116 19332 19349 19360
rect 19116 19320 19122 19332
rect 19337 19329 19349 19332
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19484 19332 19717 19360
rect 19484 19320 19490 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19978 19320 19984 19372
rect 20036 19334 20042 19372
rect 20036 19320 20116 19334
rect 19996 19306 20116 19320
rect 18966 19292 18972 19304
rect 18892 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19889 19295 19947 19301
rect 19889 19261 19901 19295
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 20088 19292 20116 19306
rect 20272 19304 20300 19400
rect 20533 19363 20591 19369
rect 20533 19358 20545 19363
rect 20457 19330 20545 19358
rect 20254 19292 20260 19304
rect 20088 19264 20260 19292
rect 19904 19224 19932 19255
rect 20088 19224 20116 19264
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 17880 19196 19334 19224
rect 19904 19196 20116 19224
rect 14918 19156 14924 19168
rect 13280 19128 14924 19156
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 16945 19159 17003 19165
rect 16945 19125 16957 19159
rect 16991 19156 17003 19159
rect 17494 19156 17500 19168
rect 16991 19128 17500 19156
rect 16991 19125 17003 19128
rect 16945 19119 17003 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19156 17647 19159
rect 18966 19156 18972 19168
rect 17635 19128 18972 19156
rect 17635 19125 17647 19128
rect 17589 19119 17647 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 19306 19156 19334 19196
rect 19886 19156 19892 19168
rect 19306 19128 19892 19156
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 20457 19156 20485 19330
rect 20533 19329 20545 19330
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 20645 19292 20673 19400
rect 20732 19400 22968 19428
rect 20732 19369 20760 19400
rect 22940 19372 22968 19400
rect 24210 19388 24216 19440
rect 24268 19428 24274 19440
rect 24489 19431 24547 19437
rect 24489 19428 24501 19431
rect 24268 19400 24501 19428
rect 24268 19388 24274 19400
rect 24489 19397 24501 19400
rect 24535 19397 24547 19431
rect 25884 19428 25912 19459
rect 25958 19456 25964 19468
rect 26016 19456 26022 19508
rect 26418 19456 26424 19508
rect 26476 19496 26482 19508
rect 26605 19499 26663 19505
rect 26605 19496 26617 19499
rect 26476 19468 26617 19496
rect 26476 19456 26482 19468
rect 26605 19465 26617 19468
rect 26651 19465 26663 19499
rect 26605 19459 26663 19465
rect 27338 19456 27344 19508
rect 27396 19496 27402 19508
rect 27433 19499 27491 19505
rect 27433 19496 27445 19499
rect 27396 19468 27445 19496
rect 27396 19456 27402 19468
rect 27433 19465 27445 19468
rect 27479 19465 27491 19499
rect 27433 19459 27491 19465
rect 28166 19456 28172 19508
rect 28224 19456 28230 19508
rect 30006 19496 30012 19508
rect 28552 19468 30012 19496
rect 24489 19391 24547 19397
rect 24596 19400 25912 19428
rect 26237 19431 26295 19437
rect 20717 19363 20775 19369
rect 20717 19329 20729 19363
rect 20763 19329 20775 19363
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20717 19323 20775 19329
rect 20870 19332 21005 19360
rect 20870 19292 20898 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 22186 19320 22192 19372
rect 22244 19320 22250 19372
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19360 22523 19363
rect 22554 19360 22560 19372
rect 22511 19332 22560 19360
rect 22511 19329 22523 19332
rect 22465 19323 22523 19329
rect 22554 19320 22560 19332
rect 22612 19320 22618 19372
rect 22922 19320 22928 19372
rect 22980 19320 22986 19372
rect 23017 19363 23075 19369
rect 23017 19329 23029 19363
rect 23063 19360 23075 19363
rect 23474 19360 23480 19372
rect 23063 19332 23480 19360
rect 23063 19329 23075 19332
rect 23017 19323 23075 19329
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 23753 19363 23811 19369
rect 23753 19329 23765 19363
rect 23799 19360 23811 19363
rect 23842 19360 23848 19372
rect 23799 19332 23848 19360
rect 23799 19329 23811 19332
rect 23753 19323 23811 19329
rect 20645 19264 20898 19292
rect 22646 19252 22652 19304
rect 22704 19252 22710 19304
rect 23768 19292 23796 19323
rect 23842 19320 23848 19332
rect 23900 19320 23906 19372
rect 23937 19363 23995 19369
rect 23937 19329 23949 19363
rect 23983 19329 23995 19363
rect 23937 19323 23995 19329
rect 24029 19363 24087 19369
rect 24029 19329 24041 19363
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 24121 19363 24179 19369
rect 24121 19329 24133 19363
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 22756 19264 23796 19292
rect 20898 19184 20904 19236
rect 20956 19184 20962 19236
rect 22756 19224 22784 19264
rect 21008 19196 22784 19224
rect 21008 19156 21036 19196
rect 23290 19184 23296 19236
rect 23348 19184 23354 19236
rect 20457 19128 21036 19156
rect 23842 19116 23848 19168
rect 23900 19156 23906 19168
rect 23952 19156 23980 19323
rect 24044 19224 24072 19323
rect 24136 19292 24164 19323
rect 24394 19320 24400 19372
rect 24452 19320 24458 19372
rect 24596 19369 24624 19400
rect 26237 19397 26249 19431
rect 26283 19428 26295 19431
rect 26283 19400 26832 19428
rect 26283 19397 26295 19400
rect 26237 19391 26295 19397
rect 26804 19372 26832 19400
rect 24581 19363 24639 19369
rect 24581 19329 24593 19363
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 25682 19320 25688 19372
rect 25740 19320 25746 19372
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19329 25927 19363
rect 25869 19323 25927 19329
rect 25884 19292 25912 19323
rect 26050 19320 26056 19372
rect 26108 19320 26114 19372
rect 26326 19360 26332 19372
rect 26160 19332 26332 19360
rect 26160 19292 26188 19332
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 26421 19363 26479 19369
rect 26421 19329 26433 19363
rect 26467 19329 26479 19363
rect 26421 19323 26479 19329
rect 26436 19292 26464 19323
rect 26602 19320 26608 19372
rect 26660 19320 26666 19372
rect 26786 19320 26792 19372
rect 26844 19320 26850 19372
rect 27157 19363 27215 19369
rect 27157 19329 27169 19363
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 24136 19264 24256 19292
rect 24118 19224 24124 19236
rect 24044 19196 24124 19224
rect 24118 19184 24124 19196
rect 24176 19184 24182 19236
rect 24228 19224 24256 19264
rect 25056 19264 26188 19292
rect 26350 19264 26464 19292
rect 26620 19292 26648 19320
rect 27172 19292 27200 19323
rect 27246 19320 27252 19372
rect 27304 19360 27310 19372
rect 27341 19363 27399 19369
rect 27341 19360 27353 19363
rect 27304 19332 27353 19360
rect 27304 19320 27310 19332
rect 27341 19329 27353 19332
rect 27387 19329 27399 19363
rect 27341 19323 27399 19329
rect 27890 19320 27896 19372
rect 27948 19360 27954 19372
rect 28077 19363 28135 19369
rect 28077 19360 28089 19363
rect 27948 19332 28089 19360
rect 27948 19320 27954 19332
rect 28077 19329 28089 19332
rect 28123 19329 28135 19363
rect 28184 19360 28212 19456
rect 28552 19369 28580 19468
rect 30006 19456 30012 19468
rect 30064 19456 30070 19508
rect 30282 19456 30288 19508
rect 30340 19456 30346 19508
rect 30466 19456 30472 19508
rect 30524 19456 30530 19508
rect 33226 19456 33232 19508
rect 33284 19456 33290 19508
rect 34422 19456 34428 19508
rect 34480 19456 34486 19508
rect 35066 19456 35072 19508
rect 35124 19456 35130 19508
rect 29178 19388 29184 19440
rect 29236 19428 29242 19440
rect 29236 19400 29592 19428
rect 29236 19388 29242 19400
rect 28261 19363 28319 19369
rect 28261 19360 28273 19363
rect 28184 19332 28273 19360
rect 28077 19323 28135 19329
rect 28261 19329 28273 19332
rect 28307 19329 28319 19363
rect 28261 19323 28319 19329
rect 28537 19363 28595 19369
rect 28537 19329 28549 19363
rect 28583 19329 28595 19363
rect 28537 19323 28595 19329
rect 28626 19320 28632 19372
rect 28684 19360 28690 19372
rect 28812 19363 28870 19369
rect 28812 19360 28824 19363
rect 28684 19332 28824 19360
rect 28684 19320 28690 19332
rect 28812 19329 28824 19332
rect 28858 19329 28870 19363
rect 28812 19323 28870 19329
rect 28994 19320 29000 19372
rect 29052 19320 29058 19372
rect 29089 19363 29147 19369
rect 29089 19329 29101 19363
rect 29135 19360 29147 19363
rect 29270 19360 29276 19372
rect 29135 19332 29276 19360
rect 29135 19329 29147 19332
rect 29089 19323 29147 19329
rect 29270 19320 29276 19332
rect 29328 19320 29334 19372
rect 29454 19320 29460 19372
rect 29512 19320 29518 19372
rect 26620 19264 27200 19292
rect 28169 19295 28227 19301
rect 24302 19224 24308 19236
rect 24228 19196 24308 19224
rect 24302 19184 24308 19196
rect 24360 19184 24366 19236
rect 23900 19128 23980 19156
rect 24136 19156 24164 19184
rect 24854 19156 24860 19168
rect 24136 19128 24860 19156
rect 23900 19116 23906 19128
rect 24854 19116 24860 19128
rect 24912 19156 24918 19168
rect 25056 19156 25084 19264
rect 26350 19224 26378 19264
rect 28169 19261 28181 19295
rect 28215 19292 28227 19295
rect 28721 19295 28779 19301
rect 28721 19292 28733 19295
rect 28215 19264 28733 19292
rect 28215 19261 28227 19264
rect 28169 19255 28227 19261
rect 28721 19261 28733 19264
rect 28767 19261 28779 19295
rect 28721 19255 28779 19261
rect 25148 19196 26378 19224
rect 28629 19227 28687 19233
rect 25148 19168 25176 19196
rect 28629 19193 28641 19227
rect 28675 19193 28687 19227
rect 29472 19224 29500 19320
rect 29564 19292 29592 19400
rect 30009 19363 30067 19369
rect 30009 19329 30021 19363
rect 30055 19360 30067 19363
rect 30300 19360 30328 19456
rect 30484 19428 30512 19456
rect 30392 19400 30512 19428
rect 30392 19369 30420 19400
rect 30742 19388 30748 19440
rect 30800 19428 30806 19440
rect 31202 19428 31208 19440
rect 30800 19400 31208 19428
rect 30800 19388 30806 19400
rect 31202 19388 31208 19400
rect 31260 19428 31266 19440
rect 31665 19431 31723 19437
rect 31260 19400 31616 19428
rect 31260 19388 31266 19400
rect 30055 19332 30328 19360
rect 30377 19363 30435 19369
rect 30055 19329 30067 19332
rect 30009 19323 30067 19329
rect 30377 19329 30389 19363
rect 30423 19329 30435 19363
rect 30377 19323 30435 19329
rect 30466 19320 30472 19372
rect 30524 19320 30530 19372
rect 31588 19369 31616 19400
rect 31665 19397 31677 19431
rect 31711 19428 31723 19431
rect 33244 19428 33272 19456
rect 33965 19431 34023 19437
rect 31711 19400 32352 19428
rect 31711 19397 31723 19400
rect 31665 19391 31723 19397
rect 31113 19363 31171 19369
rect 31113 19360 31125 19363
rect 30852 19332 31125 19360
rect 30852 19292 30880 19332
rect 31113 19329 31125 19332
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19329 31631 19363
rect 31573 19323 31631 19329
rect 31938 19320 31944 19372
rect 31996 19360 32002 19372
rect 32324 19369 32352 19400
rect 32416 19400 32720 19428
rect 32416 19372 32444 19400
rect 32125 19363 32183 19369
rect 32125 19360 32137 19363
rect 31996 19332 32137 19360
rect 31996 19320 32002 19332
rect 32125 19329 32137 19332
rect 32171 19329 32183 19363
rect 32125 19323 32183 19329
rect 32309 19363 32367 19369
rect 32309 19329 32321 19363
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 32398 19320 32404 19372
rect 32456 19320 32462 19372
rect 32582 19320 32588 19372
rect 32640 19320 32646 19372
rect 32692 19369 32720 19400
rect 32876 19400 33916 19428
rect 32876 19369 32904 19400
rect 33888 19369 33916 19400
rect 33965 19397 33977 19431
rect 34011 19428 34023 19431
rect 34011 19400 35020 19428
rect 34011 19397 34023 19400
rect 33965 19391 34023 19397
rect 32677 19363 32735 19369
rect 32677 19329 32689 19363
rect 32723 19329 32735 19363
rect 32677 19323 32735 19329
rect 32861 19363 32919 19369
rect 32861 19329 32873 19363
rect 32907 19329 32919 19363
rect 32861 19323 32919 19329
rect 32953 19363 33011 19369
rect 32953 19329 32965 19363
rect 32999 19329 33011 19363
rect 32953 19323 33011 19329
rect 33873 19363 33931 19369
rect 33873 19329 33885 19363
rect 33919 19329 33931 19363
rect 33873 19323 33931 19329
rect 29564 19264 30880 19292
rect 30852 19233 30880 19264
rect 30926 19252 30932 19304
rect 30984 19292 30990 19304
rect 31021 19295 31079 19301
rect 31021 19292 31033 19295
rect 30984 19264 31033 19292
rect 30984 19252 30990 19264
rect 31021 19261 31033 19264
rect 31067 19261 31079 19295
rect 31021 19255 31079 19261
rect 31481 19295 31539 19301
rect 31481 19261 31493 19295
rect 31527 19292 31539 19295
rect 31527 19264 31754 19292
rect 31527 19261 31539 19264
rect 31481 19255 31539 19261
rect 28629 19187 28687 19193
rect 28920 19196 29500 19224
rect 30837 19227 30895 19233
rect 24912 19128 25084 19156
rect 24912 19116 24918 19128
rect 25130 19116 25136 19168
rect 25188 19116 25194 19168
rect 28350 19116 28356 19168
rect 28408 19116 28414 19168
rect 28644 19156 28672 19187
rect 28920 19156 28948 19196
rect 30837 19193 30849 19227
rect 30883 19193 30895 19227
rect 30837 19187 30895 19193
rect 28644 19128 28948 19156
rect 29178 19116 29184 19168
rect 29236 19116 29242 19168
rect 29362 19116 29368 19168
rect 29420 19156 29426 19168
rect 30466 19156 30472 19168
rect 29420 19128 30472 19156
rect 29420 19116 29426 19128
rect 30466 19116 30472 19128
rect 30524 19156 30530 19168
rect 31294 19156 31300 19168
rect 30524 19128 31300 19156
rect 30524 19116 30530 19128
rect 31294 19116 31300 19128
rect 31352 19116 31358 19168
rect 31726 19156 31754 19264
rect 32214 19252 32220 19304
rect 32272 19292 32278 19304
rect 32968 19292 32996 19323
rect 34238 19320 34244 19372
rect 34296 19360 34302 19372
rect 34992 19369 35020 19400
rect 34609 19363 34667 19369
rect 34609 19360 34621 19363
rect 34296 19332 34621 19360
rect 34296 19320 34302 19332
rect 34609 19329 34621 19332
rect 34655 19329 34667 19363
rect 34609 19323 34667 19329
rect 34793 19363 34851 19369
rect 34793 19329 34805 19363
rect 34839 19329 34851 19363
rect 34793 19323 34851 19329
rect 34885 19363 34943 19369
rect 34885 19329 34897 19363
rect 34931 19329 34943 19363
rect 34885 19323 34943 19329
rect 34977 19363 35035 19369
rect 34977 19329 34989 19363
rect 35023 19329 35035 19363
rect 35084 19360 35112 19456
rect 35161 19363 35219 19369
rect 35161 19360 35173 19363
rect 35084 19332 35173 19360
rect 34977 19323 35035 19329
rect 35161 19329 35173 19332
rect 35207 19329 35219 19363
rect 35161 19323 35219 19329
rect 32272 19264 32996 19292
rect 32272 19252 32278 19264
rect 32401 19227 32459 19233
rect 32401 19193 32413 19227
rect 32447 19224 32459 19227
rect 34514 19224 34520 19236
rect 32447 19196 34520 19224
rect 32447 19193 32459 19196
rect 32401 19187 32459 19193
rect 34514 19184 34520 19196
rect 34572 19184 34578 19236
rect 34808 19168 34836 19323
rect 34900 19292 34928 19323
rect 34900 19264 35388 19292
rect 35360 19236 35388 19264
rect 35342 19184 35348 19236
rect 35400 19184 35406 19236
rect 33318 19156 33324 19168
rect 31726 19128 33324 19156
rect 33318 19116 33324 19128
rect 33376 19116 33382 19168
rect 34790 19116 34796 19168
rect 34848 19156 34854 19168
rect 35069 19159 35127 19165
rect 35069 19156 35081 19159
rect 34848 19128 35081 19156
rect 34848 19116 34854 19128
rect 35069 19125 35081 19128
rect 35115 19156 35127 19159
rect 35710 19156 35716 19168
rect 35115 19128 35716 19156
rect 35115 19125 35127 19128
rect 35069 19119 35127 19125
rect 35710 19116 35716 19128
rect 35768 19116 35774 19168
rect 1104 19066 38272 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38272 19066
rect 1104 18992 38272 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 2004 18924 2329 18952
rect 2004 18912 2010 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 3786 18912 3792 18964
rect 3844 18912 3850 18964
rect 4614 18912 4620 18964
rect 4672 18952 4678 18964
rect 4801 18955 4859 18961
rect 4801 18952 4813 18955
rect 4672 18924 4813 18952
rect 4672 18912 4678 18924
rect 4801 18921 4813 18924
rect 4847 18921 4859 18955
rect 4801 18915 4859 18921
rect 7006 18912 7012 18964
rect 7064 18912 7070 18964
rect 8662 18912 8668 18964
rect 8720 18912 8726 18964
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10744 18924 11069 18952
rect 10744 18912 10750 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 11885 18955 11943 18961
rect 11885 18921 11897 18955
rect 11931 18952 11943 18955
rect 12158 18952 12164 18964
rect 11931 18924 12164 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 12526 18912 12532 18964
rect 12584 18912 12590 18964
rect 15289 18955 15347 18961
rect 15289 18952 15301 18955
rect 13004 18924 15301 18952
rect 7024 18884 7052 18912
rect 5920 18856 7052 18884
rect 3234 18816 3240 18828
rect 2148 18788 3240 18816
rect 1489 18751 1547 18757
rect 1489 18717 1501 18751
rect 1535 18748 1547 18751
rect 1762 18748 1768 18760
rect 1535 18720 1768 18748
rect 1535 18717 1547 18720
rect 1489 18711 1547 18717
rect 1762 18708 1768 18720
rect 1820 18708 1826 18760
rect 2038 18708 2044 18760
rect 2096 18708 2102 18760
rect 2148 18757 2176 18788
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 5920 18825 5948 18856
rect 8754 18844 8760 18896
rect 8812 18884 8818 18896
rect 10410 18884 10416 18896
rect 8812 18856 10416 18884
rect 8812 18844 8818 18856
rect 10410 18844 10416 18856
rect 10468 18844 10474 18896
rect 10962 18844 10968 18896
rect 11020 18844 11026 18896
rect 13004 18884 13032 18924
rect 15289 18921 15301 18924
rect 15335 18952 15347 18955
rect 17586 18952 17592 18964
rect 15335 18924 17592 18952
rect 15335 18921 15347 18924
rect 15289 18915 15347 18921
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 18138 18952 18144 18964
rect 17828 18924 18144 18952
rect 17828 18912 17834 18924
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 20073 18955 20131 18961
rect 20073 18952 20085 18955
rect 19484 18924 20085 18952
rect 19484 18912 19490 18924
rect 20073 18921 20085 18924
rect 20119 18921 20131 18955
rect 20073 18915 20131 18921
rect 20162 18912 20168 18964
rect 20220 18952 20226 18964
rect 20441 18955 20499 18961
rect 20441 18952 20453 18955
rect 20220 18924 20453 18952
rect 20220 18912 20226 18924
rect 20441 18921 20453 18924
rect 20487 18921 20499 18955
rect 20441 18915 20499 18921
rect 20622 18912 20628 18964
rect 20680 18912 20686 18964
rect 21910 18912 21916 18964
rect 21968 18912 21974 18964
rect 22480 18924 23152 18952
rect 12176 18856 13032 18884
rect 5905 18819 5963 18825
rect 4080 18788 5856 18816
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18717 2559 18751
rect 2501 18711 2559 18717
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18748 2651 18751
rect 3510 18748 3516 18760
rect 2639 18720 3516 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 2056 18680 2084 18708
rect 2516 18680 2544 18711
rect 3510 18708 3516 18720
rect 3568 18708 3574 18760
rect 4080 18757 4108 18788
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 4154 18708 4160 18760
rect 4212 18708 4218 18760
rect 4246 18708 4252 18760
rect 4304 18708 4310 18760
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18748 5043 18751
rect 5031 18720 5488 18748
rect 5031 18717 5043 18720
rect 4985 18711 5043 18717
rect 2958 18680 2964 18692
rect 2056 18652 2964 18680
rect 2958 18640 2964 18652
rect 3016 18680 3022 18692
rect 4448 18680 4476 18711
rect 5350 18680 5356 18692
rect 3016 18652 5356 18680
rect 3016 18640 3022 18652
rect 5350 18640 5356 18652
rect 5408 18640 5414 18692
rect 934 18572 940 18624
rect 992 18612 998 18624
rect 1581 18615 1639 18621
rect 1581 18612 1593 18615
rect 992 18584 1593 18612
rect 992 18572 998 18584
rect 1581 18581 1593 18584
rect 1627 18581 1639 18615
rect 1581 18575 1639 18581
rect 2774 18572 2780 18624
rect 2832 18572 2838 18624
rect 5460 18621 5488 18720
rect 5828 18680 5856 18788
rect 5905 18785 5917 18819
rect 5951 18785 5963 18819
rect 5905 18779 5963 18785
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 6914 18776 6920 18828
rect 6972 18816 6978 18828
rect 12176 18825 12204 18856
rect 13078 18844 13084 18896
rect 13136 18884 13142 18896
rect 22480 18884 22508 18924
rect 23124 18896 23152 18924
rect 23290 18912 23296 18964
rect 23348 18912 23354 18964
rect 23382 18912 23388 18964
rect 23440 18912 23446 18964
rect 23658 18912 23664 18964
rect 23716 18912 23722 18964
rect 23750 18912 23756 18964
rect 23808 18912 23814 18964
rect 23934 18912 23940 18964
rect 23992 18952 23998 18964
rect 24118 18952 24124 18964
rect 23992 18924 24124 18952
rect 23992 18912 23998 18924
rect 24118 18912 24124 18924
rect 24176 18912 24182 18964
rect 26786 18952 26792 18964
rect 24596 18924 26792 18952
rect 22922 18884 22928 18896
rect 13136 18856 22508 18884
rect 22572 18856 22928 18884
rect 13136 18844 13142 18856
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 6972 18788 9168 18816
rect 6972 18776 6978 18788
rect 9140 18760 9168 18788
rect 10336 18788 11161 18816
rect 8294 18708 8300 18760
rect 8352 18708 8358 18760
rect 9122 18708 9128 18760
rect 9180 18708 9186 18760
rect 10336 18757 10364 18788
rect 11149 18785 11161 18788
rect 11195 18816 11207 18819
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11195 18788 12173 18816
rect 11195 18785 11207 18788
rect 11149 18779 11207 18785
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 10594 18748 10600 18760
rect 10551 18720 10600 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 10873 18751 10931 18757
rect 10873 18750 10885 18751
rect 10796 18722 10885 18750
rect 7193 18683 7251 18689
rect 5828 18652 7144 18680
rect 5445 18615 5503 18621
rect 5445 18581 5457 18615
rect 5491 18581 5503 18615
rect 5445 18575 5503 18581
rect 5813 18615 5871 18621
rect 5813 18581 5825 18615
rect 5859 18612 5871 18615
rect 5994 18612 6000 18624
rect 5859 18584 6000 18612
rect 5859 18581 5871 18584
rect 5813 18575 5871 18581
rect 5994 18572 6000 18584
rect 6052 18612 6058 18624
rect 6914 18612 6920 18624
rect 6052 18584 6920 18612
rect 6052 18572 6058 18584
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7116 18612 7144 18652
rect 7193 18649 7205 18683
rect 7239 18680 7251 18683
rect 7466 18680 7472 18692
rect 7239 18652 7472 18680
rect 7239 18649 7251 18652
rect 7193 18643 7251 18649
rect 7466 18640 7472 18652
rect 7524 18640 7530 18692
rect 10134 18680 10140 18692
rect 9646 18652 10140 18680
rect 9646 18612 9674 18652
rect 10134 18640 10140 18652
rect 10192 18680 10198 18692
rect 10796 18680 10824 18722
rect 10873 18717 10885 18722
rect 10919 18717 10931 18751
rect 10873 18711 10931 18717
rect 10962 18708 10968 18760
rect 11020 18748 11026 18760
rect 11440 18757 11468 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 16574 18816 16580 18828
rect 15672 18788 16580 18816
rect 13725 18761 13783 18767
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 11020 18720 11345 18748
rect 11020 18708 11026 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 11790 18708 11796 18760
rect 11848 18708 11854 18760
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 13078 18708 13084 18760
rect 13136 18748 13142 18760
rect 13438 18751 13496 18757
rect 13438 18750 13450 18751
rect 13188 18748 13450 18750
rect 13136 18722 13450 18748
rect 13136 18720 13216 18722
rect 13136 18708 13142 18720
rect 13438 18717 13450 18722
rect 13484 18717 13496 18751
rect 13725 18727 13737 18761
rect 13771 18727 13783 18761
rect 15672 18760 15700 18788
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17037 18819 17095 18825
rect 17037 18816 17049 18819
rect 16816 18788 17049 18816
rect 16816 18776 16822 18788
rect 17037 18785 17049 18788
rect 17083 18785 17095 18819
rect 17037 18779 17095 18785
rect 18138 18776 18144 18828
rect 18196 18816 18202 18828
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 18196 18788 19073 18816
rect 18196 18776 18202 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19797 18819 19855 18825
rect 19797 18816 19809 18819
rect 19061 18779 19119 18785
rect 19168 18788 19809 18816
rect 13725 18721 13783 18727
rect 13438 18711 13496 18717
rect 13740 18692 13768 18721
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 13872 18720 14105 18748
rect 13872 18708 13878 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 15197 18751 15255 18757
rect 15197 18717 15209 18751
rect 15243 18717 15255 18751
rect 15197 18711 15255 18717
rect 10192 18652 10732 18680
rect 10796 18652 12112 18680
rect 10192 18640 10198 18652
rect 7116 18584 9674 18612
rect 10410 18572 10416 18624
rect 10468 18572 10474 18624
rect 10594 18572 10600 18624
rect 10652 18572 10658 18624
rect 10704 18612 10732 18652
rect 11974 18612 11980 18624
rect 10704 18584 11980 18612
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12084 18621 12112 18652
rect 12802 18640 12808 18692
rect 12860 18640 12866 18692
rect 12986 18640 12992 18692
rect 13044 18640 13050 18692
rect 13262 18640 13268 18692
rect 13320 18640 13326 18692
rect 13722 18640 13728 18692
rect 13780 18680 13786 18692
rect 14366 18680 14372 18692
rect 13780 18652 14372 18680
rect 13780 18640 13786 18652
rect 14366 18640 14372 18652
rect 14424 18640 14430 18692
rect 14918 18640 14924 18692
rect 14976 18640 14982 18692
rect 15212 18680 15240 18711
rect 15378 18708 15384 18760
rect 15436 18708 15442 18760
rect 15654 18708 15660 18760
rect 15712 18708 15718 18760
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 16255 18720 16344 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 16022 18680 16028 18692
rect 15212 18652 16028 18680
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 12069 18615 12127 18621
rect 12069 18581 12081 18615
rect 12115 18581 12127 18615
rect 12069 18575 12127 18581
rect 12526 18572 12532 18624
rect 12584 18572 12590 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 13173 18615 13231 18621
rect 13173 18612 13185 18615
rect 13136 18584 13185 18612
rect 13136 18572 13142 18584
rect 13173 18581 13185 18584
rect 13219 18581 13231 18615
rect 13173 18575 13231 18581
rect 13630 18572 13636 18624
rect 13688 18612 13694 18624
rect 13817 18615 13875 18621
rect 13817 18612 13829 18615
rect 13688 18584 13829 18612
rect 13688 18572 13694 18584
rect 13817 18581 13829 18584
rect 13863 18612 13875 18615
rect 16316 18612 16344 18720
rect 16482 18708 16488 18760
rect 16540 18708 16546 18760
rect 16850 18708 16856 18760
rect 16908 18708 16914 18760
rect 17126 18708 17132 18760
rect 17184 18708 17190 18760
rect 17494 18708 17500 18760
rect 17552 18708 17558 18760
rect 17586 18708 17592 18760
rect 17644 18748 17650 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 17644 18720 18521 18748
rect 17644 18708 17650 18720
rect 18509 18717 18521 18720
rect 18555 18748 18567 18751
rect 19168 18748 19196 18788
rect 19797 18785 19809 18788
rect 19843 18785 19855 18819
rect 19797 18779 19855 18785
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18816 19947 18819
rect 20530 18816 20536 18828
rect 19935 18788 20536 18816
rect 19935 18785 19947 18788
rect 19889 18779 19947 18785
rect 18555 18720 19196 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19812 18748 19840 18779
rect 20530 18776 20536 18788
rect 20588 18776 20594 18828
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 22005 18819 22063 18825
rect 22005 18816 22017 18819
rect 21876 18788 22017 18816
rect 21876 18776 21882 18788
rect 22005 18785 22017 18788
rect 22051 18785 22063 18819
rect 22005 18779 22063 18785
rect 22462 18776 22468 18828
rect 22520 18776 22526 18828
rect 20806 18748 20812 18760
rect 19300 18720 19472 18748
rect 19812 18720 20812 18748
rect 19300 18708 19306 18720
rect 17862 18640 17868 18692
rect 17920 18680 17926 18692
rect 18046 18680 18052 18692
rect 17920 18652 18052 18680
rect 17920 18640 17926 18652
rect 18046 18640 18052 18652
rect 18104 18640 18110 18692
rect 18141 18683 18199 18689
rect 18141 18649 18153 18683
rect 18187 18649 18199 18683
rect 18141 18643 18199 18649
rect 13863 18584 16344 18612
rect 18156 18612 18184 18643
rect 18322 18640 18328 18692
rect 18380 18680 18386 18692
rect 18601 18683 18659 18689
rect 18601 18680 18613 18683
rect 18380 18652 18613 18680
rect 18380 18640 18386 18652
rect 18601 18649 18613 18652
rect 18647 18649 18659 18683
rect 18601 18643 18659 18649
rect 19058 18640 19064 18692
rect 19116 18640 19122 18692
rect 19076 18612 19104 18640
rect 19444 18621 19472 18720
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 22186 18708 22192 18760
rect 22244 18708 22250 18760
rect 22572 18748 22600 18856
rect 22922 18844 22928 18856
rect 22980 18844 22986 18896
rect 23106 18844 23112 18896
rect 23164 18844 23170 18896
rect 23308 18884 23336 18912
rect 24394 18884 24400 18896
rect 23308 18856 24400 18884
rect 24394 18844 24400 18856
rect 24452 18844 24458 18896
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 23198 18816 23204 18828
rect 23072 18788 23204 18816
rect 23072 18776 23078 18788
rect 23198 18776 23204 18788
rect 23256 18816 23262 18828
rect 23293 18819 23351 18825
rect 23293 18816 23305 18819
rect 23256 18788 23305 18816
rect 23256 18776 23262 18788
rect 23293 18785 23305 18788
rect 23339 18785 23351 18819
rect 23293 18779 23351 18785
rect 23842 18776 23848 18828
rect 23900 18816 23906 18828
rect 23900 18788 24164 18816
rect 23900 18776 23906 18788
rect 24136 18760 24164 18788
rect 24210 18776 24216 18828
rect 24268 18825 24274 18828
rect 24268 18816 24277 18825
rect 24596 18816 24624 18924
rect 26786 18912 26792 18924
rect 26844 18912 26850 18964
rect 28718 18912 28724 18964
rect 28776 18912 28782 18964
rect 32953 18955 33011 18961
rect 32953 18952 32965 18955
rect 28966 18924 32965 18952
rect 26697 18887 26755 18893
rect 26697 18853 26709 18887
rect 26743 18853 26755 18887
rect 26804 18884 26832 18912
rect 28966 18884 28994 18924
rect 32953 18921 32965 18924
rect 32999 18921 33011 18955
rect 32953 18915 33011 18921
rect 26804 18856 28994 18884
rect 26697 18847 26755 18853
rect 24268 18788 24624 18816
rect 24268 18779 24277 18788
rect 24268 18776 24274 18779
rect 24762 18776 24768 18828
rect 24820 18816 24826 18828
rect 26602 18816 26608 18828
rect 24820 18788 26608 18816
rect 24820 18776 24826 18788
rect 22741 18751 22799 18757
rect 22741 18748 22753 18751
rect 22572 18720 22753 18748
rect 22741 18717 22753 18720
rect 22787 18717 22799 18751
rect 22741 18711 22799 18717
rect 22830 18708 22836 18760
rect 22888 18708 22894 18760
rect 22922 18708 22928 18760
rect 22980 18708 22986 18760
rect 23109 18751 23167 18757
rect 23109 18717 23121 18751
rect 23155 18748 23167 18751
rect 23155 18720 23336 18748
rect 23155 18717 23167 18720
rect 23109 18711 23167 18717
rect 20070 18640 20076 18692
rect 20128 18680 20134 18692
rect 20257 18683 20315 18689
rect 20257 18680 20269 18683
rect 20128 18652 20269 18680
rect 20128 18640 20134 18652
rect 20257 18649 20269 18652
rect 20303 18649 20315 18683
rect 20257 18643 20315 18649
rect 20364 18652 21312 18680
rect 18156 18584 19104 18612
rect 19429 18615 19487 18621
rect 13863 18581 13875 18584
rect 13817 18575 13875 18581
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 20364 18612 20392 18652
rect 21284 18624 21312 18652
rect 21358 18640 21364 18692
rect 21416 18680 21422 18692
rect 21913 18683 21971 18689
rect 21913 18680 21925 18683
rect 21416 18652 21925 18680
rect 21416 18640 21422 18652
rect 21913 18649 21925 18652
rect 21959 18649 21971 18683
rect 23201 18683 23259 18689
rect 23201 18680 23213 18683
rect 21913 18643 21971 18649
rect 22388 18652 23213 18680
rect 19475 18584 20392 18612
rect 20467 18615 20525 18621
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 20467 18581 20479 18615
rect 20513 18612 20525 18615
rect 20622 18612 20628 18624
rect 20513 18584 20628 18612
rect 20513 18581 20525 18584
rect 20467 18575 20525 18581
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 21266 18572 21272 18624
rect 21324 18572 21330 18624
rect 22388 18621 22416 18652
rect 23201 18649 23213 18652
rect 23247 18649 23259 18683
rect 23201 18643 23259 18649
rect 22373 18615 22431 18621
rect 22373 18581 22385 18615
rect 22419 18581 22431 18615
rect 22373 18575 22431 18581
rect 22462 18572 22468 18624
rect 22520 18612 22526 18624
rect 23308 18612 23336 18720
rect 23382 18708 23388 18760
rect 23440 18748 23446 18760
rect 23477 18751 23535 18757
rect 23477 18748 23489 18751
rect 23440 18720 23489 18748
rect 23440 18708 23446 18720
rect 23477 18717 23489 18720
rect 23523 18717 23535 18751
rect 23477 18711 23535 18717
rect 23937 18751 23995 18757
rect 23937 18717 23949 18751
rect 23983 18748 23995 18751
rect 24026 18748 24032 18760
rect 23983 18720 24032 18748
rect 23983 18717 23995 18720
rect 23937 18711 23995 18717
rect 24026 18708 24032 18720
rect 24084 18708 24090 18760
rect 24118 18708 24124 18760
rect 24176 18708 24182 18760
rect 25038 18708 25044 18760
rect 25096 18748 25102 18760
rect 25317 18751 25375 18757
rect 25317 18748 25329 18751
rect 25096 18720 25329 18748
rect 25096 18708 25102 18720
rect 25317 18717 25329 18720
rect 25363 18717 25375 18751
rect 25317 18711 25375 18717
rect 25685 18751 25743 18757
rect 25685 18717 25697 18751
rect 25731 18748 25743 18751
rect 25774 18748 25780 18760
rect 25731 18720 25780 18748
rect 25731 18717 25743 18720
rect 25685 18711 25743 18717
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 25884 18757 25912 18788
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 26712 18816 26740 18847
rect 31754 18844 31760 18896
rect 31812 18884 31818 18896
rect 31849 18887 31907 18893
rect 31849 18884 31861 18887
rect 31812 18856 31861 18884
rect 31812 18844 31818 18856
rect 31849 18853 31861 18856
rect 31895 18853 31907 18887
rect 31849 18847 31907 18853
rect 32309 18887 32367 18893
rect 32309 18853 32321 18887
rect 32355 18853 32367 18887
rect 32309 18847 32367 18853
rect 31113 18819 31171 18825
rect 26712 18788 31064 18816
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 26142 18708 26148 18760
rect 26200 18708 26206 18760
rect 26513 18751 26571 18757
rect 26513 18717 26525 18751
rect 26559 18717 26571 18751
rect 26513 18711 26571 18717
rect 28629 18751 28687 18757
rect 28629 18717 28641 18751
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 24854 18640 24860 18692
rect 24912 18680 24918 18692
rect 25590 18680 25596 18692
rect 24912 18652 25596 18680
rect 24912 18640 24918 18652
rect 25590 18640 25596 18652
rect 25648 18680 25654 18692
rect 26329 18683 26387 18689
rect 26329 18680 26341 18683
rect 25648 18652 26341 18680
rect 25648 18640 25654 18652
rect 26329 18649 26341 18652
rect 26375 18649 26387 18683
rect 26329 18643 26387 18649
rect 26418 18640 26424 18692
rect 26476 18640 26482 18692
rect 22520 18584 23336 18612
rect 22520 18572 22526 18584
rect 25866 18572 25872 18624
rect 25924 18612 25930 18624
rect 26528 18612 26556 18711
rect 28644 18680 28672 18711
rect 28810 18708 28816 18760
rect 28868 18708 28874 18760
rect 29178 18708 29184 18760
rect 29236 18708 29242 18760
rect 31036 18757 31064 18788
rect 31113 18785 31125 18819
rect 31159 18816 31171 18819
rect 32324 18816 32352 18847
rect 34698 18844 34704 18896
rect 34756 18884 34762 18896
rect 34756 18856 35112 18884
rect 34756 18844 34762 18856
rect 31159 18788 32076 18816
rect 32324 18788 33732 18816
rect 31159 18785 31171 18788
rect 31113 18779 31171 18785
rect 31021 18751 31079 18757
rect 31021 18717 31033 18751
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 29196 18680 29224 18708
rect 28644 18652 29224 18680
rect 31036 18680 31064 18711
rect 31202 18708 31208 18760
rect 31260 18748 31266 18760
rect 32048 18757 32076 18788
rect 31481 18751 31539 18757
rect 31481 18748 31493 18751
rect 31260 18720 31493 18748
rect 31260 18708 31266 18720
rect 31481 18717 31493 18720
rect 31527 18717 31539 18751
rect 31481 18711 31539 18717
rect 31665 18751 31723 18757
rect 31665 18717 31677 18751
rect 31711 18748 31723 18751
rect 31757 18751 31815 18757
rect 31757 18748 31769 18751
rect 31711 18720 31769 18748
rect 31711 18717 31723 18720
rect 31665 18711 31723 18717
rect 31757 18717 31769 18720
rect 31803 18717 31815 18751
rect 31757 18711 31815 18717
rect 32033 18751 32091 18757
rect 32033 18717 32045 18751
rect 32079 18717 32091 18751
rect 32033 18711 32091 18717
rect 31297 18683 31355 18689
rect 31297 18680 31309 18683
rect 31036 18652 31309 18680
rect 31297 18649 31309 18652
rect 31343 18649 31355 18683
rect 31938 18680 31944 18692
rect 31297 18643 31355 18649
rect 31726 18652 31944 18680
rect 25924 18584 26556 18612
rect 31312 18612 31340 18643
rect 31726 18612 31754 18652
rect 31938 18640 31944 18652
rect 31996 18640 32002 18692
rect 32048 18624 32076 18711
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32309 18751 32367 18757
rect 32309 18748 32321 18751
rect 32272 18720 32321 18748
rect 32272 18708 32278 18720
rect 32309 18717 32321 18720
rect 32355 18717 32367 18751
rect 32309 18711 32367 18717
rect 32582 18708 32588 18760
rect 32640 18708 32646 18760
rect 32861 18751 32919 18757
rect 32861 18748 32873 18751
rect 32784 18720 32873 18748
rect 32600 18680 32628 18708
rect 32324 18652 32628 18680
rect 32324 18624 32352 18652
rect 32784 18624 32812 18720
rect 32861 18717 32873 18720
rect 32907 18717 32919 18751
rect 32861 18711 32919 18717
rect 32950 18640 32956 18692
rect 33008 18680 33014 18692
rect 33704 18680 33732 18788
rect 35084 18748 35112 18856
rect 35526 18844 35532 18896
rect 35584 18844 35590 18896
rect 35158 18776 35164 18828
rect 35216 18776 35222 18828
rect 35345 18819 35403 18825
rect 35345 18785 35357 18819
rect 35391 18816 35403 18819
rect 35434 18816 35440 18828
rect 35391 18788 35440 18816
rect 35391 18785 35403 18788
rect 35345 18779 35403 18785
rect 35434 18776 35440 18788
rect 35492 18776 35498 18828
rect 35805 18751 35863 18757
rect 35805 18748 35817 18751
rect 35084 18720 35817 18748
rect 35805 18717 35817 18720
rect 35851 18717 35863 18751
rect 35805 18711 35863 18717
rect 35069 18683 35127 18689
rect 35069 18680 35081 18683
rect 33008 18652 33640 18680
rect 33704 18652 35081 18680
rect 33008 18640 33014 18652
rect 31312 18584 31754 18612
rect 25924 18572 25930 18584
rect 32030 18572 32036 18624
rect 32088 18572 32094 18624
rect 32306 18572 32312 18624
rect 32364 18572 32370 18624
rect 32398 18572 32404 18624
rect 32456 18612 32462 18624
rect 32493 18615 32551 18621
rect 32493 18612 32505 18615
rect 32456 18584 32505 18612
rect 32456 18572 32462 18584
rect 32493 18581 32505 18584
rect 32539 18581 32551 18615
rect 32493 18575 32551 18581
rect 32766 18572 32772 18624
rect 32824 18572 32830 18624
rect 33612 18612 33640 18652
rect 35069 18649 35081 18652
rect 35115 18649 35127 18683
rect 35069 18643 35127 18649
rect 35529 18683 35587 18689
rect 35529 18649 35541 18683
rect 35575 18649 35587 18683
rect 35529 18643 35587 18649
rect 35544 18612 35572 18643
rect 35710 18640 35716 18692
rect 35768 18640 35774 18692
rect 36262 18612 36268 18624
rect 33612 18584 36268 18612
rect 36262 18572 36268 18584
rect 36320 18572 36326 18624
rect 1104 18522 38272 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38272 18522
rect 1104 18448 38272 18470
rect 2406 18368 2412 18420
rect 2464 18368 2470 18420
rect 2774 18408 2780 18420
rect 2746 18368 2780 18408
rect 2832 18368 2838 18420
rect 3510 18368 3516 18420
rect 3568 18368 3574 18420
rect 3605 18411 3663 18417
rect 3605 18377 3617 18411
rect 3651 18408 3663 18411
rect 4246 18408 4252 18420
rect 3651 18380 4252 18408
rect 3651 18377 3663 18380
rect 3605 18371 3663 18377
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 4540 18380 6377 18408
rect 2424 18340 2452 18368
rect 1780 18312 2452 18340
rect 1780 18281 1808 18312
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2746 18272 2774 18368
rect 3528 18340 3556 18368
rect 4540 18340 4568 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 6472 18380 7052 18408
rect 3528 18312 4568 18340
rect 2179 18244 2774 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 3234 18232 3240 18284
rect 3292 18232 3298 18284
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18272 3479 18275
rect 4062 18272 4068 18284
rect 3467 18244 4068 18272
rect 3467 18241 3479 18244
rect 3421 18235 3479 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 6472 18272 6500 18380
rect 6914 18300 6920 18352
rect 6972 18300 6978 18352
rect 7024 18349 7052 18380
rect 9122 18368 9128 18420
rect 9180 18368 9186 18420
rect 10594 18408 10600 18420
rect 10520 18380 10600 18408
rect 7009 18343 7067 18349
rect 7009 18309 7021 18343
rect 7055 18340 7067 18343
rect 8754 18340 8760 18352
rect 7055 18312 8760 18340
rect 7055 18309 7067 18312
rect 7009 18303 7067 18309
rect 8754 18300 8760 18312
rect 8812 18300 8818 18352
rect 10520 18349 10548 18380
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 10689 18411 10747 18417
rect 10689 18377 10701 18411
rect 10735 18377 10747 18411
rect 10689 18371 10747 18377
rect 12069 18411 12127 18417
rect 12069 18377 12081 18411
rect 12115 18408 12127 18411
rect 12710 18408 12716 18420
rect 12115 18380 12716 18408
rect 12115 18377 12127 18380
rect 12069 18371 12127 18377
rect 10505 18343 10563 18349
rect 10505 18309 10517 18343
rect 10551 18309 10563 18343
rect 10704 18340 10732 18371
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 15562 18368 15568 18420
rect 15620 18408 15626 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15620 18380 15669 18408
rect 15620 18368 15626 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15657 18371 15715 18377
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 16298 18408 16304 18420
rect 16080 18380 16304 18408
rect 16080 18368 16086 18380
rect 16298 18368 16304 18380
rect 16356 18368 16362 18420
rect 16482 18368 16488 18420
rect 16540 18408 16546 18420
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 16540 18380 16865 18408
rect 16540 18368 16546 18380
rect 16853 18377 16865 18380
rect 16899 18408 16911 18411
rect 17126 18408 17132 18420
rect 16899 18380 17132 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 18690 18368 18696 18420
rect 18748 18368 18754 18420
rect 19429 18411 19487 18417
rect 19429 18377 19441 18411
rect 19475 18408 19487 18411
rect 20714 18408 20720 18420
rect 19475 18380 20720 18408
rect 19475 18377 19487 18380
rect 19429 18371 19487 18377
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 25130 18408 25136 18420
rect 21876 18380 25136 18408
rect 21876 18368 21882 18380
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 25314 18368 25320 18420
rect 25372 18408 25378 18420
rect 25372 18380 31754 18408
rect 25372 18368 25378 18380
rect 11977 18343 12035 18349
rect 11977 18340 11989 18343
rect 10704 18312 11989 18340
rect 10505 18303 10563 18309
rect 11977 18309 11989 18312
rect 12023 18309 12035 18343
rect 19702 18340 19708 18352
rect 11977 18303 12035 18309
rect 12084 18312 19708 18340
rect 4212 18244 6500 18272
rect 6641 18275 6699 18281
rect 4212 18232 4218 18244
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 6822 18273 6828 18284
rect 6748 18272 6828 18273
rect 6687 18245 6828 18272
rect 6687 18244 6776 18245
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 6822 18232 6828 18245
rect 6880 18232 6886 18284
rect 7101 18275 7159 18281
rect 7101 18241 7113 18275
rect 7147 18272 7159 18275
rect 7190 18272 7196 18284
rect 7147 18244 7196 18272
rect 7147 18241 7159 18244
rect 7101 18235 7159 18241
rect 7190 18232 7196 18244
rect 7248 18272 7254 18284
rect 7837 18275 7895 18281
rect 7248 18244 7420 18272
rect 7248 18232 7254 18244
rect 3252 18204 3280 18232
rect 3878 18204 3884 18216
rect 3252 18176 3884 18204
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 6534 18207 6592 18213
rect 6534 18173 6546 18207
rect 6580 18204 6592 18207
rect 6580 18176 6684 18204
rect 6580 18173 6592 18176
rect 6534 18167 6592 18173
rect 1946 18028 1952 18080
rect 2004 18028 2010 18080
rect 2314 18028 2320 18080
rect 2372 18028 2378 18080
rect 6656 18068 6684 18176
rect 6730 18164 6736 18216
rect 6788 18204 6794 18216
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6788 18176 7297 18204
rect 6788 18164 6794 18176
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 7392 18136 7420 18244
rect 7837 18241 7849 18275
rect 7883 18272 7895 18275
rect 8570 18272 8576 18284
rect 7883 18244 8576 18272
rect 7883 18241 7895 18244
rect 7837 18235 7895 18241
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 9030 18232 9036 18284
rect 9088 18272 9094 18284
rect 9582 18272 9588 18284
rect 9088 18244 9588 18272
rect 9088 18232 9094 18244
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 10134 18232 10140 18284
rect 10192 18232 10198 18284
rect 10686 18232 10692 18284
rect 10744 18232 10750 18284
rect 10962 18232 10968 18284
rect 11020 18232 11026 18284
rect 11057 18275 11115 18281
rect 11057 18241 11069 18275
rect 11103 18241 11115 18275
rect 11057 18235 11115 18241
rect 11170 18278 11228 18284
rect 11170 18244 11182 18278
rect 11216 18275 11228 18278
rect 11216 18272 11284 18275
rect 11216 18247 11290 18272
rect 11216 18244 11228 18247
rect 11256 18244 11290 18247
rect 11170 18238 11228 18244
rect 10321 18207 10379 18213
rect 10321 18173 10333 18207
rect 10367 18204 10379 18207
rect 10410 18204 10416 18216
rect 10367 18176 10416 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 10410 18164 10416 18176
rect 10468 18204 10474 18216
rect 10594 18204 10600 18216
rect 10468 18176 10600 18204
rect 10468 18164 10474 18176
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 10704 18204 10732 18232
rect 11072 18204 11100 18235
rect 10704 18176 11100 18204
rect 11262 18204 11290 18244
rect 11330 18232 11336 18284
rect 11388 18232 11394 18284
rect 11790 18232 11796 18284
rect 11848 18232 11854 18284
rect 12084 18272 12112 18312
rect 19702 18300 19708 18312
rect 19760 18300 19766 18352
rect 20533 18343 20591 18349
rect 20533 18309 20545 18343
rect 20579 18340 20591 18343
rect 20898 18340 20904 18352
rect 20579 18312 20904 18340
rect 20579 18309 20591 18312
rect 20533 18303 20591 18309
rect 20898 18300 20904 18312
rect 20956 18300 20962 18352
rect 21910 18300 21916 18352
rect 21968 18340 21974 18352
rect 23842 18340 23848 18352
rect 21968 18312 23848 18340
rect 21968 18300 21974 18312
rect 23842 18300 23848 18312
rect 23900 18340 23906 18352
rect 24486 18340 24492 18352
rect 23900 18312 24492 18340
rect 23900 18300 23906 18312
rect 24486 18300 24492 18312
rect 24544 18300 24550 18352
rect 28350 18300 28356 18352
rect 28408 18340 28414 18352
rect 31726 18340 31754 18380
rect 32030 18368 32036 18420
rect 32088 18408 32094 18420
rect 32125 18411 32183 18417
rect 32125 18408 32137 18411
rect 32088 18380 32137 18408
rect 32088 18368 32094 18380
rect 32125 18377 32137 18380
rect 32171 18377 32183 18411
rect 32125 18371 32183 18377
rect 32769 18411 32827 18417
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 35158 18408 35164 18420
rect 32815 18380 35164 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 35158 18368 35164 18380
rect 35216 18368 35222 18420
rect 35526 18368 35532 18420
rect 35584 18368 35590 18420
rect 35069 18343 35127 18349
rect 28408 18312 28948 18340
rect 31726 18312 34836 18340
rect 28408 18300 28414 18312
rect 11992 18244 12112 18272
rect 11808 18204 11836 18232
rect 11992 18216 12020 18244
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 13630 18272 13636 18284
rect 12584 18244 13636 18272
rect 12584 18232 12590 18244
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 11262 18176 11836 18204
rect 11974 18164 11980 18216
rect 12032 18164 12038 18216
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12161 18207 12219 18213
rect 12161 18204 12173 18207
rect 12124 18176 12173 18204
rect 12124 18164 12130 18176
rect 12161 18173 12173 18176
rect 12207 18173 12219 18207
rect 12161 18167 12219 18173
rect 13078 18164 13084 18216
rect 13136 18204 13142 18216
rect 13814 18204 13820 18216
rect 13136 18176 13820 18204
rect 13136 18164 13142 18176
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 15580 18204 15608 18235
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18272 15899 18275
rect 15930 18272 15936 18284
rect 15887 18244 15936 18272
rect 15887 18241 15899 18244
rect 15841 18235 15899 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18272 16083 18275
rect 16114 18272 16120 18284
rect 16071 18244 16120 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 16114 18232 16120 18244
rect 16172 18272 16178 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 16172 18244 17049 18272
rect 16172 18232 16178 18244
rect 17037 18241 17049 18244
rect 17083 18272 17095 18275
rect 17586 18272 17592 18284
rect 17083 18244 17592 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 18141 18275 18199 18281
rect 18141 18272 18153 18275
rect 17696 18244 18153 18272
rect 16482 18204 16488 18216
rect 15580 18176 16488 18204
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16669 18207 16727 18213
rect 16669 18204 16681 18207
rect 16632 18176 16681 18204
rect 16632 18164 16638 18176
rect 16669 18173 16681 18176
rect 16715 18173 16727 18207
rect 16669 18167 16727 18173
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17494 18204 17500 18216
rect 16816 18176 17500 18204
rect 16816 18164 16822 18176
rect 17494 18164 17500 18176
rect 17552 18204 17558 18216
rect 17696 18204 17724 18244
rect 18141 18241 18153 18244
rect 18187 18241 18199 18275
rect 18141 18235 18199 18241
rect 18506 18232 18512 18284
rect 18564 18232 18570 18284
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 18966 18272 18972 18284
rect 18656 18244 18972 18272
rect 18656 18232 18662 18244
rect 18966 18232 18972 18244
rect 19024 18272 19030 18284
rect 19061 18275 19119 18281
rect 19061 18272 19073 18275
rect 19024 18244 19073 18272
rect 19024 18232 19030 18244
rect 19061 18241 19073 18244
rect 19107 18241 19119 18275
rect 19061 18235 19119 18241
rect 19242 18232 19248 18284
rect 19300 18232 19306 18284
rect 20070 18232 20076 18284
rect 20128 18272 20134 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 20128 18244 20177 18272
rect 20128 18232 20134 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20349 18275 20407 18281
rect 20349 18272 20361 18275
rect 20312 18244 20361 18272
rect 20312 18232 20318 18244
rect 20349 18241 20361 18244
rect 20395 18272 20407 18275
rect 20806 18272 20812 18284
rect 20395 18244 20812 18272
rect 20395 18241 20407 18244
rect 20349 18235 20407 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 17552 18176 17724 18204
rect 17552 18164 17558 18176
rect 18046 18164 18052 18216
rect 18104 18164 18110 18216
rect 18414 18164 18420 18216
rect 18472 18204 18478 18216
rect 20916 18204 20944 18300
rect 23382 18232 23388 18284
rect 23440 18272 23446 18284
rect 27154 18272 27160 18284
rect 23440 18244 27160 18272
rect 23440 18232 23446 18244
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 28920 18281 28948 18312
rect 28537 18275 28595 18281
rect 28537 18241 28549 18275
rect 28583 18241 28595 18275
rect 28537 18235 28595 18241
rect 28905 18275 28963 18281
rect 28905 18241 28917 18275
rect 28951 18241 28963 18275
rect 28905 18235 28963 18241
rect 18472 18176 20944 18204
rect 18472 18164 18478 18176
rect 22186 18164 22192 18216
rect 22244 18204 22250 18216
rect 26694 18204 26700 18216
rect 22244 18176 26700 18204
rect 22244 18164 22250 18176
rect 26694 18164 26700 18176
rect 26752 18204 26758 18216
rect 27706 18204 27712 18216
rect 26752 18176 27712 18204
rect 26752 18164 26758 18176
rect 27706 18164 27712 18176
rect 27764 18164 27770 18216
rect 28350 18164 28356 18216
rect 28408 18164 28414 18216
rect 28552 18204 28580 18235
rect 30190 18232 30196 18284
rect 30248 18272 30254 18284
rect 32585 18275 32643 18281
rect 32585 18272 32597 18275
rect 30248 18244 32597 18272
rect 30248 18232 30254 18244
rect 32585 18241 32597 18244
rect 32631 18241 32643 18275
rect 32585 18235 32643 18241
rect 32861 18275 32919 18281
rect 32861 18241 32873 18275
rect 32907 18272 32919 18275
rect 32907 18244 33088 18272
rect 32907 18241 32919 18244
rect 32861 18235 32919 18241
rect 30098 18204 30104 18216
rect 28552 18176 30104 18204
rect 30098 18164 30104 18176
rect 30156 18164 30162 18216
rect 31110 18164 31116 18216
rect 31168 18164 31174 18216
rect 31754 18164 31760 18216
rect 31812 18204 31818 18216
rect 32398 18204 32404 18216
rect 31812 18176 32404 18204
rect 31812 18164 31818 18176
rect 32398 18164 32404 18176
rect 32456 18164 32462 18216
rect 32493 18207 32551 18213
rect 32493 18173 32505 18207
rect 32539 18204 32551 18207
rect 32953 18207 33011 18213
rect 32953 18204 32965 18207
rect 32539 18176 32965 18204
rect 32539 18173 32551 18176
rect 32493 18167 32551 18173
rect 32953 18173 32965 18176
rect 32999 18173 33011 18207
rect 32953 18167 33011 18173
rect 9582 18136 9588 18148
rect 7392 18108 9588 18136
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 10137 18139 10195 18145
rect 10137 18136 10149 18139
rect 9732 18108 10149 18136
rect 9732 18096 9738 18108
rect 10137 18105 10149 18108
rect 10183 18105 10195 18139
rect 10137 18099 10195 18105
rect 11054 18096 11060 18148
rect 11112 18136 11118 18148
rect 11609 18139 11667 18145
rect 11609 18136 11621 18139
rect 11112 18108 11621 18136
rect 11112 18096 11118 18108
rect 11609 18105 11621 18108
rect 11655 18105 11667 18139
rect 12986 18136 12992 18148
rect 11609 18099 11667 18105
rect 11808 18108 12992 18136
rect 11808 18068 11836 18108
rect 12986 18096 12992 18108
rect 13044 18096 13050 18148
rect 15562 18096 15568 18148
rect 15620 18136 15626 18148
rect 28813 18139 28871 18145
rect 28813 18136 28825 18139
rect 15620 18108 28825 18136
rect 15620 18096 15626 18108
rect 28813 18105 28825 18108
rect 28859 18105 28871 18139
rect 31128 18136 31156 18164
rect 32214 18136 32220 18148
rect 31128 18108 32220 18136
rect 28813 18099 28871 18105
rect 32214 18096 32220 18108
rect 32272 18096 32278 18148
rect 32416 18136 32444 18164
rect 33060 18136 33088 18244
rect 34698 18232 34704 18284
rect 34756 18232 34762 18284
rect 34808 18272 34836 18312
rect 35069 18309 35081 18343
rect 35115 18340 35127 18343
rect 35544 18340 35572 18368
rect 35115 18312 35572 18340
rect 35115 18309 35127 18312
rect 35069 18303 35127 18309
rect 37553 18275 37611 18281
rect 37553 18272 37565 18275
rect 34808 18244 37565 18272
rect 37553 18241 37565 18244
rect 37599 18241 37611 18275
rect 37553 18235 37611 18241
rect 34790 18164 34796 18216
rect 34848 18164 34854 18216
rect 32416 18108 33088 18136
rect 33410 18096 33416 18148
rect 33468 18136 33474 18148
rect 34701 18139 34759 18145
rect 34701 18136 34713 18139
rect 33468 18108 34713 18136
rect 33468 18096 33474 18108
rect 34701 18105 34713 18108
rect 34747 18105 34759 18139
rect 34701 18099 34759 18105
rect 6656 18040 11836 18068
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 13722 18068 13728 18080
rect 11940 18040 13728 18068
rect 11940 18028 11946 18040
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 15746 18028 15752 18080
rect 15804 18068 15810 18080
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 15804 18040 15945 18068
rect 15804 18028 15810 18040
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 17126 18068 17132 18080
rect 16356 18040 17132 18068
rect 16356 18028 16362 18040
rect 17126 18028 17132 18040
rect 17184 18068 17190 18080
rect 17221 18071 17279 18077
rect 17221 18068 17233 18071
rect 17184 18040 17233 18068
rect 17184 18028 17190 18040
rect 17221 18037 17233 18040
rect 17267 18068 17279 18071
rect 17862 18068 17868 18080
rect 17267 18040 17868 18068
rect 17267 18037 17279 18040
rect 17221 18031 17279 18037
rect 17862 18028 17868 18040
rect 17920 18068 17926 18080
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 17920 18040 18521 18068
rect 17920 18028 17926 18040
rect 18509 18037 18521 18040
rect 18555 18068 18567 18071
rect 18782 18068 18788 18080
rect 18555 18040 18788 18068
rect 18555 18037 18567 18040
rect 18509 18031 18567 18037
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 19058 18028 19064 18080
rect 19116 18028 19122 18080
rect 21818 18028 21824 18080
rect 21876 18068 21882 18080
rect 23382 18068 23388 18080
rect 21876 18040 23388 18068
rect 21876 18028 21882 18040
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 26602 18028 26608 18080
rect 26660 18068 26666 18080
rect 30466 18068 30472 18080
rect 26660 18040 30472 18068
rect 26660 18028 26666 18040
rect 30466 18028 30472 18040
rect 30524 18068 30530 18080
rect 30650 18068 30656 18080
rect 30524 18040 30656 18068
rect 30524 18028 30530 18040
rect 30650 18028 30656 18040
rect 30708 18028 30714 18080
rect 32766 18028 32772 18080
rect 32824 18068 32830 18080
rect 33428 18068 33456 18096
rect 32824 18040 33456 18068
rect 37829 18071 37887 18077
rect 32824 18028 32830 18040
rect 37829 18037 37841 18071
rect 37875 18068 37887 18071
rect 37875 18040 38424 18068
rect 37875 18037 37887 18040
rect 37829 18031 37887 18037
rect 38396 18012 38424 18040
rect 1104 17978 38272 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38272 17978
rect 38378 17960 38384 18012
rect 38436 17960 38442 18012
rect 1104 17904 38272 17926
rect 4448 17836 6684 17864
rect 4448 17796 4476 17836
rect 6656 17808 6684 17836
rect 7558 17824 7564 17876
rect 7616 17864 7622 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7616 17836 7665 17864
rect 7616 17824 7622 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 9582 17824 9588 17876
rect 9640 17824 9646 17876
rect 10134 17824 10140 17876
rect 10192 17864 10198 17876
rect 10321 17867 10379 17873
rect 10321 17864 10333 17867
rect 10192 17836 10333 17864
rect 10192 17824 10198 17836
rect 10321 17833 10333 17836
rect 10367 17833 10379 17867
rect 10321 17827 10379 17833
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 11330 17864 11336 17876
rect 10744 17836 11336 17864
rect 10744 17824 10750 17836
rect 11330 17824 11336 17836
rect 11388 17824 11394 17876
rect 11422 17824 11428 17876
rect 11480 17824 11486 17876
rect 11790 17824 11796 17876
rect 11848 17864 11854 17876
rect 12161 17867 12219 17873
rect 12161 17864 12173 17867
rect 11848 17836 12173 17864
rect 11848 17824 11854 17836
rect 12161 17833 12173 17836
rect 12207 17833 12219 17867
rect 15378 17864 15384 17876
rect 12161 17827 12219 17833
rect 14476 17836 15384 17864
rect 4356 17768 4476 17796
rect 3050 17688 3056 17740
rect 3108 17688 3114 17740
rect 4246 17728 4252 17740
rect 4172 17700 4252 17728
rect 3970 17620 3976 17672
rect 4028 17620 4034 17672
rect 4172 17669 4200 17700
rect 4246 17688 4252 17700
rect 4304 17688 4310 17740
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4356 17660 4384 17768
rect 6638 17756 6644 17808
rect 6696 17756 6702 17808
rect 9601 17796 9629 17824
rect 9861 17799 9919 17805
rect 9861 17796 9873 17799
rect 9601 17768 9873 17796
rect 9861 17765 9873 17768
rect 9907 17765 9919 17799
rect 11609 17799 11667 17805
rect 11609 17796 11621 17799
rect 9861 17759 9919 17765
rect 9968 17768 11621 17796
rect 7466 17688 7472 17740
rect 7524 17688 7530 17740
rect 8018 17688 8024 17740
rect 8076 17728 8082 17740
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 8076 17700 8217 17728
rect 8076 17688 8082 17700
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 8662 17688 8668 17740
rect 8720 17688 8726 17740
rect 9217 17731 9275 17737
rect 9217 17697 9229 17731
rect 9263 17728 9275 17731
rect 9674 17728 9680 17740
rect 9263 17700 9680 17728
rect 9263 17697 9275 17700
rect 9217 17691 9275 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 4157 17623 4215 17629
rect 4310 17632 4384 17660
rect 4310 17601 4338 17632
rect 4430 17620 4436 17672
rect 4488 17620 4494 17672
rect 4540 17669 4660 17670
rect 4525 17663 4660 17669
rect 4525 17629 4537 17663
rect 4571 17660 4660 17663
rect 4571 17642 4936 17660
rect 4571 17629 4583 17642
rect 4632 17632 4936 17642
rect 4525 17623 4583 17629
rect 4908 17604 4936 17632
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 5261 17663 5319 17669
rect 5261 17660 5273 17663
rect 5224 17632 5273 17660
rect 5224 17620 5230 17632
rect 5261 17629 5273 17632
rect 5307 17629 5319 17663
rect 5261 17623 5319 17629
rect 4065 17595 4123 17601
rect 4065 17561 4077 17595
rect 4111 17561 4123 17595
rect 4065 17555 4123 17561
rect 4295 17595 4353 17601
rect 4295 17561 4307 17595
rect 4341 17561 4353 17595
rect 4295 17555 4353 17561
rect 4617 17595 4675 17601
rect 4617 17561 4629 17595
rect 4663 17561 4675 17595
rect 4617 17555 4675 17561
rect 2498 17484 2504 17536
rect 2556 17484 2562 17536
rect 2866 17484 2872 17536
rect 2924 17484 2930 17536
rect 2961 17527 3019 17533
rect 2961 17493 2973 17527
rect 3007 17524 3019 17527
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3007 17496 3801 17524
rect 3007 17493 3019 17496
rect 2961 17487 3019 17493
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 4080 17524 4108 17555
rect 4632 17524 4660 17555
rect 4890 17552 4896 17604
rect 4948 17552 4954 17604
rect 5074 17552 5080 17604
rect 5132 17592 5138 17604
rect 5537 17595 5595 17601
rect 5537 17592 5549 17595
rect 5132 17564 5549 17592
rect 5132 17552 5138 17564
rect 5537 17561 5549 17564
rect 5583 17561 5595 17595
rect 5537 17555 5595 17561
rect 5994 17552 6000 17604
rect 6052 17552 6058 17604
rect 7101 17595 7159 17601
rect 7101 17561 7113 17595
rect 7147 17592 7159 17595
rect 7190 17592 7196 17604
rect 7147 17564 7196 17592
rect 7147 17561 7159 17564
rect 7101 17555 7159 17561
rect 7190 17552 7196 17564
rect 7248 17552 7254 17604
rect 7285 17595 7343 17601
rect 7285 17561 7297 17595
rect 7331 17561 7343 17595
rect 8036 17592 8064 17688
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8680 17660 8708 17688
rect 9968 17672 9996 17768
rect 11609 17765 11621 17768
rect 11655 17765 11667 17799
rect 11609 17759 11667 17765
rect 10778 17688 10784 17740
rect 10836 17688 10842 17740
rect 10965 17731 11023 17737
rect 10965 17697 10977 17731
rect 11011 17728 11023 17731
rect 11146 17728 11152 17740
rect 11011 17700 11152 17728
rect 11011 17697 11023 17700
rect 10965 17691 11023 17697
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 11348 17700 14105 17728
rect 8159 17632 8708 17660
rect 9585 17663 9643 17669
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 9585 17629 9597 17663
rect 9631 17629 9643 17663
rect 9585 17623 9643 17629
rect 8662 17592 8668 17604
rect 8036 17564 8668 17592
rect 7285 17555 7343 17561
rect 4080 17496 4660 17524
rect 3789 17487 3847 17493
rect 5442 17484 5448 17536
rect 5500 17524 5506 17536
rect 7009 17527 7067 17533
rect 7009 17524 7021 17527
rect 5500 17496 7021 17524
rect 5500 17484 5506 17496
rect 7009 17493 7021 17496
rect 7055 17524 7067 17527
rect 7300 17524 7328 17555
rect 8662 17552 8668 17564
rect 8720 17552 8726 17604
rect 9600 17592 9628 17623
rect 9950 17620 9956 17672
rect 10008 17620 10014 17672
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 11348 17660 11376 17700
rect 14093 17697 14105 17700
rect 14139 17697 14151 17731
rect 14476 17728 14504 17836
rect 15378 17824 15384 17836
rect 15436 17864 15442 17876
rect 16209 17867 16267 17873
rect 15436 17836 15608 17864
rect 15436 17824 15442 17836
rect 15580 17808 15608 17836
rect 16209 17833 16221 17867
rect 16255 17864 16267 17867
rect 16942 17864 16948 17876
rect 16255 17836 16948 17864
rect 16255 17833 16267 17836
rect 16209 17827 16267 17833
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 18506 17824 18512 17876
rect 18564 17824 18570 17876
rect 20349 17867 20407 17873
rect 20349 17833 20361 17867
rect 20395 17864 20407 17867
rect 20990 17864 20996 17876
rect 20395 17836 20996 17864
rect 20395 17833 20407 17836
rect 20349 17827 20407 17833
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 27154 17824 27160 17876
rect 27212 17864 27218 17876
rect 30374 17864 30380 17876
rect 27212 17836 30380 17864
rect 27212 17824 27218 17836
rect 30374 17824 30380 17836
rect 30432 17824 30438 17876
rect 31202 17824 31208 17876
rect 31260 17864 31266 17876
rect 32306 17864 32312 17876
rect 31260 17836 32312 17864
rect 31260 17824 31266 17836
rect 32306 17824 32312 17836
rect 32364 17824 32370 17876
rect 33321 17867 33379 17873
rect 33321 17864 33333 17867
rect 32692 17836 33333 17864
rect 15286 17796 15292 17808
rect 14093 17691 14151 17697
rect 14384 17700 14504 17728
rect 14568 17768 15292 17796
rect 11287 17632 11376 17660
rect 11425 17663 11483 17669
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11425 17629 11437 17663
rect 11471 17660 11483 17663
rect 11514 17660 11520 17672
rect 11471 17632 11520 17660
rect 11471 17629 11483 17632
rect 11425 17623 11483 17629
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 11698 17620 11704 17672
rect 11756 17660 11762 17672
rect 14384 17669 14412 17700
rect 14568 17672 14596 17768
rect 15286 17756 15292 17768
rect 15344 17756 15350 17808
rect 15562 17756 15568 17808
rect 15620 17796 15626 17808
rect 18524 17796 18552 17824
rect 15620 17768 18552 17796
rect 15620 17756 15626 17768
rect 14752 17700 15240 17728
rect 14369 17663 14427 17669
rect 11756 17632 12020 17660
rect 11756 17620 11762 17632
rect 9766 17592 9772 17604
rect 9600 17564 9772 17592
rect 9766 17552 9772 17564
rect 9824 17552 9830 17604
rect 11992 17601 12020 17632
rect 14369 17629 14381 17663
rect 14415 17629 14427 17663
rect 14369 17623 14427 17629
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17629 14519 17663
rect 14461 17623 14519 17629
rect 10689 17595 10747 17601
rect 10689 17561 10701 17595
rect 10735 17592 10747 17595
rect 11793 17595 11851 17601
rect 11793 17592 11805 17595
rect 10735 17564 11805 17592
rect 10735 17561 10747 17564
rect 10689 17555 10747 17561
rect 11793 17561 11805 17564
rect 11839 17561 11851 17595
rect 11793 17555 11851 17561
rect 11977 17595 12035 17601
rect 11977 17561 11989 17595
rect 12023 17592 12035 17595
rect 13078 17592 13084 17604
rect 12023 17564 13084 17592
rect 12023 17561 12035 17564
rect 11977 17555 12035 17561
rect 7055 17496 7328 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 8018 17484 8024 17536
rect 8076 17484 8082 17536
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 10410 17524 10416 17536
rect 9640 17496 10416 17524
rect 9640 17484 9646 17496
rect 10410 17484 10416 17496
rect 10468 17484 10474 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11698 17524 11704 17536
rect 11020 17496 11704 17524
rect 11020 17484 11026 17496
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 11808 17524 11836 17555
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 13262 17552 13268 17604
rect 13320 17592 13326 17604
rect 14476 17592 14504 17623
rect 14550 17620 14556 17672
rect 14608 17620 14614 17672
rect 14752 17669 14780 17700
rect 15212 17672 15240 17700
rect 15488 17700 16620 17728
rect 14737 17663 14795 17669
rect 14737 17629 14749 17663
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 14936 17592 14964 17623
rect 15010 17620 15016 17672
rect 15068 17620 15074 17672
rect 15194 17620 15200 17672
rect 15252 17620 15258 17672
rect 15488 17592 15516 17700
rect 15565 17663 15623 17669
rect 15565 17629 15577 17663
rect 15611 17660 15623 17663
rect 15654 17660 15660 17672
rect 15611 17632 15660 17660
rect 15611 17629 15623 17632
rect 15565 17623 15623 17629
rect 13320 17564 15516 17592
rect 13320 17552 13326 17564
rect 12158 17524 12164 17536
rect 11808 17496 12164 17524
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14182 17524 14188 17536
rect 14056 17496 14188 17524
rect 14056 17484 14062 17496
rect 14182 17484 14188 17496
rect 14240 17524 14246 17536
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 14240 17496 14933 17524
rect 14240 17484 14246 17496
rect 14921 17493 14933 17496
rect 14967 17493 14979 17527
rect 14921 17487 14979 17493
rect 15378 17484 15384 17536
rect 15436 17484 15442 17536
rect 15580 17524 15608 17623
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 15746 17620 15752 17672
rect 15804 17620 15810 17672
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15856 17592 15884 17623
rect 16390 17620 16396 17672
rect 16448 17620 16454 17672
rect 16482 17620 16488 17672
rect 16540 17620 16546 17672
rect 16592 17660 16620 17700
rect 16666 17688 16672 17740
rect 16724 17688 16730 17740
rect 16776 17737 16804 17768
rect 18690 17756 18696 17808
rect 18748 17796 18754 17808
rect 20714 17796 20720 17808
rect 18748 17768 20720 17796
rect 18748 17756 18754 17768
rect 20714 17756 20720 17768
rect 20772 17756 20778 17808
rect 23290 17756 23296 17808
rect 23348 17796 23354 17808
rect 23348 17768 24716 17796
rect 23348 17756 23354 17768
rect 16761 17731 16819 17737
rect 16761 17697 16773 17731
rect 16807 17697 16819 17731
rect 16761 17691 16819 17697
rect 16868 17700 18460 17728
rect 16868 17660 16896 17700
rect 18432 17672 18460 17700
rect 18506 17688 18512 17740
rect 18564 17728 18570 17740
rect 19794 17728 19800 17740
rect 18564 17700 19800 17728
rect 18564 17688 18570 17700
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 19886 17688 19892 17740
rect 19944 17728 19950 17740
rect 20254 17728 20260 17740
rect 19944 17700 20260 17728
rect 19944 17688 19950 17700
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 20732 17700 21312 17728
rect 16592 17632 16896 17660
rect 18138 17620 18144 17672
rect 18196 17620 18202 17672
rect 18414 17620 18420 17672
rect 18472 17620 18478 17672
rect 19334 17620 19340 17672
rect 19392 17620 19398 17672
rect 20070 17660 20076 17672
rect 19465 17632 20076 17660
rect 16500 17592 16528 17620
rect 15856 17564 16528 17592
rect 16574 17552 16580 17604
rect 16632 17592 16638 17604
rect 16942 17592 16948 17604
rect 16632 17564 16948 17592
rect 16632 17552 16638 17564
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 19465 17592 19493 17632
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20530 17620 20536 17672
rect 20588 17660 20594 17672
rect 20732 17669 20760 17700
rect 20625 17663 20683 17669
rect 20625 17660 20637 17663
rect 20588 17632 20637 17660
rect 20588 17620 20594 17632
rect 20625 17629 20637 17632
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17660 20867 17663
rect 20898 17660 20904 17672
rect 20855 17632 20904 17660
rect 20855 17629 20867 17632
rect 20809 17623 20867 17629
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17629 21051 17663
rect 20993 17623 21051 17629
rect 18248 17564 19493 17592
rect 19521 17595 19579 17601
rect 15930 17524 15936 17536
rect 15580 17496 15936 17524
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 18248 17533 18276 17564
rect 19521 17561 19533 17595
rect 19567 17592 19579 17595
rect 19567 17564 20208 17592
rect 19567 17561 19579 17564
rect 19521 17555 19579 17561
rect 18233 17527 18291 17533
rect 18233 17524 18245 17527
rect 16080 17496 18245 17524
rect 16080 17484 16086 17496
rect 18233 17493 18245 17496
rect 18279 17493 18291 17527
rect 18233 17487 18291 17493
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 19536 17524 19564 17555
rect 18472 17496 19564 17524
rect 18472 17484 18478 17496
rect 19610 17484 19616 17536
rect 19668 17524 19674 17536
rect 19705 17527 19763 17533
rect 19705 17524 19717 17527
rect 19668 17496 19717 17524
rect 19668 17484 19674 17496
rect 19705 17493 19717 17496
rect 19751 17493 19763 17527
rect 20180 17524 20208 17564
rect 20254 17552 20260 17604
rect 20312 17592 20318 17604
rect 21008 17592 21036 17623
rect 21284 17604 21312 17700
rect 23842 17688 23848 17740
rect 23900 17688 23906 17740
rect 24121 17731 24179 17737
rect 24121 17697 24133 17731
rect 24167 17728 24179 17731
rect 24489 17731 24547 17737
rect 24489 17728 24501 17731
rect 24167 17700 24501 17728
rect 24167 17697 24179 17700
rect 24121 17691 24179 17697
rect 24489 17697 24501 17700
rect 24535 17697 24547 17731
rect 24489 17691 24547 17697
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 24210 17660 24216 17672
rect 23799 17632 24216 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 24210 17620 24216 17632
rect 24268 17620 24274 17672
rect 24578 17620 24584 17672
rect 24636 17620 24642 17672
rect 24688 17660 24716 17768
rect 24946 17756 24952 17808
rect 25004 17756 25010 17808
rect 25777 17799 25835 17805
rect 25777 17765 25789 17799
rect 25823 17765 25835 17799
rect 25777 17759 25835 17765
rect 26421 17799 26479 17805
rect 26421 17765 26433 17799
rect 26467 17796 26479 17799
rect 28902 17796 28908 17808
rect 26467 17768 26648 17796
rect 26467 17765 26479 17768
rect 26421 17759 26479 17765
rect 25130 17688 25136 17740
rect 25188 17728 25194 17740
rect 25317 17731 25375 17737
rect 25317 17728 25329 17731
rect 25188 17700 25329 17728
rect 25188 17688 25194 17700
rect 25317 17697 25329 17700
rect 25363 17697 25375 17731
rect 25792 17728 25820 17759
rect 26620 17737 26648 17768
rect 27448 17768 28908 17796
rect 25961 17731 26019 17737
rect 25961 17728 25973 17731
rect 25792 17700 25973 17728
rect 25317 17691 25375 17697
rect 25961 17697 25973 17700
rect 26007 17697 26019 17731
rect 25961 17691 26019 17697
rect 26605 17731 26663 17737
rect 26605 17697 26617 17731
rect 26651 17697 26663 17731
rect 27448 17728 27476 17768
rect 28902 17756 28908 17768
rect 28960 17756 28966 17808
rect 29917 17799 29975 17805
rect 29917 17765 29929 17799
rect 29963 17796 29975 17799
rect 30006 17796 30012 17808
rect 29963 17768 30012 17796
rect 29963 17765 29975 17768
rect 29917 17759 29975 17765
rect 30006 17756 30012 17768
rect 30064 17756 30070 17808
rect 32214 17756 32220 17808
rect 32272 17756 32278 17808
rect 26605 17691 26663 17697
rect 26804 17700 27476 17728
rect 25409 17663 25467 17669
rect 25409 17660 25421 17663
rect 24688 17632 25421 17660
rect 25409 17629 25421 17632
rect 25455 17660 25467 17663
rect 25590 17660 25596 17672
rect 25455 17632 25596 17660
rect 25455 17629 25467 17632
rect 25409 17623 25467 17629
rect 25590 17620 25596 17632
rect 25648 17620 25654 17672
rect 26053 17663 26111 17669
rect 26053 17629 26065 17663
rect 26099 17629 26111 17663
rect 26053 17623 26111 17629
rect 26697 17663 26755 17669
rect 26697 17629 26709 17663
rect 26743 17629 26755 17663
rect 26697 17623 26755 17629
rect 20312 17564 21036 17592
rect 20312 17552 20318 17564
rect 21266 17552 21272 17604
rect 21324 17552 21330 17604
rect 23201 17595 23259 17601
rect 23201 17561 23213 17595
rect 23247 17592 23259 17595
rect 24762 17592 24768 17604
rect 23247 17564 24768 17592
rect 23247 17561 23259 17564
rect 23201 17555 23259 17561
rect 24762 17552 24768 17564
rect 24820 17552 24826 17604
rect 24946 17552 24952 17604
rect 25004 17592 25010 17604
rect 26068 17592 26096 17623
rect 25004 17564 26096 17592
rect 25004 17552 25010 17564
rect 26602 17552 26608 17604
rect 26660 17592 26666 17604
rect 26712 17592 26740 17623
rect 26660 17564 26740 17592
rect 26660 17552 26666 17564
rect 23934 17524 23940 17536
rect 20180 17496 23940 17524
rect 19705 17487 19763 17493
rect 23934 17484 23940 17496
rect 23992 17524 23998 17536
rect 26804 17524 26832 17700
rect 27448 17669 27476 17700
rect 27614 17688 27620 17740
rect 27672 17728 27678 17740
rect 28353 17731 28411 17737
rect 28353 17728 28365 17731
rect 27672 17700 28365 17728
rect 27672 17688 27678 17700
rect 28353 17697 28365 17700
rect 28399 17697 28411 17731
rect 29454 17728 29460 17740
rect 28353 17691 28411 17697
rect 28644 17700 29460 17728
rect 27249 17663 27307 17669
rect 27249 17660 27261 17663
rect 27080 17632 27261 17660
rect 27080 17533 27108 17632
rect 27249 17629 27261 17632
rect 27295 17629 27307 17663
rect 27249 17623 27307 17629
rect 27433 17663 27491 17669
rect 27433 17629 27445 17663
rect 27479 17660 27491 17663
rect 27525 17663 27583 17669
rect 27525 17660 27537 17663
rect 27479 17632 27537 17660
rect 27479 17629 27491 17632
rect 27433 17623 27491 17629
rect 27525 17629 27537 17632
rect 27571 17629 27583 17663
rect 27525 17623 27583 17629
rect 27982 17620 27988 17672
rect 28040 17620 28046 17672
rect 28644 17669 28672 17700
rect 29454 17688 29460 17700
rect 29512 17688 29518 17740
rect 30116 17700 30420 17728
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17629 28687 17663
rect 28629 17623 28687 17629
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17629 28871 17663
rect 28813 17623 28871 17629
rect 27341 17595 27399 17601
rect 27341 17561 27353 17595
rect 27387 17592 27399 17595
rect 28828 17592 28856 17623
rect 29822 17620 29828 17672
rect 29880 17620 29886 17672
rect 29914 17620 29920 17672
rect 29972 17660 29978 17672
rect 30009 17663 30067 17669
rect 30009 17660 30021 17663
rect 29972 17632 30021 17660
rect 29972 17620 29978 17632
rect 30009 17629 30021 17632
rect 30055 17629 30067 17663
rect 30009 17623 30067 17629
rect 27387 17564 28856 17592
rect 29840 17592 29868 17620
rect 30116 17592 30144 17700
rect 30285 17663 30343 17669
rect 30285 17660 30297 17663
rect 30208 17632 30297 17660
rect 30208 17604 30236 17632
rect 30285 17629 30297 17632
rect 30331 17629 30343 17663
rect 30285 17623 30343 17629
rect 29840 17564 30144 17592
rect 27387 17561 27399 17564
rect 27341 17555 27399 17561
rect 30190 17552 30196 17604
rect 30248 17552 30254 17604
rect 30392 17592 30420 17700
rect 31386 17688 31392 17740
rect 31444 17688 31450 17740
rect 31754 17688 31760 17740
rect 31812 17728 31818 17740
rect 32232 17728 32260 17756
rect 32692 17728 32720 17836
rect 33321 17833 33333 17836
rect 33367 17833 33379 17867
rect 33321 17827 33379 17833
rect 33689 17867 33747 17873
rect 33689 17833 33701 17867
rect 33735 17864 33747 17867
rect 33778 17864 33784 17876
rect 33735 17836 33784 17864
rect 33735 17833 33747 17836
rect 33689 17827 33747 17833
rect 32769 17799 32827 17805
rect 32769 17765 32781 17799
rect 32815 17796 32827 17799
rect 33704 17796 33732 17827
rect 33778 17824 33784 17836
rect 33836 17824 33842 17876
rect 32815 17768 33732 17796
rect 33980 17768 34468 17796
rect 32815 17765 32827 17768
rect 32769 17759 32827 17765
rect 31812 17700 31857 17728
rect 32232 17700 33088 17728
rect 31812 17688 31818 17700
rect 30466 17620 30472 17672
rect 30524 17620 30530 17672
rect 31570 17620 31576 17672
rect 31628 17620 31634 17672
rect 31662 17620 31668 17672
rect 31720 17620 31726 17672
rect 31846 17620 31852 17672
rect 31904 17660 31910 17672
rect 32490 17660 32496 17672
rect 31904 17632 32496 17660
rect 31904 17620 31910 17632
rect 32490 17620 32496 17632
rect 32548 17660 32554 17672
rect 32858 17660 32864 17672
rect 32548 17632 32864 17660
rect 32548 17620 32554 17632
rect 32858 17620 32864 17632
rect 32916 17620 32922 17672
rect 33060 17669 33088 17700
rect 33134 17688 33140 17740
rect 33192 17728 33198 17740
rect 33781 17731 33839 17737
rect 33781 17728 33793 17731
rect 33192 17700 33793 17728
rect 33192 17688 33198 17700
rect 33781 17697 33793 17700
rect 33827 17728 33839 17731
rect 33980 17728 34008 17768
rect 34440 17737 34468 17768
rect 34241 17731 34299 17737
rect 34241 17728 34253 17731
rect 33827 17700 34008 17728
rect 34072 17700 34253 17728
rect 33827 17697 33839 17700
rect 33781 17691 33839 17697
rect 33045 17663 33103 17669
rect 33045 17629 33057 17663
rect 33091 17629 33103 17663
rect 33410 17660 33416 17672
rect 33368 17635 33416 17660
rect 33045 17623 33103 17629
rect 33367 17629 33416 17635
rect 30392 17564 32720 17592
rect 32692 17536 32720 17564
rect 32766 17552 32772 17604
rect 32824 17552 32830 17604
rect 33134 17592 33140 17604
rect 33060 17564 33140 17592
rect 23992 17496 26832 17524
rect 27065 17527 27123 17533
rect 23992 17484 23998 17496
rect 27065 17493 27077 17527
rect 27111 17493 27123 17527
rect 27065 17487 27123 17493
rect 28718 17484 28724 17536
rect 28776 17524 28782 17536
rect 30377 17527 30435 17533
rect 30377 17524 30389 17527
rect 28776 17496 30389 17524
rect 28776 17484 28782 17496
rect 30377 17493 30389 17496
rect 30423 17524 30435 17527
rect 31662 17524 31668 17536
rect 30423 17496 31668 17524
rect 30423 17493 30435 17496
rect 30377 17487 30435 17493
rect 31662 17484 31668 17496
rect 31720 17484 31726 17536
rect 32674 17484 32680 17536
rect 32732 17524 32738 17536
rect 32953 17527 33011 17533
rect 32953 17524 32965 17527
rect 32732 17496 32965 17524
rect 32732 17484 32738 17496
rect 32953 17493 32965 17496
rect 32999 17524 33011 17527
rect 33060 17524 33088 17564
rect 33134 17552 33140 17564
rect 33192 17552 33198 17604
rect 33367 17595 33379 17629
rect 33413 17620 33416 17629
rect 33468 17620 33474 17672
rect 33689 17663 33747 17669
rect 33689 17629 33701 17663
rect 33735 17660 33747 17663
rect 34072 17660 34100 17700
rect 34241 17697 34253 17700
rect 34287 17697 34299 17731
rect 34241 17691 34299 17697
rect 34425 17731 34483 17737
rect 34425 17697 34437 17731
rect 34471 17697 34483 17731
rect 34425 17691 34483 17697
rect 33735 17632 34100 17660
rect 34149 17663 34207 17669
rect 33735 17629 33747 17632
rect 33689 17623 33747 17629
rect 34149 17629 34161 17663
rect 34195 17629 34207 17663
rect 34149 17623 34207 17629
rect 33413 17595 33425 17620
rect 33367 17589 33425 17595
rect 32999 17496 33088 17524
rect 33505 17527 33563 17533
rect 32999 17493 33011 17496
rect 32953 17487 33011 17493
rect 33505 17493 33517 17527
rect 33551 17524 33563 17527
rect 33704 17524 33732 17623
rect 33778 17552 33784 17604
rect 33836 17592 33842 17604
rect 34164 17592 34192 17623
rect 33836 17564 34192 17592
rect 33836 17552 33842 17564
rect 33551 17496 33732 17524
rect 33551 17493 33563 17496
rect 33505 17487 33563 17493
rect 34054 17484 34060 17536
rect 34112 17484 34118 17536
rect 34422 17484 34428 17536
rect 34480 17484 34486 17536
rect 1104 17434 38272 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38272 17434
rect 1104 17360 38272 17382
rect 5166 17320 5172 17332
rect 1412 17292 5172 17320
rect 1412 17196 1440 17292
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 5353 17323 5411 17329
rect 5353 17289 5365 17323
rect 5399 17289 5411 17323
rect 5353 17283 5411 17289
rect 3970 17212 3976 17264
rect 4028 17212 4034 17264
rect 4525 17255 4583 17261
rect 4525 17221 4537 17255
rect 4571 17221 4583 17255
rect 4525 17215 4583 17221
rect 1394 17144 1400 17196
rect 1452 17144 1458 17196
rect 2774 17144 2780 17196
rect 2832 17144 2838 17196
rect 1670 17076 1676 17128
rect 1728 17076 1734 17128
rect 3881 17119 3939 17125
rect 3881 17085 3893 17119
rect 3927 17116 3939 17119
rect 3988 17116 4016 17212
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4540 17184 4568 17215
rect 4706 17212 4712 17264
rect 4764 17261 4770 17264
rect 4764 17255 4783 17261
rect 4771 17221 4783 17255
rect 4764 17215 4783 17221
rect 4764 17212 4770 17215
rect 4203 17156 4568 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 3927 17088 4016 17116
rect 3927 17085 3939 17088
rect 3881 17079 3939 17085
rect 4062 17076 4068 17128
rect 4120 17076 4126 17128
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17085 4399 17119
rect 4540 17116 4568 17156
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17184 5319 17187
rect 5368 17184 5396 17283
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 5500 17292 5733 17320
rect 5500 17280 5506 17292
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 5721 17283 5779 17289
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 10965 17323 11023 17329
rect 10965 17320 10977 17323
rect 10836 17292 10977 17320
rect 10836 17280 10842 17292
rect 10965 17289 10977 17292
rect 11011 17289 11023 17323
rect 10965 17283 11023 17289
rect 11054 17280 11060 17332
rect 11112 17280 11118 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11241 17323 11299 17329
rect 11241 17320 11253 17323
rect 11204 17292 11253 17320
rect 11204 17280 11210 17292
rect 11241 17289 11253 17292
rect 11287 17289 11299 17323
rect 11241 17283 11299 17289
rect 11422 17280 11428 17332
rect 11480 17320 11486 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11480 17292 11621 17320
rect 11480 17280 11486 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 12158 17280 12164 17332
rect 12216 17280 12222 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 13354 17320 13360 17332
rect 13219 17292 13360 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 14366 17280 14372 17332
rect 14424 17280 14430 17332
rect 16114 17280 16120 17332
rect 16172 17320 16178 17332
rect 16209 17323 16267 17329
rect 16209 17320 16221 17323
rect 16172 17292 16221 17320
rect 16172 17280 16178 17292
rect 16209 17289 16221 17292
rect 16255 17320 16267 17323
rect 16482 17320 16488 17332
rect 16255 17292 16488 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 16666 17280 16672 17332
rect 16724 17320 16730 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 16724 17292 17417 17320
rect 16724 17280 16730 17292
rect 17405 17289 17417 17292
rect 17451 17289 17463 17323
rect 17405 17283 17463 17289
rect 5307 17156 5396 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 4798 17116 4804 17128
rect 4540 17088 4804 17116
rect 4341 17079 4399 17085
rect 3970 17008 3976 17060
rect 4028 17048 4034 17060
rect 4154 17048 4160 17060
rect 4028 17020 4160 17048
rect 4028 17008 4034 17020
rect 4154 17008 4160 17020
rect 4212 17048 4218 17060
rect 4264 17048 4292 17079
rect 4212 17020 4292 17048
rect 4356 17048 4384 17079
rect 4798 17076 4804 17088
rect 4856 17116 4862 17128
rect 5460 17116 5488 17280
rect 9766 17252 9772 17264
rect 9508 17224 9772 17252
rect 9214 17144 9220 17196
rect 9272 17144 9278 17196
rect 9508 17193 9536 17224
rect 9766 17212 9772 17224
rect 9824 17252 9830 17264
rect 11072 17252 11100 17280
rect 11440 17252 11468 17280
rect 12176 17252 12204 17280
rect 9824 17224 11100 17252
rect 11164 17224 11468 17252
rect 11624 17224 12204 17252
rect 9824 17212 9830 17224
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 9586 17187 9644 17193
rect 9586 17153 9598 17187
rect 9632 17184 9644 17187
rect 9674 17184 9680 17196
rect 9632 17156 9680 17184
rect 9632 17153 9644 17156
rect 9586 17147 9644 17153
rect 4856 17088 5488 17116
rect 4856 17076 4862 17088
rect 5810 17076 5816 17128
rect 5868 17076 5874 17128
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17116 6055 17119
rect 6086 17116 6092 17128
rect 6043 17088 6092 17116
rect 6043 17085 6055 17088
rect 5997 17079 6055 17085
rect 4356 17020 4752 17048
rect 4212 17008 4218 17020
rect 2866 16940 2872 16992
rect 2924 16980 2930 16992
rect 3145 16983 3203 16989
rect 3145 16980 3157 16983
rect 2924 16952 3157 16980
rect 2924 16940 2930 16952
rect 3145 16949 3157 16952
rect 3191 16980 3203 16983
rect 4356 16980 4384 17020
rect 4724 16989 4752 17020
rect 4890 17008 4896 17060
rect 4948 17008 4954 17060
rect 5000 17020 5488 17048
rect 3191 16952 4384 16980
rect 4709 16983 4767 16989
rect 3191 16949 3203 16952
rect 3145 16943 3203 16949
rect 4709 16949 4721 16983
rect 4755 16980 4767 16983
rect 5000 16980 5028 17020
rect 5460 16992 5488 17020
rect 4755 16952 5028 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 5074 16940 5080 16992
rect 5132 16940 5138 16992
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 6012 16980 6040 17079
rect 6086 17076 6092 17088
rect 6144 17076 6150 17128
rect 9416 17116 9444 17147
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 10888 17116 10916 17147
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 11164 17193 11192 17224
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 11020 17156 11069 17184
rect 11020 17144 11026 17156
rect 11057 17153 11069 17156
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17153 11207 17187
rect 11149 17147 11207 17153
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11296 17156 11345 17184
rect 11296 17144 11302 17156
rect 11333 17153 11345 17156
rect 11379 17153 11391 17187
rect 11333 17147 11391 17153
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11480 17156 11529 17184
rect 11480 17144 11486 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 11624 17116 11652 17224
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 12897 17255 12955 17261
rect 12897 17252 12909 17255
rect 12400 17224 12909 17252
rect 12400 17212 12406 17224
rect 12897 17221 12909 17224
rect 12943 17221 12955 17255
rect 12897 17215 12955 17221
rect 13446 17212 13452 17264
rect 13504 17212 13510 17264
rect 14384 17252 14412 17280
rect 15286 17252 15292 17264
rect 14384 17224 15292 17252
rect 15286 17212 15292 17224
rect 15344 17252 15350 17264
rect 15344 17224 15608 17252
rect 15344 17212 15350 17224
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 11793 17187 11851 17193
rect 11793 17153 11805 17187
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 9416 17088 10824 17116
rect 10888 17088 11652 17116
rect 11808 17116 11836 17147
rect 11974 17144 11980 17196
rect 12032 17144 12038 17196
rect 12069 17187 12127 17193
rect 12069 17153 12081 17187
rect 12115 17184 12127 17187
rect 12158 17184 12164 17196
rect 12115 17156 12164 17184
rect 12115 17153 12127 17156
rect 12069 17147 12127 17153
rect 12084 17116 12112 17147
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12434 17184 12440 17196
rect 12299 17156 12440 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 11808 17088 12112 17116
rect 6638 17008 6644 17060
rect 6696 17048 6702 17060
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 6696 17020 9873 17048
rect 6696 17008 6702 17020
rect 9861 17017 9873 17020
rect 9907 17017 9919 17051
rect 9861 17011 9919 17017
rect 9950 17008 9956 17060
rect 10008 17008 10014 17060
rect 10796 17048 10824 17088
rect 12268 17060 12296 17147
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 13078 17144 13084 17196
rect 13136 17144 13142 17196
rect 13305 17187 13363 17193
rect 13305 17153 13317 17187
rect 13351 17184 13363 17187
rect 14921 17187 14979 17193
rect 13351 17156 14872 17184
rect 13351 17153 13363 17156
rect 13305 17147 13363 17153
rect 10796 17020 12020 17048
rect 5592 16952 6040 16980
rect 5592 16940 5598 16952
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 9968 16980 9996 17008
rect 9272 16952 9996 16980
rect 9272 16940 9278 16952
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 11480 16952 11897 16980
rect 11480 16940 11486 16952
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 11992 16980 12020 17020
rect 12250 17008 12256 17060
rect 12308 17008 12314 17060
rect 14182 16980 14188 16992
rect 11992 16952 14188 16980
rect 11885 16943 11943 16949
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 14737 16983 14795 16989
rect 14737 16980 14749 16983
rect 14424 16952 14749 16980
rect 14424 16940 14430 16952
rect 14737 16949 14749 16952
rect 14783 16949 14795 16983
rect 14844 16980 14872 17156
rect 14921 17153 14933 17187
rect 14967 17184 14979 17187
rect 15378 17184 15384 17196
rect 14967 17156 15384 17184
rect 14967 17153 14979 17156
rect 14921 17147 14979 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 15580 17193 15608 17224
rect 15838 17212 15844 17264
rect 15896 17252 15902 17264
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15896 17224 15945 17252
rect 15896 17212 15902 17224
rect 15933 17221 15945 17224
rect 15979 17252 15991 17255
rect 16390 17252 16396 17264
rect 15979 17224 16396 17252
rect 15979 17221 15991 17224
rect 15933 17215 15991 17221
rect 15746 17193 15752 17196
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 15719 17187 15752 17193
rect 15719 17153 15731 17187
rect 15719 17147 15752 17153
rect 15746 17144 15752 17147
rect 15804 17144 15810 17196
rect 16022 17144 16028 17196
rect 16080 17144 16086 17196
rect 16316 17193 16344 17224
rect 16390 17212 16396 17224
rect 16448 17252 16454 17264
rect 17420 17252 17448 17283
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 18690 17320 18696 17332
rect 17552 17292 18696 17320
rect 17552 17280 17558 17292
rect 16448 17224 17356 17252
rect 17420 17224 17724 17252
rect 16448 17212 16454 17224
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16540 17156 16865 17184
rect 16540 17144 16546 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17000 17156 17233 17184
rect 17000 17144 17006 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17328 17184 17356 17224
rect 17696 17193 17724 17224
rect 18230 17212 18236 17264
rect 18288 17252 18294 17264
rect 18414 17252 18420 17264
rect 18288 17224 18420 17252
rect 18288 17212 18294 17224
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 17497 17187 17555 17193
rect 17497 17184 17509 17187
rect 17328 17156 17509 17184
rect 17221 17147 17279 17153
rect 17497 17153 17509 17156
rect 17543 17153 17555 17187
rect 17497 17147 17555 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 18322 17184 18328 17196
rect 17681 17147 17739 17153
rect 17880 17156 18328 17184
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 15252 17088 16436 17116
rect 15252 17076 15258 17088
rect 15105 17051 15163 17057
rect 15105 17017 15117 17051
rect 15151 17048 15163 17051
rect 16025 17051 16083 17057
rect 16025 17048 16037 17051
rect 15151 17020 16037 17048
rect 15151 17017 15163 17020
rect 15105 17011 15163 17017
rect 16025 17017 16037 17020
rect 16071 17017 16083 17051
rect 16025 17011 16083 17017
rect 16298 16980 16304 16992
rect 14844 16952 16304 16980
rect 14737 16943 14795 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 16408 16980 16436 17088
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 16761 17119 16819 17125
rect 16761 17116 16773 17119
rect 16724 17088 16773 17116
rect 16724 17076 16730 17088
rect 16761 17085 16773 17088
rect 16807 17116 16819 17119
rect 17880 17116 17908 17156
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 18616 17193 18644 17292
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 18874 17280 18880 17332
rect 18932 17280 18938 17332
rect 19886 17280 19892 17332
rect 19944 17280 19950 17332
rect 20254 17280 20260 17332
rect 20312 17280 20318 17332
rect 20622 17320 20628 17332
rect 20371 17292 20628 17320
rect 19904 17252 19932 17280
rect 19981 17255 20039 17261
rect 19981 17252 19993 17255
rect 19306 17224 19748 17252
rect 19904 17224 19993 17252
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 16807 17088 17908 17116
rect 16807 17085 16819 17088
rect 16761 17079 16819 17085
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18230 17116 18236 17128
rect 18012 17088 18236 17116
rect 18012 17076 18018 17088
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 18340 17048 18368 17144
rect 18693 17119 18751 17125
rect 18693 17085 18705 17119
rect 18739 17116 18751 17119
rect 18874 17116 18880 17128
rect 18739 17088 18880 17116
rect 18739 17085 18751 17088
rect 18693 17079 18751 17085
rect 18874 17076 18880 17088
rect 18932 17076 18938 17128
rect 19306 17048 19334 17224
rect 19720 17193 19748 17224
rect 19981 17221 19993 17224
rect 20027 17221 20039 17255
rect 19981 17215 20039 17221
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 19706 17187 19764 17193
rect 19706 17153 19718 17187
rect 19752 17153 19764 17187
rect 19706 17147 19764 17153
rect 19628 17116 19656 17147
rect 19886 17144 19892 17196
rect 19944 17144 19950 17196
rect 20070 17144 20076 17196
rect 20128 17193 20134 17196
rect 20371 17193 20399 17292
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17289 21051 17323
rect 20993 17283 21051 17289
rect 20714 17212 20720 17264
rect 20772 17212 20778 17264
rect 21008 17252 21036 17283
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 24213 17323 24271 17329
rect 21416 17292 23520 17320
rect 21416 17280 21422 17292
rect 21008 17224 22692 17252
rect 20128 17184 20136 17193
rect 20349 17187 20407 17193
rect 20128 17156 20173 17184
rect 20128 17147 20136 17156
rect 20349 17153 20361 17187
rect 20395 17153 20407 17187
rect 20349 17147 20407 17153
rect 20497 17187 20555 17193
rect 20497 17153 20509 17187
rect 20543 17184 20555 17187
rect 20543 17153 20576 17184
rect 20497 17147 20576 17153
rect 20128 17144 20134 17147
rect 19628 17088 20300 17116
rect 17052 17020 17632 17048
rect 18340 17020 19334 17048
rect 17052 16980 17080 17020
rect 16408 16952 17080 16980
rect 17126 16940 17132 16992
rect 17184 16940 17190 16992
rect 17494 16940 17500 16992
rect 17552 16940 17558 16992
rect 17604 16980 17632 17020
rect 19886 17008 19892 17060
rect 19944 17008 19950 17060
rect 19904 16980 19932 17008
rect 17604 16952 19932 16980
rect 20272 16980 20300 17088
rect 20371 17060 20399 17147
rect 20548 17116 20576 17147
rect 20622 17144 20628 17196
rect 20680 17144 20686 17196
rect 20898 17193 20904 17196
rect 20855 17187 20904 17193
rect 20855 17153 20867 17187
rect 20901 17153 20904 17187
rect 20855 17147 20904 17153
rect 20898 17144 20904 17147
rect 20956 17144 20962 17196
rect 20990 17144 20996 17196
rect 21048 17144 21054 17196
rect 21174 17144 21180 17196
rect 21232 17144 21238 17196
rect 21284 17193 21312 17224
rect 22664 17193 22692 17224
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17153 21327 17187
rect 22189 17187 22247 17193
rect 22189 17184 22201 17187
rect 21269 17147 21327 17153
rect 21376 17156 22201 17184
rect 21008 17116 21036 17144
rect 20548 17088 21036 17116
rect 21082 17076 21088 17128
rect 21140 17076 21146 17128
rect 21192 17116 21220 17144
rect 21376 17116 21404 17156
rect 22189 17153 22201 17156
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 22649 17187 22707 17193
rect 22649 17153 22661 17187
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 23201 17187 23259 17193
rect 23201 17153 23213 17187
rect 23247 17184 23259 17187
rect 23382 17184 23388 17196
rect 23247 17156 23388 17184
rect 23247 17153 23259 17156
rect 23201 17147 23259 17153
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 23492 17184 23520 17292
rect 24213 17289 24225 17323
rect 24259 17320 24271 17323
rect 24578 17320 24584 17332
rect 24259 17292 24584 17320
rect 24259 17289 24271 17292
rect 24213 17283 24271 17289
rect 24578 17280 24584 17292
rect 24636 17280 24642 17332
rect 25590 17280 25596 17332
rect 25648 17320 25654 17332
rect 28074 17320 28080 17332
rect 25648 17292 28080 17320
rect 25648 17280 25654 17292
rect 28074 17280 28080 17292
rect 28132 17280 28138 17332
rect 28350 17280 28356 17332
rect 28408 17280 28414 17332
rect 29012 17292 29224 17320
rect 29012 17252 29040 17292
rect 29196 17264 29224 17292
rect 29454 17280 29460 17332
rect 29512 17280 29518 17332
rect 31386 17280 31392 17332
rect 31444 17280 31450 17332
rect 31570 17280 31576 17332
rect 31628 17280 31634 17332
rect 31662 17280 31668 17332
rect 31720 17320 31726 17332
rect 31849 17323 31907 17329
rect 31849 17320 31861 17323
rect 31720 17292 31861 17320
rect 31720 17280 31726 17292
rect 31849 17289 31861 17292
rect 31895 17289 31907 17323
rect 31849 17283 31907 17289
rect 34054 17280 34060 17332
rect 34112 17320 34118 17332
rect 34149 17323 34207 17329
rect 34149 17320 34161 17323
rect 34112 17292 34161 17320
rect 34112 17280 34118 17292
rect 34149 17289 34161 17292
rect 34195 17289 34207 17323
rect 34149 17283 34207 17289
rect 28276 17224 29040 17252
rect 23845 17187 23903 17193
rect 23845 17184 23857 17187
rect 23492 17156 23857 17184
rect 23845 17153 23857 17156
rect 23891 17184 23903 17187
rect 24302 17184 24308 17196
rect 23891 17156 24308 17184
rect 23891 17153 23903 17156
rect 23845 17147 23903 17153
rect 24302 17144 24308 17156
rect 24360 17144 24366 17196
rect 28276 17193 28304 17224
rect 29086 17212 29092 17264
rect 29144 17212 29150 17264
rect 29178 17212 29184 17264
rect 29236 17252 29242 17264
rect 29289 17255 29347 17261
rect 29289 17252 29301 17255
rect 29236 17224 29301 17252
rect 29236 17212 29242 17224
rect 29289 17221 29301 17224
rect 29335 17221 29347 17255
rect 29289 17215 29347 17221
rect 30466 17212 30472 17264
rect 30524 17252 30530 17264
rect 31404 17252 31432 17280
rect 34164 17252 34192 17283
rect 34422 17280 34428 17332
rect 34480 17280 34486 17332
rect 34701 17323 34759 17329
rect 34701 17289 34713 17323
rect 34747 17320 34759 17323
rect 34747 17292 34836 17320
rect 34747 17289 34759 17292
rect 34701 17283 34759 17289
rect 34333 17255 34391 17261
rect 34333 17252 34345 17255
rect 30524 17224 31340 17252
rect 31404 17224 32352 17252
rect 34164 17224 34345 17252
rect 30524 17212 30530 17224
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28169 17187 28227 17193
rect 28169 17153 28181 17187
rect 28215 17153 28227 17187
rect 28169 17147 28227 17153
rect 28261 17187 28319 17193
rect 28261 17153 28273 17187
rect 28307 17153 28319 17187
rect 28261 17147 28319 17153
rect 21192 17088 21404 17116
rect 21542 17076 21548 17128
rect 21600 17116 21606 17128
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21600 17088 21925 17116
rect 21600 17076 21606 17088
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 23014 17076 23020 17128
rect 23072 17116 23078 17128
rect 23109 17119 23167 17125
rect 23109 17116 23121 17119
rect 23072 17088 23121 17116
rect 23072 17076 23078 17088
rect 23109 17085 23121 17088
rect 23155 17085 23167 17119
rect 23109 17079 23167 17085
rect 23569 17119 23627 17125
rect 23569 17085 23581 17119
rect 23615 17116 23627 17119
rect 23753 17119 23811 17125
rect 23753 17116 23765 17119
rect 23615 17088 23765 17116
rect 23615 17085 23627 17088
rect 23569 17079 23627 17085
rect 23753 17085 23765 17088
rect 23799 17085 23811 17119
rect 23753 17079 23811 17085
rect 24210 17076 24216 17128
rect 24268 17116 24274 17128
rect 25682 17116 25688 17128
rect 24268 17088 25688 17116
rect 24268 17076 24274 17088
rect 25682 17076 25688 17088
rect 25740 17116 25746 17128
rect 27062 17116 27068 17128
rect 25740 17088 27068 17116
rect 25740 17076 25746 17088
rect 27062 17076 27068 17088
rect 27120 17076 27126 17128
rect 28000 17116 28028 17147
rect 28184 17116 28212 17147
rect 28626 17144 28632 17196
rect 28684 17144 28690 17196
rect 28718 17144 28724 17196
rect 28776 17144 28782 17196
rect 28810 17144 28816 17196
rect 28868 17144 28874 17196
rect 28994 17144 29000 17196
rect 29052 17144 29058 17196
rect 31202 17144 31208 17196
rect 31260 17144 31266 17196
rect 31312 17184 31340 17224
rect 31389 17187 31447 17193
rect 31389 17184 31401 17187
rect 31312 17156 31401 17184
rect 31389 17153 31401 17156
rect 31435 17153 31447 17187
rect 31389 17147 31447 17153
rect 31570 17144 31576 17196
rect 31628 17144 31634 17196
rect 31665 17187 31723 17193
rect 31665 17153 31677 17187
rect 31711 17184 31723 17187
rect 31754 17184 31760 17196
rect 31711 17156 31760 17184
rect 31711 17153 31723 17156
rect 31665 17147 31723 17153
rect 31754 17144 31760 17156
rect 31812 17144 31818 17196
rect 32324 17193 32352 17224
rect 34333 17221 34345 17224
rect 34379 17221 34391 17255
rect 34333 17215 34391 17221
rect 31941 17187 31999 17193
rect 31941 17153 31953 17187
rect 31987 17153 31999 17187
rect 31941 17147 31999 17153
rect 32125 17187 32183 17193
rect 32125 17153 32137 17187
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32309 17187 32367 17193
rect 32309 17153 32321 17187
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 33965 17187 34023 17193
rect 33965 17153 33977 17187
rect 34011 17153 34023 17187
rect 33965 17147 34023 17153
rect 34241 17187 34299 17193
rect 34241 17153 34253 17187
rect 34287 17184 34299 17187
rect 34440 17184 34468 17280
rect 34514 17212 34520 17264
rect 34572 17261 34578 17264
rect 34572 17255 34591 17261
rect 34579 17221 34591 17255
rect 34572 17215 34591 17221
rect 34808 17252 34836 17292
rect 34808 17224 35388 17252
rect 34572 17212 34578 17215
rect 34808 17193 34836 17224
rect 34287 17156 34468 17184
rect 34287 17153 34299 17156
rect 34241 17147 34299 17153
rect 31588 17116 31616 17144
rect 31956 17116 31984 17147
rect 28000 17088 28120 17116
rect 28184 17088 28304 17116
rect 31588 17088 31984 17116
rect 20346 17008 20352 17060
rect 20404 17008 20410 17060
rect 20438 17008 20444 17060
rect 20496 17048 20502 17060
rect 20496 17020 21588 17048
rect 20496 17008 20502 17020
rect 21174 16980 21180 16992
rect 20272 16952 21180 16980
rect 21174 16940 21180 16952
rect 21232 16980 21238 16992
rect 21453 16983 21511 16989
rect 21453 16980 21465 16983
rect 21232 16952 21465 16980
rect 21232 16940 21238 16952
rect 21453 16949 21465 16952
rect 21499 16949 21511 16983
rect 21560 16980 21588 17020
rect 22646 17008 22652 17060
rect 22704 17008 22710 17060
rect 27982 17008 27988 17060
rect 28040 17008 28046 17060
rect 24118 16980 24124 16992
rect 21560 16952 24124 16980
rect 21453 16943 21511 16949
rect 24118 16940 24124 16952
rect 24176 16940 24182 16992
rect 28092 16980 28120 17088
rect 28276 17048 28304 17088
rect 31665 17051 31723 17057
rect 28276 17020 29316 17048
rect 29178 16980 29184 16992
rect 28092 16952 29184 16980
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 29288 16989 29316 17020
rect 31665 17017 31677 17051
rect 31711 17048 31723 17051
rect 32140 17048 32168 17147
rect 33980 17116 34008 17147
rect 34330 17116 34336 17128
rect 33980 17088 34336 17116
rect 34330 17076 34336 17088
rect 34388 17076 34394 17128
rect 34440 17116 34468 17156
rect 34793 17187 34851 17193
rect 34793 17153 34805 17187
rect 34839 17153 34851 17187
rect 35253 17187 35311 17193
rect 35253 17184 35265 17187
rect 34793 17147 34851 17153
rect 34992 17156 35265 17184
rect 34992 17128 35020 17156
rect 35253 17153 35265 17156
rect 35299 17153 35311 17187
rect 35253 17147 35311 17153
rect 34514 17116 34520 17128
rect 34440 17088 34520 17116
rect 34514 17076 34520 17088
rect 34572 17076 34578 17128
rect 34698 17076 34704 17128
rect 34756 17116 34762 17128
rect 34885 17119 34943 17125
rect 34885 17116 34897 17119
rect 34756 17088 34897 17116
rect 34756 17076 34762 17088
rect 34885 17085 34897 17088
rect 34931 17085 34943 17119
rect 34885 17079 34943 17085
rect 34974 17076 34980 17128
rect 35032 17076 35038 17128
rect 35360 17125 35388 17224
rect 35526 17212 35532 17264
rect 35584 17212 35590 17264
rect 35345 17119 35403 17125
rect 35345 17085 35357 17119
rect 35391 17085 35403 17119
rect 35345 17079 35403 17085
rect 35529 17119 35587 17125
rect 35529 17085 35541 17119
rect 35575 17085 35587 17119
rect 35529 17079 35587 17085
rect 31711 17020 32168 17048
rect 31711 17017 31723 17020
rect 31665 17011 31723 17017
rect 32398 17008 32404 17060
rect 32456 17008 32462 17060
rect 35161 17051 35219 17057
rect 35161 17048 35173 17051
rect 32508 17020 35173 17048
rect 29273 16983 29331 16989
rect 29273 16949 29285 16983
rect 29319 16980 29331 16983
rect 32508 16980 32536 17020
rect 35161 17017 35173 17020
rect 35207 17017 35219 17051
rect 35544 17048 35572 17079
rect 35161 17011 35219 17017
rect 35360 17020 35572 17048
rect 35360 16992 35388 17020
rect 29319 16952 32536 16980
rect 33965 16983 34023 16989
rect 29319 16949 29331 16952
rect 29273 16943 29331 16949
rect 33965 16949 33977 16983
rect 34011 16980 34023 16983
rect 34422 16980 34428 16992
rect 34011 16952 34428 16980
rect 34011 16949 34023 16952
rect 33965 16943 34023 16949
rect 34422 16940 34428 16952
rect 34480 16940 34486 16992
rect 34514 16940 34520 16992
rect 34572 16940 34578 16992
rect 34606 16940 34612 16992
rect 34664 16980 34670 16992
rect 34793 16983 34851 16989
rect 34793 16980 34805 16983
rect 34664 16952 34805 16980
rect 34664 16940 34670 16952
rect 34793 16949 34805 16952
rect 34839 16980 34851 16983
rect 34974 16980 34980 16992
rect 34839 16952 34980 16980
rect 34839 16949 34851 16952
rect 34793 16943 34851 16949
rect 34974 16940 34980 16952
rect 35032 16940 35038 16992
rect 35342 16940 35348 16992
rect 35400 16940 35406 16992
rect 1104 16890 38272 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38272 16890
rect 1104 16816 38272 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1949 16779 2007 16785
rect 1949 16776 1961 16779
rect 1728 16748 1961 16776
rect 1728 16736 1734 16748
rect 1949 16745 1961 16748
rect 1995 16745 2007 16779
rect 1949 16739 2007 16745
rect 2498 16736 2504 16788
rect 2556 16736 2562 16788
rect 3050 16736 3056 16788
rect 3108 16776 3114 16788
rect 3108 16748 5120 16776
rect 3108 16736 3114 16748
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 2516 16572 2544 16736
rect 4706 16708 4712 16720
rect 4632 16680 4712 16708
rect 4522 16600 4528 16652
rect 4580 16640 4586 16652
rect 4632 16649 4660 16680
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 5092 16708 5120 16748
rect 5166 16736 5172 16788
rect 5224 16776 5230 16788
rect 5224 16748 6914 16776
rect 5224 16736 5230 16748
rect 5534 16708 5540 16720
rect 5092 16680 5540 16708
rect 5534 16668 5540 16680
rect 5592 16668 5598 16720
rect 5810 16668 5816 16720
rect 5868 16668 5874 16720
rect 6886 16708 6914 16748
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7248 16748 10180 16776
rect 7248 16736 7254 16748
rect 6886 16680 6960 16708
rect 6932 16652 6960 16680
rect 8478 16668 8484 16720
rect 8536 16708 8542 16720
rect 8665 16711 8723 16717
rect 8665 16708 8677 16711
rect 8536 16680 8677 16708
rect 8536 16668 8542 16680
rect 8665 16677 8677 16680
rect 8711 16677 8723 16711
rect 8665 16671 8723 16677
rect 4617 16643 4675 16649
rect 4617 16640 4629 16643
rect 4580 16612 4629 16640
rect 4580 16600 4586 16612
rect 4617 16609 4629 16612
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 5077 16643 5135 16649
rect 5077 16609 5089 16643
rect 5123 16640 5135 16643
rect 6273 16643 6331 16649
rect 6273 16640 6285 16643
rect 5123 16612 6285 16640
rect 5123 16609 5135 16612
rect 5077 16603 5135 16609
rect 6273 16609 6285 16612
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 6457 16643 6515 16649
rect 6457 16609 6469 16643
rect 6503 16640 6515 16643
rect 6730 16640 6736 16652
rect 6503 16612 6736 16640
rect 6503 16609 6515 16612
rect 6457 16603 6515 16609
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 6914 16600 6920 16652
rect 6972 16600 6978 16652
rect 9125 16643 9183 16649
rect 9125 16609 9137 16643
rect 9171 16640 9183 16643
rect 9214 16640 9220 16652
rect 9171 16612 9220 16640
rect 9171 16609 9183 16612
rect 9125 16603 9183 16609
rect 9214 16600 9220 16612
rect 9272 16640 9278 16652
rect 10042 16640 10048 16652
rect 9272 16612 10048 16640
rect 9272 16600 9278 16612
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 10152 16640 10180 16748
rect 15378 16736 15384 16788
rect 15436 16776 15442 16788
rect 16482 16776 16488 16788
rect 15436 16748 16488 16776
rect 15436 16736 15442 16748
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 20438 16776 20444 16788
rect 18196 16748 18736 16776
rect 18196 16736 18202 16748
rect 18708 16717 18736 16748
rect 19168 16748 20444 16776
rect 18693 16711 18751 16717
rect 12406 16680 17540 16708
rect 12406 16640 12434 16680
rect 10152 16612 12434 16640
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 13081 16643 13139 16649
rect 13081 16640 13093 16643
rect 12860 16612 13093 16640
rect 12860 16600 12866 16612
rect 13081 16609 13093 16612
rect 13127 16609 13139 16643
rect 13722 16640 13728 16652
rect 13081 16603 13139 16609
rect 13188 16612 13728 16640
rect 2179 16544 2544 16572
rect 4709 16575 4767 16581
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 4798 16572 4804 16584
rect 4755 16544 4804 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 8294 16532 8300 16584
rect 8352 16532 8358 16584
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 9309 16575 9367 16581
rect 9309 16572 9321 16575
rect 9088 16544 9321 16572
rect 9088 16532 9094 16544
rect 9309 16541 9321 16544
rect 9355 16572 9367 16575
rect 9490 16572 9496 16584
rect 9355 16544 9496 16572
rect 9355 16541 9367 16544
rect 9309 16535 9367 16541
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16572 13047 16575
rect 13188 16572 13216 16612
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14366 16600 14372 16652
rect 14424 16600 14430 16652
rect 15470 16640 15476 16652
rect 14752 16612 15476 16640
rect 14752 16581 14780 16612
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 17512 16640 17540 16680
rect 18064 16680 18644 16708
rect 18064 16649 18092 16680
rect 18049 16643 18107 16649
rect 17512 16612 18000 16640
rect 13035 16544 13216 16572
rect 14461 16575 14519 16581
rect 13035 16541 13047 16544
rect 12989 16535 13047 16541
rect 14461 16541 14473 16575
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 14737 16575 14795 16581
rect 14737 16541 14749 16575
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 7190 16464 7196 16516
rect 7248 16464 7254 16516
rect 13078 16464 13084 16516
rect 13136 16464 13142 16516
rect 6178 16396 6184 16448
rect 6236 16396 6242 16448
rect 9122 16396 9128 16448
rect 9180 16436 9186 16448
rect 9398 16436 9404 16448
rect 9180 16408 9404 16436
rect 9180 16396 9186 16408
rect 9398 16396 9404 16408
rect 9456 16436 9462 16448
rect 9493 16439 9551 16445
rect 9493 16436 9505 16439
rect 9456 16408 9505 16436
rect 9456 16396 9462 16408
rect 9493 16405 9505 16408
rect 9539 16405 9551 16439
rect 9493 16399 9551 16405
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 12529 16439 12587 16445
rect 12529 16436 12541 16439
rect 9640 16408 12541 16436
rect 9640 16396 9646 16408
rect 12529 16405 12541 16408
rect 12575 16405 12587 16439
rect 12529 16399 12587 16405
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 12894 16436 12900 16448
rect 12676 16408 12900 16436
rect 12676 16396 12682 16408
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 13096 16436 13124 16464
rect 14476 16448 14504 16535
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 16482 16572 16488 16584
rect 15344 16544 16488 16572
rect 15344 16532 15350 16544
rect 16482 16532 16488 16544
rect 16540 16572 16546 16584
rect 16758 16572 16764 16584
rect 16540 16544 16764 16572
rect 16540 16532 16546 16544
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17972 16572 18000 16612
rect 18049 16609 18061 16643
rect 18095 16609 18107 16643
rect 18049 16603 18107 16609
rect 18141 16643 18199 16649
rect 18141 16609 18153 16643
rect 18187 16640 18199 16643
rect 18506 16640 18512 16652
rect 18187 16612 18512 16640
rect 18187 16609 18199 16612
rect 18141 16603 18199 16609
rect 18156 16572 18184 16603
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 18616 16640 18644 16680
rect 18693 16677 18705 16711
rect 18739 16677 18751 16711
rect 18693 16671 18751 16677
rect 19168 16640 19196 16748
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 20530 16736 20536 16788
rect 20588 16776 20594 16788
rect 20990 16776 20996 16788
rect 20588 16748 20996 16776
rect 20588 16736 20594 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21174 16736 21180 16788
rect 21232 16736 21238 16788
rect 26878 16776 26884 16788
rect 22480 16748 26884 16776
rect 19610 16668 19616 16720
rect 19668 16708 19674 16720
rect 20346 16708 20352 16720
rect 19668 16680 20352 16708
rect 19668 16668 19674 16680
rect 20346 16668 20352 16680
rect 20404 16668 20410 16720
rect 22480 16708 22508 16748
rect 26878 16736 26884 16748
rect 26936 16736 26942 16788
rect 32398 16776 32404 16788
rect 28966 16748 32404 16776
rect 20457 16680 22508 16708
rect 22557 16711 22615 16717
rect 18616 16612 19196 16640
rect 19245 16643 19303 16649
rect 19245 16609 19257 16643
rect 19291 16640 19303 16643
rect 20457 16640 20485 16680
rect 22557 16677 22569 16711
rect 22603 16708 22615 16711
rect 24946 16708 24952 16720
rect 22603 16680 24952 16708
rect 22603 16677 22615 16680
rect 22557 16671 22615 16677
rect 24946 16668 24952 16680
rect 25004 16668 25010 16720
rect 28966 16708 28994 16748
rect 32398 16736 32404 16748
rect 32456 16736 32462 16788
rect 34698 16736 34704 16788
rect 34756 16776 34762 16788
rect 35161 16779 35219 16785
rect 35161 16776 35173 16779
rect 34756 16748 35173 16776
rect 34756 16736 34762 16748
rect 35161 16745 35173 16748
rect 35207 16776 35219 16779
rect 35342 16776 35348 16788
rect 35207 16748 35348 16776
rect 35207 16745 35219 16748
rect 35161 16739 35219 16745
rect 35342 16736 35348 16748
rect 35400 16736 35406 16788
rect 25056 16680 28994 16708
rect 19291 16612 20485 16640
rect 19291 16609 19303 16612
rect 19245 16603 19303 16609
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 22813 16643 22871 16649
rect 22813 16640 22825 16643
rect 20588 16612 22825 16640
rect 20588 16600 20594 16612
rect 22813 16609 22825 16612
rect 22859 16609 22871 16643
rect 22813 16603 22871 16609
rect 17972 16544 18184 16572
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 18782 16572 18788 16584
rect 18463 16544 18788 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 18782 16532 18788 16544
rect 18840 16572 18846 16584
rect 19058 16572 19064 16584
rect 18840 16544 19064 16572
rect 18840 16532 18846 16544
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 19705 16575 19763 16581
rect 19705 16572 19717 16575
rect 19484 16544 19717 16572
rect 19484 16532 19490 16544
rect 19705 16541 19717 16544
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 19852 16544 19901 16572
rect 19852 16532 19858 16544
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20073 16575 20131 16581
rect 20073 16572 20085 16575
rect 20036 16544 20085 16572
rect 20036 16532 20042 16544
rect 20073 16541 20085 16544
rect 20119 16541 20131 16575
rect 20073 16535 20131 16541
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 15654 16504 15660 16516
rect 14884 16476 15660 16504
rect 14884 16464 14890 16476
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 17328 16476 17908 16504
rect 17328 16448 17356 16476
rect 14185 16439 14243 16445
rect 14185 16436 14197 16439
rect 13096 16408 14197 16436
rect 14185 16405 14197 16408
rect 14231 16405 14243 16439
rect 14185 16399 14243 16405
rect 14458 16396 14464 16448
rect 14516 16396 14522 16448
rect 14550 16396 14556 16448
rect 14608 16436 14614 16448
rect 17310 16436 17316 16448
rect 14608 16408 17316 16436
rect 14608 16396 14614 16408
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 17586 16396 17592 16448
rect 17644 16396 17650 16448
rect 17880 16436 17908 16476
rect 17954 16464 17960 16516
rect 18012 16464 18018 16516
rect 19610 16504 19616 16516
rect 18801 16476 19616 16504
rect 18801 16436 18829 16476
rect 19610 16464 19616 16476
rect 19668 16464 19674 16516
rect 17880 16408 18829 16436
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 20088 16436 20116 16535
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 20496 16544 20637 16572
rect 20496 16532 20502 16544
rect 20625 16541 20637 16544
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20772 16544 20852 16572
rect 20772 16532 20778 16544
rect 20824 16513 20852 16544
rect 21174 16532 21180 16584
rect 21232 16572 21238 16584
rect 21453 16575 21511 16581
rect 21453 16572 21465 16575
rect 21232 16544 21465 16572
rect 21232 16532 21238 16544
rect 21453 16541 21465 16544
rect 21499 16541 21511 16575
rect 22828 16572 22856 16603
rect 23106 16600 23112 16652
rect 23164 16600 23170 16652
rect 24118 16600 24124 16652
rect 24176 16640 24182 16652
rect 25056 16640 25084 16680
rect 24176 16612 25084 16640
rect 24176 16600 24182 16612
rect 27246 16600 27252 16652
rect 27304 16640 27310 16652
rect 28626 16640 28632 16652
rect 27304 16612 28632 16640
rect 27304 16600 27310 16612
rect 28626 16600 28632 16612
rect 28684 16640 28690 16652
rect 32490 16640 32496 16652
rect 28684 16612 32496 16640
rect 28684 16600 28690 16612
rect 32490 16600 32496 16612
rect 32548 16600 32554 16652
rect 34790 16600 34796 16652
rect 34848 16600 34854 16652
rect 25866 16572 25872 16584
rect 21453 16535 21511 16541
rect 21560 16544 22692 16572
rect 22828 16544 25872 16572
rect 20809 16507 20867 16513
rect 20809 16473 20821 16507
rect 20855 16473 20867 16507
rect 20809 16467 20867 16473
rect 21025 16507 21083 16513
rect 21025 16473 21037 16507
rect 21071 16504 21083 16507
rect 21266 16504 21272 16516
rect 21071 16476 21272 16504
rect 21071 16473 21083 16476
rect 21025 16467 21083 16473
rect 21266 16464 21272 16476
rect 21324 16464 21330 16516
rect 21560 16436 21588 16544
rect 22002 16464 22008 16516
rect 22060 16464 22066 16516
rect 22554 16464 22560 16516
rect 22612 16464 22618 16516
rect 22664 16504 22692 16544
rect 25866 16532 25872 16544
rect 25924 16532 25930 16584
rect 31205 16575 31263 16581
rect 31205 16541 31217 16575
rect 31251 16572 31263 16575
rect 32122 16572 32128 16584
rect 31251 16544 32128 16572
rect 31251 16541 31263 16544
rect 31205 16535 31263 16541
rect 32122 16532 32128 16544
rect 32180 16532 32186 16584
rect 33318 16532 33324 16584
rect 33376 16572 33382 16584
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 33376 16544 34897 16572
rect 33376 16532 33382 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 23017 16507 23075 16513
rect 23017 16504 23029 16507
rect 22664 16476 23029 16504
rect 23017 16473 23029 16476
rect 23063 16504 23075 16507
rect 24854 16504 24860 16516
rect 23063 16476 24860 16504
rect 23063 16473 23075 16476
rect 23017 16467 23075 16473
rect 24854 16464 24860 16476
rect 24912 16464 24918 16516
rect 20088 16408 21588 16436
rect 22922 16396 22928 16448
rect 22980 16396 22986 16448
rect 30374 16396 30380 16448
rect 30432 16436 30438 16448
rect 31389 16439 31447 16445
rect 31389 16436 31401 16439
rect 30432 16408 31401 16436
rect 30432 16396 30438 16408
rect 31389 16405 31401 16408
rect 31435 16405 31447 16439
rect 31389 16399 31447 16405
rect 1104 16346 38272 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38272 16346
rect 1104 16272 38272 16294
rect 3988 16204 4844 16232
rect 1486 16124 1492 16176
rect 1544 16124 1550 16176
rect 3988 16108 4016 16204
rect 4709 16167 4767 16173
rect 4709 16164 4721 16167
rect 4356 16136 4721 16164
rect 3970 16056 3976 16108
rect 4028 16056 4034 16108
rect 4062 16056 4068 16108
rect 4120 16056 4126 16108
rect 4356 16105 4384 16136
rect 4709 16133 4721 16136
rect 4755 16133 4767 16167
rect 4709 16127 4767 16133
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 4522 16056 4528 16108
rect 4580 16056 4586 16108
rect 4816 16105 4844 16204
rect 6178 16192 6184 16244
rect 6236 16192 6242 16244
rect 7190 16192 7196 16244
rect 7248 16232 7254 16244
rect 7653 16235 7711 16241
rect 7653 16232 7665 16235
rect 7248 16204 7665 16232
rect 7248 16192 7254 16204
rect 7653 16201 7665 16204
rect 7699 16201 7711 16235
rect 7653 16195 7711 16201
rect 8478 16192 8484 16244
rect 8536 16192 8542 16244
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 15197 16235 15255 16241
rect 15197 16232 15209 16235
rect 8628 16204 15209 16232
rect 8628 16192 8634 16204
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 992 15864 1593 15892
rect 992 15852 998 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 4080 15892 4108 16056
rect 4249 16031 4307 16037
rect 4249 15997 4261 16031
rect 4295 16028 4307 16031
rect 4540 16028 4568 16056
rect 4295 16000 4568 16028
rect 4632 16028 4660 16059
rect 4632 16000 4844 16028
rect 4295 15997 4307 16000
rect 4249 15991 4307 15997
rect 4341 15963 4399 15969
rect 4341 15929 4353 15963
rect 4387 15960 4399 15963
rect 4706 15960 4712 15972
rect 4387 15932 4712 15960
rect 4387 15929 4399 15932
rect 4341 15923 4399 15929
rect 4706 15920 4712 15932
rect 4764 15920 4770 15972
rect 4816 15892 4844 16000
rect 4080 15864 4844 15892
rect 6196 15892 6224 16192
rect 6822 16124 6828 16176
rect 6880 16164 6886 16176
rect 6880 16136 9536 16164
rect 6880 16124 6886 16136
rect 7837 16099 7895 16105
rect 7837 16096 7849 16099
rect 7484 16068 7849 16096
rect 7484 15960 7512 16068
rect 7837 16065 7849 16068
rect 7883 16065 7895 16099
rect 7837 16059 7895 16065
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16096 8447 16099
rect 9122 16096 9128 16108
rect 8435 16068 9128 16096
rect 8435 16065 8447 16068
rect 8389 16059 8447 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9306 16056 9312 16108
rect 9364 16056 9370 16108
rect 9508 16105 9536 16136
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9493 16099 9551 16105
rect 9493 16065 9505 16099
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 8662 15988 8668 16040
rect 8720 15988 8726 16040
rect 9416 16028 9444 16059
rect 8956 16000 9444 16028
rect 8021 15963 8079 15969
rect 8021 15960 8033 15963
rect 7484 15932 8033 15960
rect 8021 15929 8033 15932
rect 8067 15929 8079 15963
rect 8021 15923 8079 15929
rect 8478 15920 8484 15972
rect 8536 15960 8542 15972
rect 8754 15960 8760 15972
rect 8536 15932 8760 15960
rect 8536 15920 8542 15932
rect 8754 15920 8760 15932
rect 8812 15960 8818 15972
rect 8956 15960 8984 16000
rect 8812 15932 8984 15960
rect 8812 15920 8818 15932
rect 9030 15920 9036 15972
rect 9088 15920 9094 15972
rect 9122 15920 9128 15972
rect 9180 15960 9186 15972
rect 9600 15960 9628 16204
rect 15197 16201 15209 16204
rect 15243 16201 15255 16235
rect 18874 16232 18880 16244
rect 15197 16195 15255 16201
rect 16132 16204 18880 16232
rect 12158 16124 12164 16176
rect 12216 16164 12222 16176
rect 12216 16136 13860 16164
rect 12216 16124 12222 16136
rect 9674 16056 9680 16108
rect 9732 16056 9738 16108
rect 12986 16056 12992 16108
rect 13044 16056 13050 16108
rect 13832 16096 13860 16136
rect 13906 16124 13912 16176
rect 13964 16124 13970 16176
rect 16132 16105 16160 16204
rect 18874 16192 18880 16204
rect 18932 16192 18938 16244
rect 30098 16192 30104 16244
rect 30156 16192 30162 16244
rect 34330 16192 34336 16244
rect 34388 16192 34394 16244
rect 16942 16124 16948 16176
rect 17000 16124 17006 16176
rect 17236 16136 17540 16164
rect 17236 16105 17264 16136
rect 17512 16108 17540 16136
rect 17880 16136 19334 16164
rect 17880 16108 17908 16136
rect 16117 16099 16175 16105
rect 16117 16096 16129 16099
rect 13832 16068 16129 16096
rect 16117 16065 16129 16068
rect 16163 16065 16175 16099
rect 16117 16059 16175 16065
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 12802 15988 12808 16040
rect 12860 15988 12866 16040
rect 13078 15988 13084 16040
rect 13136 15988 13142 16040
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 15997 13231 16031
rect 13173 15991 13231 15997
rect 12621 15963 12679 15969
rect 12621 15960 12633 15963
rect 9180 15932 9628 15960
rect 12406 15932 12633 15960
rect 9180 15920 9186 15932
rect 12406 15892 12434 15932
rect 12621 15929 12633 15932
rect 12667 15929 12679 15963
rect 12820 15960 12848 15988
rect 13188 15960 13216 15991
rect 16022 15988 16028 16040
rect 16080 16028 16086 16040
rect 16206 16028 16212 16040
rect 16080 16000 16212 16028
rect 16080 15988 16086 16000
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 17328 16028 17356 16059
rect 16500 16000 17356 16028
rect 16500 15969 16528 16000
rect 16485 15963 16543 15969
rect 12820 15932 16344 15960
rect 12621 15923 12679 15929
rect 6196 15864 12434 15892
rect 1581 15855 1639 15861
rect 16206 15852 16212 15904
rect 16264 15852 16270 15904
rect 16316 15892 16344 15932
rect 16485 15929 16497 15963
rect 16531 15929 16543 15963
rect 16485 15923 16543 15929
rect 16850 15920 16856 15972
rect 16908 15960 16914 15972
rect 17420 15960 17448 16059
rect 17494 16056 17500 16108
rect 17552 16056 17558 16108
rect 17589 16099 17647 16105
rect 17589 16065 17601 16099
rect 17635 16096 17647 16099
rect 17678 16096 17684 16108
rect 17635 16068 17684 16096
rect 17635 16065 17647 16068
rect 17589 16059 17647 16065
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 17770 16056 17776 16108
rect 17828 16056 17834 16108
rect 17862 16056 17868 16108
rect 17920 16056 17926 16108
rect 18966 16056 18972 16108
rect 19024 16056 19030 16108
rect 19306 16096 19334 16136
rect 20622 16124 20628 16176
rect 20680 16164 20686 16176
rect 20809 16167 20867 16173
rect 20809 16164 20821 16167
rect 20680 16136 20821 16164
rect 20680 16124 20686 16136
rect 20809 16133 20821 16136
rect 20855 16133 20867 16167
rect 20809 16127 20867 16133
rect 24964 16136 26556 16164
rect 24964 16108 24992 16136
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19306 16068 19901 16096
rect 19889 16065 19901 16068
rect 19935 16096 19947 16099
rect 20438 16096 20444 16108
rect 19935 16068 20444 16096
rect 19935 16065 19947 16068
rect 19889 16059 19947 16065
rect 20438 16056 20444 16068
rect 20496 16096 20502 16108
rect 20898 16096 20904 16108
rect 20496 16068 20904 16096
rect 20496 16056 20502 16068
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 24302 16056 24308 16108
rect 24360 16056 24366 16108
rect 24578 16056 24584 16108
rect 24636 16096 24642 16108
rect 24857 16099 24915 16105
rect 24857 16096 24869 16099
rect 24636 16068 24869 16096
rect 24636 16056 24642 16068
rect 24857 16065 24869 16068
rect 24903 16065 24915 16099
rect 24857 16059 24915 16065
rect 24872 16028 24900 16059
rect 24946 16056 24952 16108
rect 25004 16056 25010 16108
rect 25130 16056 25136 16108
rect 25188 16096 25194 16108
rect 26528 16105 26556 16136
rect 27154 16124 27160 16176
rect 27212 16164 27218 16176
rect 29362 16164 29368 16176
rect 27212 16136 29368 16164
rect 27212 16124 27218 16136
rect 29362 16124 29368 16136
rect 29420 16164 29426 16176
rect 30377 16167 30435 16173
rect 30377 16164 30389 16167
rect 29420 16136 29868 16164
rect 29420 16124 29426 16136
rect 25593 16099 25651 16105
rect 25593 16096 25605 16099
rect 25188 16068 25605 16096
rect 25188 16056 25194 16068
rect 25593 16065 25605 16068
rect 25639 16096 25651 16099
rect 25869 16099 25927 16105
rect 25869 16096 25881 16099
rect 25639 16068 25881 16096
rect 25639 16065 25651 16068
rect 25593 16059 25651 16065
rect 25869 16065 25881 16068
rect 25915 16065 25927 16099
rect 25869 16059 25927 16065
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16065 26111 16099
rect 26053 16059 26111 16065
rect 26513 16099 26571 16105
rect 26513 16065 26525 16099
rect 26559 16065 26571 16099
rect 26513 16059 26571 16065
rect 25409 16031 25467 16037
rect 25409 16028 25421 16031
rect 24872 16000 25421 16028
rect 25409 15997 25421 16000
rect 25455 16028 25467 16031
rect 26068 16028 26096 16059
rect 29086 16056 29092 16108
rect 29144 16096 29150 16108
rect 29840 16105 29868 16136
rect 30024 16136 30389 16164
rect 30024 16105 30052 16136
rect 30377 16133 30389 16136
rect 30423 16133 30435 16167
rect 30377 16127 30435 16133
rect 29181 16099 29239 16105
rect 29181 16096 29193 16099
rect 29144 16068 29193 16096
rect 29144 16056 29150 16068
rect 29181 16065 29193 16068
rect 29227 16096 29239 16099
rect 29641 16099 29699 16105
rect 29641 16096 29653 16099
rect 29227 16068 29653 16096
rect 29227 16065 29239 16068
rect 29181 16059 29239 16065
rect 29641 16065 29653 16068
rect 29687 16065 29699 16099
rect 29641 16059 29699 16065
rect 29825 16099 29883 16105
rect 29825 16065 29837 16099
rect 29871 16065 29883 16099
rect 29825 16059 29883 16065
rect 30009 16099 30067 16105
rect 30009 16065 30021 16099
rect 30055 16065 30067 16099
rect 30009 16059 30067 16065
rect 30193 16099 30251 16105
rect 30193 16065 30205 16099
rect 30239 16096 30251 16099
rect 30282 16096 30288 16108
rect 30239 16068 30288 16096
rect 30239 16065 30251 16068
rect 30193 16059 30251 16065
rect 30282 16056 30288 16068
rect 30340 16056 30346 16108
rect 30561 16099 30619 16105
rect 30561 16065 30573 16099
rect 30607 16065 30619 16099
rect 30561 16059 30619 16065
rect 30745 16099 30803 16105
rect 30745 16065 30757 16099
rect 30791 16065 30803 16099
rect 30745 16059 30803 16065
rect 30837 16099 30895 16105
rect 30837 16065 30849 16099
rect 30883 16096 30895 16099
rect 32858 16096 32864 16108
rect 30883 16068 32864 16096
rect 30883 16065 30895 16068
rect 30837 16059 30895 16065
rect 25455 16000 26096 16028
rect 25455 15997 25467 16000
rect 25409 15991 25467 15997
rect 26234 15988 26240 16040
rect 26292 16028 26298 16040
rect 26329 16031 26387 16037
rect 26329 16028 26341 16031
rect 26292 16000 26341 16028
rect 26292 15988 26298 16000
rect 26329 15997 26341 16000
rect 26375 15997 26387 16031
rect 26329 15991 26387 15997
rect 26418 15988 26424 16040
rect 26476 16028 26482 16040
rect 26697 16031 26755 16037
rect 26697 16028 26709 16031
rect 26476 16000 26709 16028
rect 26476 15988 26482 16000
rect 26697 15997 26709 16000
rect 26743 16028 26755 16031
rect 30576 16028 30604 16059
rect 26743 16000 30604 16028
rect 26743 15997 26755 16000
rect 26697 15991 26755 15997
rect 30760 15972 30788 16059
rect 32858 16056 32864 16068
rect 32916 16056 32922 16108
rect 33962 16056 33968 16108
rect 34020 16056 34026 16108
rect 37642 16056 37648 16108
rect 37700 16056 37706 16108
rect 33870 15988 33876 16040
rect 33928 15988 33934 16040
rect 20622 15960 20628 15972
rect 16908 15932 20628 15960
rect 16908 15920 16914 15932
rect 20622 15920 20628 15932
rect 20680 15920 20686 15972
rect 25777 15963 25835 15969
rect 25777 15929 25789 15963
rect 25823 15960 25835 15963
rect 26510 15960 26516 15972
rect 25823 15932 26516 15960
rect 25823 15929 25835 15932
rect 25777 15923 25835 15929
rect 26510 15920 26516 15932
rect 26568 15920 26574 15972
rect 26878 15920 26884 15972
rect 26936 15960 26942 15972
rect 27890 15960 27896 15972
rect 26936 15932 27896 15960
rect 26936 15920 26942 15932
rect 27890 15920 27896 15932
rect 27948 15920 27954 15972
rect 30374 15920 30380 15972
rect 30432 15960 30438 15972
rect 30742 15960 30748 15972
rect 30432 15932 30748 15960
rect 30432 15920 30438 15932
rect 30742 15920 30748 15932
rect 30800 15920 30806 15972
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 16316 15864 17877 15892
rect 17865 15861 17877 15864
rect 17911 15892 17923 15895
rect 18690 15892 18696 15904
rect 17911 15864 18696 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 18690 15852 18696 15864
rect 18748 15852 18754 15904
rect 24397 15895 24455 15901
rect 24397 15861 24409 15895
rect 24443 15892 24455 15895
rect 24670 15892 24676 15904
rect 24443 15864 24676 15892
rect 24443 15861 24455 15864
rect 24397 15855 24455 15861
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 25961 15895 26019 15901
rect 25961 15861 25973 15895
rect 26007 15892 26019 15895
rect 27154 15892 27160 15904
rect 26007 15864 27160 15892
rect 26007 15861 26019 15864
rect 25961 15855 26019 15861
rect 27154 15852 27160 15864
rect 27212 15852 27218 15904
rect 29546 15852 29552 15904
rect 29604 15852 29610 15904
rect 29733 15895 29791 15901
rect 29733 15861 29745 15895
rect 29779 15892 29791 15895
rect 29822 15892 29828 15904
rect 29779 15864 29828 15892
rect 29779 15861 29791 15864
rect 29733 15855 29791 15861
rect 29822 15852 29828 15864
rect 29880 15852 29886 15904
rect 37826 15852 37832 15904
rect 37884 15852 37890 15904
rect 1104 15802 38272 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38272 15802
rect 1104 15728 38272 15750
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 3145 15691 3203 15697
rect 3145 15688 3157 15691
rect 3016 15660 3157 15688
rect 3016 15648 3022 15660
rect 3145 15657 3157 15660
rect 3191 15688 3203 15691
rect 3970 15688 3976 15700
rect 3191 15660 3976 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4706 15648 4712 15700
rect 4764 15648 4770 15700
rect 6730 15648 6736 15700
rect 6788 15648 6794 15700
rect 9582 15688 9588 15700
rect 6840 15660 9588 15688
rect 4724 15620 4752 15648
rect 4264 15592 4752 15620
rect 1394 15512 1400 15564
rect 1452 15512 1458 15564
rect 4264 15561 4292 15592
rect 4249 15555 4307 15561
rect 4249 15521 4261 15555
rect 4295 15521 4307 15555
rect 4249 15515 4307 15521
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4614 15552 4620 15564
rect 4479 15524 4620 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4614 15512 4620 15524
rect 4672 15552 4678 15564
rect 6748 15552 6776 15648
rect 4672 15524 6776 15552
rect 4672 15512 4678 15524
rect 2774 15444 2780 15496
rect 2832 15444 2838 15496
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 6840 15484 6868 15660
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 13817 15691 13875 15697
rect 13817 15657 13829 15691
rect 13863 15688 13875 15691
rect 14550 15688 14556 15700
rect 13863 15660 14556 15688
rect 13863 15657 13875 15660
rect 13817 15651 13875 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 14734 15648 14740 15700
rect 14792 15688 14798 15700
rect 16393 15691 16451 15697
rect 16393 15688 16405 15691
rect 14792 15660 16405 15688
rect 14792 15648 14798 15660
rect 16393 15657 16405 15660
rect 16439 15688 16451 15691
rect 17126 15688 17132 15700
rect 16439 15660 17132 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 17313 15691 17371 15697
rect 17313 15657 17325 15691
rect 17359 15688 17371 15691
rect 17402 15688 17408 15700
rect 17359 15660 17408 15688
rect 17359 15657 17371 15660
rect 17313 15651 17371 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 17497 15691 17555 15697
rect 17497 15657 17509 15691
rect 17543 15688 17555 15691
rect 17770 15688 17776 15700
rect 17543 15660 17776 15688
rect 17543 15657 17555 15660
rect 17497 15651 17555 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 18046 15648 18052 15700
rect 18104 15688 18110 15700
rect 19337 15691 19395 15697
rect 19337 15688 19349 15691
rect 18104 15660 19349 15688
rect 18104 15648 18110 15660
rect 19337 15657 19349 15660
rect 19383 15688 19395 15691
rect 20898 15688 20904 15700
rect 19383 15660 20904 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 20898 15648 20904 15660
rect 20956 15688 20962 15700
rect 21542 15688 21548 15700
rect 20956 15660 21548 15688
rect 20956 15648 20962 15660
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 22554 15688 22560 15700
rect 22066 15660 22560 15688
rect 12805 15623 12863 15629
rect 12805 15589 12817 15623
rect 12851 15620 12863 15623
rect 12986 15620 12992 15632
rect 12851 15592 12992 15620
rect 12851 15589 12863 15592
rect 12805 15583 12863 15589
rect 12986 15580 12992 15592
rect 13044 15620 13050 15632
rect 22066 15620 22094 15660
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 25130 15648 25136 15700
rect 25188 15688 25194 15700
rect 26329 15691 26387 15697
rect 26329 15688 26341 15691
rect 25188 15660 26341 15688
rect 25188 15648 25194 15660
rect 26329 15657 26341 15660
rect 26375 15688 26387 15691
rect 26375 15660 27568 15688
rect 26375 15657 26387 15660
rect 26329 15651 26387 15657
rect 13044 15592 16804 15620
rect 13044 15580 13050 15592
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 6932 15524 8953 15552
rect 6932 15496 6960 15524
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9364 15524 12572 15552
rect 9364 15512 9370 15524
rect 4203 15456 6868 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 6914 15444 6920 15496
rect 6972 15444 6978 15496
rect 8754 15444 8760 15496
rect 8812 15444 8818 15496
rect 10336 15470 10364 15524
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 1670 15376 1676 15428
rect 1728 15376 1734 15428
rect 9217 15419 9275 15425
rect 9217 15385 9229 15419
rect 9263 15385 9275 15419
rect 9217 15379 9275 15385
rect 10965 15419 11023 15425
rect 10965 15385 10977 15419
rect 11011 15385 11023 15419
rect 10965 15379 11023 15385
rect 3786 15308 3792 15360
rect 3844 15308 3850 15360
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15348 8631 15351
rect 9232 15348 9260 15379
rect 8619 15320 9260 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10980 15348 11008 15379
rect 11330 15376 11336 15428
rect 11388 15376 11394 15428
rect 12544 15416 12572 15524
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 14734 15552 14740 15564
rect 14516 15524 14740 15552
rect 14516 15512 14522 15524
rect 14734 15512 14740 15524
rect 14792 15512 14798 15564
rect 15010 15512 15016 15564
rect 15068 15512 15074 15564
rect 15470 15512 15476 15564
rect 15528 15512 15534 15564
rect 16206 15552 16212 15564
rect 15672 15524 16212 15552
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 15672 15493 15700 15524
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16482 15512 16488 15564
rect 16540 15552 16546 15564
rect 16776 15552 16804 15592
rect 17420 15592 22094 15620
rect 17420 15552 17448 15592
rect 24394 15580 24400 15632
rect 24452 15620 24458 15632
rect 26418 15620 26424 15632
rect 24452 15592 26424 15620
rect 24452 15580 24458 15592
rect 26418 15580 26424 15592
rect 26476 15580 26482 15632
rect 26789 15623 26847 15629
rect 26789 15589 26801 15623
rect 26835 15589 26847 15623
rect 26789 15583 26847 15589
rect 16540 15524 16712 15552
rect 16776 15524 17448 15552
rect 16540 15512 16546 15524
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 13320 15456 13461 15484
rect 13320 15444 13326 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15453 14427 15487
rect 14369 15447 14427 15453
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 13078 15416 13084 15428
rect 12544 15402 13084 15416
rect 12558 15388 13084 15402
rect 13078 15376 13084 15388
rect 13136 15376 13142 15428
rect 11974 15348 11980 15360
rect 10008 15320 11980 15348
rect 10008 15308 10014 15320
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 13648 15348 13676 15447
rect 14384 15360 14412 15447
rect 14660 15416 14688 15447
rect 15838 15444 15844 15496
rect 15896 15444 15902 15496
rect 16684 15493 16712 15524
rect 18874 15512 18880 15564
rect 18932 15552 18938 15564
rect 20990 15552 20996 15564
rect 18932 15524 20996 15552
rect 18932 15512 18938 15524
rect 20990 15512 20996 15524
rect 21048 15552 21054 15564
rect 21048 15524 21128 15552
rect 21048 15512 21054 15524
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 16669 15487 16727 15493
rect 16669 15453 16681 15487
rect 16715 15453 16727 15487
rect 16669 15447 16727 15453
rect 16761 15487 16819 15493
rect 16761 15453 16773 15487
rect 16807 15484 16819 15487
rect 16850 15484 16856 15496
rect 16807 15456 16856 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 14660 15388 15700 15416
rect 15672 15360 15700 15388
rect 12952 15320 13676 15348
rect 12952 15308 12958 15320
rect 14366 15308 14372 15360
rect 14424 15308 14430 15360
rect 15654 15308 15660 15360
rect 15712 15308 15718 15360
rect 15838 15308 15844 15360
rect 15896 15348 15902 15360
rect 15948 15348 15976 15447
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18966 15484 18972 15496
rect 18104 15456 18972 15484
rect 18104 15444 18110 15456
rect 18966 15444 18972 15456
rect 19024 15484 19030 15496
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 19024 15456 19349 15484
rect 19024 15444 19030 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 19337 15447 19395 15453
rect 20438 15444 20444 15496
rect 20496 15444 20502 15496
rect 20622 15444 20628 15496
rect 20680 15444 20686 15496
rect 20898 15444 20904 15496
rect 20956 15444 20962 15496
rect 21100 15493 21128 15524
rect 21910 15512 21916 15564
rect 21968 15552 21974 15564
rect 26804 15552 26832 15583
rect 26878 15580 26884 15632
rect 26936 15580 26942 15632
rect 27154 15580 27160 15632
rect 27212 15580 27218 15632
rect 27172 15552 27200 15580
rect 21968 15524 22692 15552
rect 21968 15512 21974 15524
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15484 21235 15487
rect 21266 15484 21272 15496
rect 21223 15456 21272 15484
rect 21223 15453 21235 15456
rect 21177 15447 21235 15453
rect 21266 15444 21272 15456
rect 21324 15444 21330 15496
rect 21928 15484 21956 15512
rect 22664 15493 22692 15524
rect 22940 15524 23612 15552
rect 26804 15524 27200 15552
rect 22940 15493 22968 15524
rect 23584 15496 23612 15524
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 21928 15456 22017 15484
rect 22005 15453 22017 15456
rect 22051 15453 22063 15487
rect 22373 15487 22431 15493
rect 22373 15484 22385 15487
rect 22005 15447 22063 15453
rect 22112 15456 22385 15484
rect 16114 15376 16120 15428
rect 16172 15376 16178 15428
rect 16298 15376 16304 15428
rect 16356 15416 16362 15428
rect 17129 15419 17187 15425
rect 17129 15416 17141 15419
rect 16356 15388 17141 15416
rect 16356 15376 16362 15388
rect 17129 15385 17141 15388
rect 17175 15416 17187 15419
rect 17770 15416 17776 15428
rect 17175 15388 17776 15416
rect 17175 15385 17187 15388
rect 17129 15379 17187 15385
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 20640 15416 20668 15444
rect 22112 15416 22140 15456
rect 22373 15453 22385 15456
rect 22419 15453 22431 15487
rect 22373 15447 22431 15453
rect 22649 15487 22707 15493
rect 22649 15453 22661 15487
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 20640 15388 22140 15416
rect 22189 15419 22247 15425
rect 22189 15385 22201 15419
rect 22235 15385 22247 15419
rect 22189 15379 22247 15385
rect 15896 15320 15976 15348
rect 15896 15308 15902 15320
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 16945 15351 17003 15357
rect 16945 15348 16957 15351
rect 16632 15320 16957 15348
rect 16632 15308 16638 15320
rect 16945 15317 16957 15320
rect 16991 15317 17003 15351
rect 16945 15311 17003 15317
rect 17310 15308 17316 15360
rect 17368 15357 17374 15360
rect 17368 15351 17387 15357
rect 17375 15317 17387 15351
rect 17368 15311 17387 15317
rect 17368 15308 17374 15311
rect 20714 15308 20720 15360
rect 20772 15308 20778 15360
rect 22204 15348 22232 15379
rect 22278 15376 22284 15428
rect 22336 15376 22342 15428
rect 22940 15416 22968 15447
rect 23198 15444 23204 15496
rect 23256 15444 23262 15496
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 22388 15388 22968 15416
rect 23400 15416 23428 15447
rect 23474 15444 23480 15496
rect 23532 15444 23538 15496
rect 23566 15444 23572 15496
rect 23624 15444 23630 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 24857 15487 24915 15493
rect 24857 15484 24869 15487
rect 24728 15456 24869 15484
rect 24728 15444 24734 15456
rect 24857 15453 24869 15456
rect 24903 15453 24915 15487
rect 24857 15447 24915 15453
rect 24872 15416 24900 15447
rect 24946 15444 24952 15496
rect 25004 15484 25010 15496
rect 25498 15484 25504 15496
rect 25004 15456 25504 15484
rect 25004 15444 25010 15456
rect 25498 15444 25504 15456
rect 25556 15444 25562 15496
rect 26326 15444 26332 15496
rect 26384 15484 26390 15496
rect 26697 15487 26755 15493
rect 26697 15484 26709 15487
rect 26384 15456 26709 15484
rect 26384 15444 26390 15456
rect 26697 15453 26709 15456
rect 26743 15453 26755 15487
rect 26697 15447 26755 15453
rect 26970 15444 26976 15496
rect 27028 15444 27034 15496
rect 27540 15493 27568 15660
rect 29546 15648 29552 15700
rect 29604 15648 29610 15700
rect 30650 15648 30656 15700
rect 30708 15688 30714 15700
rect 33321 15691 33379 15697
rect 30708 15660 33088 15688
rect 30708 15648 30714 15660
rect 27617 15555 27675 15561
rect 27617 15521 27629 15555
rect 27663 15552 27675 15555
rect 28166 15552 28172 15564
rect 27663 15524 28172 15552
rect 27663 15521 27675 15524
rect 27617 15515 27675 15521
rect 28166 15512 28172 15524
rect 28224 15512 28230 15564
rect 29564 15552 29592 15648
rect 30374 15580 30380 15632
rect 30432 15580 30438 15632
rect 32493 15623 32551 15629
rect 32493 15589 32505 15623
rect 32539 15589 32551 15623
rect 32493 15583 32551 15589
rect 29733 15555 29791 15561
rect 29733 15552 29745 15555
rect 29564 15524 29745 15552
rect 29733 15521 29745 15524
rect 29779 15521 29791 15555
rect 29733 15515 29791 15521
rect 30742 15512 30748 15564
rect 30800 15512 30806 15564
rect 30929 15555 30987 15561
rect 30929 15521 30941 15555
rect 30975 15552 30987 15555
rect 30975 15524 31432 15552
rect 30975 15521 30987 15524
rect 30929 15515 30987 15521
rect 27525 15487 27583 15493
rect 27525 15453 27537 15487
rect 27571 15484 27583 15487
rect 27571 15456 27844 15484
rect 27571 15453 27583 15456
rect 27525 15447 27583 15453
rect 26234 15416 26240 15428
rect 23400 15388 24808 15416
rect 24872 15388 26240 15416
rect 22388 15348 22416 15388
rect 22204 15320 22416 15348
rect 22557 15351 22615 15357
rect 22557 15317 22569 15351
rect 22603 15348 22615 15351
rect 23934 15348 23940 15360
rect 22603 15320 23940 15348
rect 22603 15317 22615 15320
rect 22557 15311 22615 15317
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 24780 15348 24808 15388
rect 26234 15376 26240 15388
rect 26292 15376 26298 15428
rect 27706 15416 27712 15428
rect 26436 15388 27712 15416
rect 26436 15348 26464 15388
rect 27706 15376 27712 15388
rect 27764 15376 27770 15428
rect 27816 15416 27844 15456
rect 27890 15444 27896 15496
rect 27948 15484 27954 15496
rect 28629 15487 28687 15493
rect 28629 15484 28641 15487
rect 27948 15456 28641 15484
rect 27948 15444 27954 15456
rect 28629 15453 28641 15456
rect 28675 15484 28687 15487
rect 29086 15484 29092 15496
rect 28675 15456 29092 15484
rect 28675 15453 28687 15456
rect 28629 15447 28687 15453
rect 29086 15444 29092 15456
rect 29144 15444 29150 15496
rect 29822 15444 29828 15496
rect 29880 15484 29886 15496
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29880 15456 29929 15484
rect 29880 15444 29886 15456
rect 29917 15453 29929 15456
rect 29963 15484 29975 15487
rect 30285 15487 30343 15493
rect 30285 15486 30297 15487
rect 30116 15484 30297 15486
rect 29963 15458 30297 15484
rect 29963 15456 30144 15458
rect 29963 15453 29975 15456
rect 29917 15447 29975 15453
rect 30285 15453 30297 15458
rect 30331 15453 30343 15487
rect 30285 15447 30343 15453
rect 30469 15487 30527 15493
rect 30469 15453 30481 15487
rect 30515 15486 30527 15487
rect 30515 15484 30604 15486
rect 30760 15484 30788 15512
rect 31404 15493 31432 15524
rect 32030 15512 32036 15564
rect 32088 15512 32094 15564
rect 32508 15552 32536 15583
rect 32953 15555 33011 15561
rect 32953 15552 32965 15555
rect 32508 15524 32965 15552
rect 32953 15521 32965 15524
rect 32999 15521 33011 15555
rect 32953 15515 33011 15521
rect 31205 15487 31263 15493
rect 31205 15484 31217 15487
rect 30515 15458 30696 15484
rect 30515 15453 30527 15458
rect 30576 15456 30696 15458
rect 30760 15456 31217 15484
rect 30469 15447 30527 15453
rect 28902 15416 28908 15428
rect 27816 15388 28908 15416
rect 28902 15376 28908 15388
rect 28960 15416 28966 15428
rect 30300 15416 30328 15447
rect 30561 15419 30619 15425
rect 30561 15416 30573 15419
rect 28960 15388 30236 15416
rect 30300 15388 30573 15416
rect 28960 15376 28966 15388
rect 24780 15320 26464 15348
rect 26513 15351 26571 15357
rect 26513 15317 26525 15351
rect 26559 15348 26571 15351
rect 27798 15348 27804 15360
rect 26559 15320 27804 15348
rect 26559 15317 26571 15320
rect 26513 15311 26571 15317
rect 27798 15308 27804 15320
rect 27856 15308 27862 15360
rect 27893 15351 27951 15357
rect 27893 15317 27905 15351
rect 27939 15348 27951 15351
rect 27982 15348 27988 15360
rect 27939 15320 27988 15348
rect 27939 15317 27951 15320
rect 27893 15311 27951 15317
rect 27982 15308 27988 15320
rect 28040 15308 28046 15360
rect 28718 15308 28724 15360
rect 28776 15308 28782 15360
rect 30098 15308 30104 15360
rect 30156 15308 30162 15360
rect 30208 15348 30236 15388
rect 30561 15385 30573 15388
rect 30607 15385 30619 15419
rect 30561 15379 30619 15385
rect 30668 15416 30696 15456
rect 31205 15453 31217 15456
rect 31251 15453 31263 15487
rect 31205 15447 31263 15453
rect 31389 15487 31447 15493
rect 31389 15453 31401 15487
rect 31435 15453 31447 15487
rect 31389 15447 31447 15453
rect 32125 15487 32183 15493
rect 32125 15453 32137 15487
rect 32171 15484 32183 15487
rect 32398 15484 32404 15496
rect 32171 15456 32404 15484
rect 32171 15453 32183 15456
rect 32125 15447 32183 15453
rect 32398 15444 32404 15456
rect 32456 15444 32462 15496
rect 33060 15493 33088 15660
rect 33321 15657 33333 15691
rect 33367 15688 33379 15691
rect 33870 15688 33876 15700
rect 33367 15660 33876 15688
rect 33367 15657 33379 15660
rect 33321 15651 33379 15657
rect 33870 15648 33876 15660
rect 33928 15648 33934 15700
rect 33045 15487 33103 15493
rect 33045 15453 33057 15487
rect 33091 15453 33103 15487
rect 33045 15447 33103 15453
rect 30745 15419 30803 15425
rect 30745 15416 30757 15419
rect 30668 15388 30757 15416
rect 30668 15348 30696 15388
rect 30745 15385 30757 15388
rect 30791 15385 30803 15419
rect 30745 15379 30803 15385
rect 30208 15320 30696 15348
rect 31573 15351 31631 15357
rect 31573 15317 31585 15351
rect 31619 15348 31631 15351
rect 32950 15348 32956 15360
rect 31619 15320 32956 15348
rect 31619 15317 31631 15320
rect 31573 15311 31631 15317
rect 32950 15308 32956 15320
rect 33008 15308 33014 15360
rect 1104 15258 38272 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38272 15258
rect 1104 15184 38272 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1728 15116 1961 15144
rect 1728 15104 1734 15116
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 2593 15147 2651 15153
rect 2593 15113 2605 15147
rect 2639 15113 2651 15147
rect 2593 15107 2651 15113
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2608 15008 2636 15107
rect 2958 15104 2964 15156
rect 3016 15104 3022 15156
rect 3053 15147 3111 15153
rect 3053 15113 3065 15147
rect 3099 15144 3111 15147
rect 3786 15144 3792 15156
rect 3099 15116 3792 15144
rect 3099 15113 3111 15116
rect 3053 15107 3111 15113
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 6822 15144 6828 15156
rect 4755 15116 6828 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7374 15104 7380 15156
rect 7432 15144 7438 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 7432 15116 8125 15144
rect 7432 15104 7438 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8113 15107 8171 15113
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 9493 15147 9551 15153
rect 9493 15144 9505 15147
rect 8812 15116 9505 15144
rect 8812 15104 8818 15116
rect 9493 15113 9505 15116
rect 9539 15113 9551 15147
rect 9493 15107 9551 15113
rect 9950 15104 9956 15156
rect 10008 15104 10014 15156
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 11330 15144 11336 15156
rect 10919 15116 11336 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 6914 15076 6920 15088
rect 6380 15048 6920 15076
rect 6380 15020 6408 15048
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 8294 15076 8300 15088
rect 7866 15048 8300 15076
rect 8294 15036 8300 15048
rect 8352 15076 8358 15088
rect 9306 15076 9312 15088
rect 8352 15048 9312 15076
rect 8352 15036 8358 15048
rect 9306 15036 9312 15048
rect 9364 15036 9370 15088
rect 2179 14980 2636 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 3878 14968 3884 15020
rect 3936 15008 3942 15020
rect 4341 15011 4399 15017
rect 4341 15008 4353 15011
rect 3936 14980 4353 15008
rect 3936 14968 3942 14980
rect 4341 14977 4353 14980
rect 4387 14977 4399 15011
rect 4341 14971 4399 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4706 15008 4712 15020
rect 4571 14980 4712 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 3050 14900 3056 14952
rect 3108 14940 3114 14952
rect 3145 14943 3203 14949
rect 3145 14940 3157 14943
rect 3108 14912 3157 14940
rect 3108 14900 3114 14912
rect 3145 14909 3157 14912
rect 3191 14909 3203 14943
rect 3145 14903 3203 14909
rect 4356 14804 4384 14971
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 6362 14968 6368 15020
rect 6420 14968 6426 15020
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9456 14980 9873 15008
rect 9456 14968 9462 14980
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 11532 15008 11560 15107
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11848 15116 11897 15144
rect 11848 15104 11854 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 11977 15147 12035 15153
rect 11977 15113 11989 15147
rect 12023 15144 12035 15147
rect 12986 15144 12992 15156
rect 12023 15116 12992 15144
rect 12023 15113 12035 15116
rect 11977 15107 12035 15113
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 16114 15144 16120 15156
rect 13403 15116 16120 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 16206 15104 16212 15156
rect 16264 15104 16270 15156
rect 16390 15104 16396 15156
rect 16448 15104 16454 15156
rect 18230 15144 18236 15156
rect 16868 15116 18236 15144
rect 13004 15048 15240 15076
rect 13004 15020 13032 15048
rect 11103 14980 11560 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 12986 14968 12992 15020
rect 13044 14968 13050 15020
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 15008 13231 15011
rect 13262 15008 13268 15020
rect 13219 14980 13268 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13262 14968 13268 14980
rect 13320 15008 13326 15020
rect 13633 15011 13691 15017
rect 13633 15008 13645 15011
rect 13320 14980 13645 15008
rect 13320 14968 13326 14980
rect 13633 14977 13645 14980
rect 13679 15008 13691 15011
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 13679 14980 14565 15008
rect 13679 14977 13691 14980
rect 13633 14971 13691 14977
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 14826 14968 14832 15020
rect 14884 14968 14890 15020
rect 15212 15017 15240 15048
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 16025 15079 16083 15085
rect 16025 15076 16037 15079
rect 15712 15048 16037 15076
rect 15712 15036 15718 15048
rect 16025 15045 16037 15048
rect 16071 15076 16083 15079
rect 16408 15076 16436 15104
rect 16071 15048 16436 15076
rect 16071 15045 16083 15048
rect 16025 15039 16083 15045
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15746 15008 15752 15020
rect 15243 14980 15752 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 6638 14900 6644 14952
rect 6696 14900 6702 14952
rect 10137 14943 10195 14949
rect 10137 14909 10149 14943
rect 10183 14940 10195 14943
rect 11330 14940 11336 14952
rect 10183 14912 11336 14940
rect 10183 14909 10195 14912
rect 10137 14903 10195 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 12066 14900 12072 14952
rect 12124 14900 12130 14952
rect 12526 14900 12532 14952
rect 12584 14940 12590 14952
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 12584 14912 14289 14940
rect 12584 14900 12590 14912
rect 14277 14909 14289 14912
rect 14323 14940 14335 14943
rect 14844 14940 14872 14968
rect 16868 14940 16896 15116
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 20162 15104 20168 15156
rect 20220 15104 20226 15156
rect 20645 15116 21312 15144
rect 17034 15036 17040 15088
rect 17092 15076 17098 15088
rect 17494 15076 17500 15088
rect 17092 15048 17500 15076
rect 17092 15036 17098 15048
rect 17494 15036 17500 15048
rect 17552 15076 17558 15088
rect 19797 15079 19855 15085
rect 17552 15048 18000 15076
rect 17552 15036 17558 15048
rect 16942 14968 16948 15020
rect 17000 15008 17006 15020
rect 17681 15011 17739 15017
rect 17681 15008 17693 15011
rect 17000 14980 17693 15008
rect 17000 14968 17006 14980
rect 17681 14977 17693 14980
rect 17727 15008 17739 15011
rect 17862 15008 17868 15020
rect 17727 14980 17868 15008
rect 17727 14977 17739 14980
rect 17681 14971 17739 14977
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 17972 15017 18000 15048
rect 19797 15045 19809 15079
rect 19843 15076 19855 15079
rect 19978 15076 19984 15088
rect 19843 15048 19984 15076
rect 19843 15045 19855 15048
rect 19797 15039 19855 15045
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 17957 15011 18015 15017
rect 17957 14977 17969 15011
rect 18003 14977 18015 15011
rect 17957 14971 18015 14977
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 18104 14980 18153 15008
rect 18104 14968 18110 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18782 14968 18788 15020
rect 18840 14968 18846 15020
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 14323 14912 14872 14940
rect 15028 14912 16896 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 7650 14832 7656 14884
rect 7708 14872 7714 14884
rect 9858 14872 9864 14884
rect 7708 14844 9864 14872
rect 7708 14832 7714 14844
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 15028 14816 15056 14912
rect 17218 14900 17224 14952
rect 17276 14900 17282 14952
rect 17497 14943 17555 14949
rect 17497 14909 17509 14943
rect 17543 14940 17555 14943
rect 18230 14940 18236 14952
rect 17543 14912 18236 14940
rect 17543 14909 17555 14912
rect 17497 14903 17555 14909
rect 18230 14900 18236 14912
rect 18288 14940 18294 14952
rect 19168 14940 19196 14971
rect 18288 14912 19196 14940
rect 18288 14900 18294 14912
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 15657 14875 15715 14881
rect 15657 14872 15669 14875
rect 15436 14844 15669 14872
rect 15436 14832 15442 14844
rect 15657 14841 15669 14844
rect 15703 14841 15715 14875
rect 15657 14835 15715 14841
rect 16666 14832 16672 14884
rect 16724 14832 16730 14884
rect 17236 14872 17264 14900
rect 17865 14875 17923 14881
rect 17865 14872 17877 14875
rect 17236 14844 17877 14872
rect 17865 14841 17877 14844
rect 17911 14841 17923 14875
rect 20088 14872 20116 14971
rect 20438 14968 20444 15020
rect 20496 15008 20502 15020
rect 20645 15008 20673 15116
rect 20714 15036 20720 15088
rect 20772 15076 20778 15088
rect 20772 15048 21036 15076
rect 20772 15036 20778 15048
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 20496 14980 20821 15008
rect 20496 14968 20502 14980
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 20898 14968 20904 15020
rect 20956 14968 20962 15020
rect 21008 15017 21036 15048
rect 21284 15017 21312 15116
rect 24302 15104 24308 15156
rect 24360 15104 24366 15156
rect 25498 15104 25504 15156
rect 25556 15104 25562 15156
rect 26421 15147 26479 15153
rect 26421 15113 26433 15147
rect 26467 15144 26479 15147
rect 26970 15144 26976 15156
rect 26467 15116 26976 15144
rect 26467 15113 26479 15116
rect 26421 15107 26479 15113
rect 26970 15104 26976 15116
rect 27028 15104 27034 15156
rect 27062 15104 27068 15156
rect 27120 15144 27126 15156
rect 27617 15147 27675 15153
rect 27617 15144 27629 15147
rect 27120 15116 27629 15144
rect 27120 15104 27126 15116
rect 27617 15113 27629 15116
rect 27663 15113 27675 15147
rect 33413 15147 33471 15153
rect 33413 15144 33425 15147
rect 27617 15107 27675 15113
rect 27816 15116 33425 15144
rect 24320 15076 24348 15104
rect 25516 15076 25544 15104
rect 26053 15079 26111 15085
rect 26053 15076 26065 15079
rect 24320 15048 24808 15076
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21192 14940 21220 14971
rect 23382 14968 23388 15020
rect 23440 14968 23446 15020
rect 24578 15008 24584 15020
rect 23492 14980 24584 15008
rect 23492 14952 23520 14980
rect 24578 14968 24584 14980
rect 24636 14968 24642 15020
rect 24780 15017 24808 15048
rect 25516 15048 26065 15076
rect 25516 15017 25544 15048
rect 25792 15017 25820 15048
rect 26053 15045 26065 15048
rect 26099 15045 26111 15079
rect 26053 15039 26111 15045
rect 26234 15036 26240 15088
rect 26292 15036 26298 15088
rect 26510 15036 26516 15088
rect 26568 15076 26574 15088
rect 26605 15079 26663 15085
rect 26605 15076 26617 15079
rect 26568 15048 26617 15076
rect 26568 15036 26574 15048
rect 26605 15045 26617 15048
rect 26651 15045 26663 15079
rect 26605 15039 26663 15045
rect 27816 15017 27844 15116
rect 33413 15113 33425 15116
rect 33459 15113 33471 15147
rect 33413 15107 33471 15113
rect 27982 15036 27988 15088
rect 28040 15076 28046 15088
rect 28350 15076 28356 15088
rect 28040 15048 28356 15076
rect 28040 15036 28046 15048
rect 28350 15036 28356 15048
rect 28408 15076 28414 15088
rect 28997 15079 29055 15085
rect 28408 15048 28488 15076
rect 28408 15036 28414 15048
rect 24765 15011 24823 15017
rect 24765 14977 24777 15011
rect 24811 14977 24823 15011
rect 24765 14971 24823 14977
rect 25501 15011 25559 15017
rect 25501 14977 25513 15011
rect 25547 14977 25559 15011
rect 25501 14971 25559 14977
rect 25685 15011 25743 15017
rect 25685 14977 25697 15011
rect 25731 14977 25743 15011
rect 25685 14971 25743 14977
rect 25777 15011 25835 15017
rect 25777 14977 25789 15011
rect 25823 14977 25835 15011
rect 25777 14971 25835 14977
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 14977 26019 15011
rect 25961 14971 26019 14977
rect 27801 15011 27859 15017
rect 27801 14977 27813 15011
rect 27847 14977 27859 15011
rect 27801 14971 27859 14977
rect 21008 14912 21220 14940
rect 21008 14884 21036 14912
rect 23474 14900 23480 14952
rect 23532 14900 23538 14952
rect 23937 14943 23995 14949
rect 23937 14909 23949 14943
rect 23983 14940 23995 14943
rect 24118 14940 24124 14952
rect 23983 14912 24124 14940
rect 23983 14909 23995 14912
rect 23937 14903 23995 14909
rect 24118 14900 24124 14912
rect 24176 14900 24182 14952
rect 24949 14943 25007 14949
rect 24949 14909 24961 14943
rect 24995 14940 25007 14943
rect 25700 14940 25728 14971
rect 25866 14940 25872 14952
rect 24995 14912 25872 14940
rect 24995 14909 25007 14912
rect 24949 14903 25007 14909
rect 25866 14900 25872 14912
rect 25924 14940 25930 14952
rect 25976 14940 26004 14971
rect 27890 14968 27896 15020
rect 27948 14968 27954 15020
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 15008 28135 15011
rect 28258 15008 28264 15020
rect 28123 14980 28264 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 28460 15019 28488 15048
rect 28552 15048 28948 15076
rect 28445 15013 28503 15019
rect 28445 14979 28457 15013
rect 28491 14979 28503 15013
rect 28445 14973 28503 14979
rect 28552 14949 28580 15048
rect 28813 15011 28871 15017
rect 28813 14977 28825 15011
rect 28859 14977 28871 15011
rect 28920 15008 28948 15048
rect 28997 15045 29009 15079
rect 29043 15076 29055 15079
rect 30650 15076 30656 15088
rect 29043 15048 30656 15076
rect 29043 15045 29055 15048
rect 28997 15039 29055 15045
rect 30650 15036 30656 15048
rect 30708 15036 30714 15088
rect 30852 15048 31340 15076
rect 28920 14980 29040 15008
rect 28813 14971 28871 14977
rect 28537 14943 28595 14949
rect 25924 14912 28120 14940
rect 25924 14900 25930 14912
rect 20162 14872 20168 14884
rect 17865 14835 17923 14841
rect 17972 14844 20168 14872
rect 5442 14804 5448 14816
rect 4356 14776 5448 14804
rect 5442 14764 5448 14776
rect 5500 14804 5506 14816
rect 7282 14804 7288 14816
rect 5500 14776 7288 14804
rect 5500 14764 5506 14776
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 15010 14764 15016 14816
rect 15068 14764 15074 14816
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 15252 14776 16037 14804
rect 15252 14764 15258 14776
rect 16025 14773 16037 14776
rect 16071 14804 16083 14807
rect 16482 14804 16488 14816
rect 16071 14776 16488 14804
rect 16071 14773 16083 14776
rect 16025 14767 16083 14773
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16684 14804 16712 14832
rect 17972 14804 18000 14844
rect 20162 14832 20168 14844
rect 20220 14832 20226 14884
rect 20990 14832 20996 14884
rect 21048 14832 21054 14884
rect 24136 14872 24164 14900
rect 25038 14872 25044 14884
rect 24136 14844 25044 14872
rect 25038 14832 25044 14844
rect 25096 14872 25102 14884
rect 25096 14844 27936 14872
rect 25096 14832 25102 14844
rect 16684 14776 18000 14804
rect 18233 14807 18291 14813
rect 18233 14773 18245 14807
rect 18279 14804 18291 14807
rect 18322 14804 18328 14816
rect 18279 14776 18328 14804
rect 18279 14773 18291 14776
rect 18233 14767 18291 14773
rect 18322 14764 18328 14776
rect 18380 14804 18386 14816
rect 19610 14804 19616 14816
rect 18380 14776 19616 14804
rect 18380 14764 18386 14776
rect 19610 14764 19616 14776
rect 19668 14804 19674 14816
rect 20254 14804 20260 14816
rect 19668 14776 20260 14804
rect 19668 14764 19674 14776
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 20530 14764 20536 14816
rect 20588 14764 20594 14816
rect 21082 14764 21088 14816
rect 21140 14804 21146 14816
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 21140 14776 21373 14804
rect 21140 14764 21146 14776
rect 21361 14773 21373 14776
rect 21407 14773 21419 14807
rect 21361 14767 21419 14773
rect 25590 14764 25596 14816
rect 25648 14764 25654 14816
rect 25774 14764 25780 14816
rect 25832 14764 25838 14816
rect 26694 14764 26700 14816
rect 26752 14764 26758 14816
rect 27908 14804 27936 14844
rect 27982 14832 27988 14884
rect 28040 14832 28046 14884
rect 28092 14872 28120 14912
rect 28537 14909 28549 14943
rect 28583 14909 28595 14943
rect 28537 14903 28595 14909
rect 28626 14900 28632 14952
rect 28684 14900 28690 14952
rect 28828 14872 28856 14971
rect 29012 14940 29040 14980
rect 29086 14968 29092 15020
rect 29144 15008 29150 15020
rect 29181 15011 29239 15017
rect 29181 15008 29193 15011
rect 29144 14980 29193 15008
rect 29144 14968 29150 14980
rect 29181 14977 29193 14980
rect 29227 14977 29239 15011
rect 29181 14971 29239 14977
rect 29362 14968 29368 15020
rect 29420 14968 29426 15020
rect 29564 14980 30144 15008
rect 29564 14952 29592 14980
rect 29012 14912 29316 14940
rect 28092 14844 28856 14872
rect 29288 14872 29316 14912
rect 29546 14900 29552 14952
rect 29604 14900 29610 14952
rect 30006 14900 30012 14952
rect 30064 14900 30070 14952
rect 30024 14872 30052 14900
rect 29288 14844 30052 14872
rect 30116 14872 30144 14980
rect 30558 14968 30564 15020
rect 30616 14968 30622 15020
rect 30852 15017 30880 15048
rect 30837 15011 30895 15017
rect 30837 14977 30849 15011
rect 30883 14977 30895 15011
rect 30837 14971 30895 14977
rect 31021 15011 31079 15017
rect 31021 14977 31033 15011
rect 31067 14977 31079 15011
rect 31312 15008 31340 15048
rect 32858 15036 32864 15088
rect 32916 15036 32922 15088
rect 33042 15036 33048 15088
rect 33100 15036 33106 15088
rect 33245 15079 33303 15085
rect 33245 15076 33257 15079
rect 33152 15048 33257 15076
rect 31754 15008 31760 15020
rect 31312 14980 31760 15008
rect 31021 14971 31079 14977
rect 30193 14943 30251 14949
rect 30193 14909 30205 14943
rect 30239 14940 30251 14943
rect 30576 14940 30604 14968
rect 31036 14940 31064 14971
rect 31754 14968 31760 14980
rect 31812 14968 31818 15020
rect 32876 15008 32904 15036
rect 33152 15008 33180 15048
rect 33245 15045 33257 15048
rect 33291 15076 33303 15079
rect 33781 15079 33839 15085
rect 33781 15076 33793 15079
rect 33291 15048 33793 15076
rect 33291 15045 33303 15048
rect 33245 15039 33303 15045
rect 33781 15045 33793 15048
rect 33827 15045 33839 15079
rect 33781 15039 33839 15045
rect 32876 14980 33180 15008
rect 33410 14968 33416 15020
rect 33468 15008 33474 15020
rect 33505 15011 33563 15017
rect 33505 15008 33517 15011
rect 33468 14980 33517 15008
rect 33468 14968 33474 14980
rect 33505 14977 33517 14980
rect 33551 14977 33563 15011
rect 33505 14971 33563 14977
rect 30239 14912 31064 14940
rect 30239 14909 30251 14912
rect 30193 14903 30251 14909
rect 32950 14900 32956 14952
rect 33008 14940 33014 14952
rect 33781 14943 33839 14949
rect 33781 14940 33793 14943
rect 33008 14912 33793 14940
rect 33008 14900 33014 14912
rect 33781 14909 33793 14912
rect 33827 14909 33839 14943
rect 33781 14903 33839 14909
rect 30282 14872 30288 14884
rect 30116 14844 30288 14872
rect 30282 14832 30288 14844
rect 30340 14872 30346 14884
rect 30340 14844 31754 14872
rect 30340 14832 30346 14844
rect 28626 14804 28632 14816
rect 27908 14776 28632 14804
rect 28626 14764 28632 14776
rect 28684 14764 28690 14816
rect 30837 14807 30895 14813
rect 30837 14773 30849 14807
rect 30883 14804 30895 14807
rect 30926 14804 30932 14816
rect 30883 14776 30932 14804
rect 30883 14773 30895 14776
rect 30837 14767 30895 14773
rect 30926 14764 30932 14776
rect 30984 14764 30990 14816
rect 31726 14804 31754 14844
rect 33226 14804 33232 14816
rect 31726 14776 33232 14804
rect 33226 14764 33232 14776
rect 33284 14764 33290 14816
rect 33594 14764 33600 14816
rect 33652 14764 33658 14816
rect 1104 14714 38272 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38272 14714
rect 1104 14640 38272 14662
rect 6365 14603 6423 14609
rect 6365 14569 6377 14603
rect 6411 14600 6423 14603
rect 6454 14600 6460 14612
rect 6411 14572 6460 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6638 14600 6644 14612
rect 6595 14572 6644 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 13262 14560 13268 14612
rect 13320 14560 13326 14612
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 14366 14600 14372 14612
rect 13964 14572 14372 14600
rect 13964 14560 13970 14572
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 15470 14560 15476 14612
rect 15528 14560 15534 14612
rect 16758 14560 16764 14612
rect 16816 14560 16822 14612
rect 18877 14603 18935 14609
rect 18877 14569 18889 14603
rect 18923 14600 18935 14603
rect 19150 14600 19156 14612
rect 18923 14572 19156 14600
rect 18923 14569 18935 14572
rect 18877 14563 18935 14569
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 19610 14560 19616 14612
rect 19668 14560 19674 14612
rect 20070 14560 20076 14612
rect 20128 14560 20134 14612
rect 22281 14603 22339 14609
rect 22281 14569 22293 14603
rect 22327 14600 22339 14603
rect 23382 14600 23388 14612
rect 22327 14572 23388 14600
rect 22327 14569 22339 14572
rect 22281 14563 22339 14569
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 23477 14603 23535 14609
rect 23477 14569 23489 14603
rect 23523 14600 23535 14603
rect 27246 14600 27252 14612
rect 23523 14572 27252 14600
rect 23523 14569 23535 14572
rect 23477 14563 23535 14569
rect 27246 14560 27252 14572
rect 27304 14560 27310 14612
rect 27341 14603 27399 14609
rect 27341 14569 27353 14603
rect 27387 14600 27399 14603
rect 27982 14600 27988 14612
rect 27387 14572 27988 14600
rect 27387 14569 27399 14572
rect 27341 14563 27399 14569
rect 27982 14560 27988 14572
rect 28040 14560 28046 14612
rect 28166 14560 28172 14612
rect 28224 14560 28230 14612
rect 28350 14560 28356 14612
rect 28408 14560 28414 14612
rect 31941 14603 31999 14609
rect 28966 14572 31800 14600
rect 6472 14532 6500 14560
rect 6822 14532 6828 14544
rect 6472 14504 6828 14532
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 6362 14464 6368 14476
rect 4663 14436 6368 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 6472 14436 7052 14464
rect 3786 14356 3792 14408
rect 3844 14396 3850 14408
rect 3881 14399 3939 14405
rect 3881 14396 3893 14399
rect 3844 14368 3893 14396
rect 3844 14356 3850 14368
rect 3881 14365 3893 14368
rect 3927 14365 3939 14399
rect 3881 14359 3939 14365
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 5994 14356 6000 14408
rect 6052 14396 6058 14408
rect 6472 14396 6500 14436
rect 6052 14368 6500 14396
rect 6733 14399 6791 14405
rect 6052 14356 6058 14368
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 7024 14396 7052 14436
rect 7374 14424 7380 14476
rect 7432 14424 7438 14476
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 8662 14464 8668 14476
rect 7616 14436 8668 14464
rect 7616 14424 7622 14436
rect 8662 14424 8668 14436
rect 8720 14424 8726 14476
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 14292 14436 15117 14464
rect 8294 14396 8300 14408
rect 6779 14368 6960 14396
rect 7024 14368 8300 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 4080 14328 4108 14356
rect 4798 14328 4804 14340
rect 4080 14300 4804 14328
rect 4798 14288 4804 14300
rect 4856 14288 4862 14340
rect 4890 14288 4896 14340
rect 4948 14288 4954 14340
rect 3970 14220 3976 14272
rect 4028 14220 4034 14272
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 6012 14260 6040 14356
rect 6932 14269 6960 14368
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 14292 14405 14320 14436
rect 15105 14433 15117 14436
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14464 15439 14467
rect 15488 14464 15516 14560
rect 15746 14492 15752 14544
rect 15804 14492 15810 14544
rect 20088 14532 20116 14560
rect 17420 14504 20116 14532
rect 16574 14464 16580 14476
rect 15427 14436 15516 14464
rect 16040 14436 16580 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 11112 14368 11529 14396
rect 11112 14356 11118 14368
rect 11517 14365 11529 14368
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14396 14703 14399
rect 14918 14396 14924 14408
rect 14691 14368 14924 14396
rect 14691 14365 14703 14368
rect 14645 14359 14703 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 15010 14356 15016 14408
rect 15068 14356 15074 14408
rect 15286 14356 15292 14408
rect 15344 14356 15350 14408
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 11790 14288 11796 14340
rect 11848 14288 11854 14340
rect 13078 14328 13084 14340
rect 13018 14300 13084 14328
rect 13078 14288 13084 14300
rect 13136 14328 13142 14340
rect 13446 14328 13452 14340
rect 13136 14300 13452 14328
rect 13136 14288 13142 14300
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 15028 14328 15056 14356
rect 15488 14328 15516 14359
rect 15028 14300 15516 14328
rect 4120 14232 6040 14260
rect 6917 14263 6975 14269
rect 4120 14220 4126 14232
rect 6917 14229 6929 14263
rect 6963 14229 6975 14263
rect 6917 14223 6975 14229
rect 7285 14263 7343 14269
rect 7285 14229 7297 14263
rect 7331 14260 7343 14263
rect 10134 14260 10140 14272
rect 7331 14232 10140 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 12434 14260 12440 14272
rect 11756 14232 12440 14260
rect 11756 14220 11762 14232
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 14826 14220 14832 14272
rect 14884 14220 14890 14272
rect 15580 14260 15608 14359
rect 15930 14356 15936 14408
rect 15988 14356 15994 14408
rect 16040 14405 16068 14436
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 17420 14464 17448 14504
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 28368 14532 28396 14560
rect 20772 14504 21220 14532
rect 20772 14492 20778 14504
rect 21192 14476 21220 14504
rect 27816 14504 28396 14532
rect 17144 14436 17448 14464
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14365 16083 14399
rect 16025 14359 16083 14365
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14396 16175 14399
rect 16206 14396 16212 14408
rect 16163 14368 16212 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 16592 14396 16620 14424
rect 16439 14368 16620 14396
rect 16669 14399 16727 14405
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 16669 14365 16681 14399
rect 16715 14396 16727 14399
rect 17144 14396 17172 14436
rect 17494 14424 17500 14476
rect 17552 14424 17558 14476
rect 17678 14424 17684 14476
rect 17736 14464 17742 14476
rect 18782 14464 18788 14476
rect 17736 14436 18788 14464
rect 17736 14424 17742 14436
rect 18782 14424 18788 14436
rect 18840 14424 18846 14476
rect 19058 14424 19064 14476
rect 19116 14464 19122 14476
rect 20898 14464 20904 14476
rect 19116 14436 19656 14464
rect 19116 14424 19122 14436
rect 16715 14368 17172 14396
rect 16715 14365 16727 14368
rect 16669 14359 16727 14365
rect 17218 14356 17224 14408
rect 17276 14396 17282 14408
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17276 14368 17785 14396
rect 17276 14356 17282 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 15838 14288 15844 14340
rect 15896 14328 15902 14340
rect 17788 14328 17816 14359
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 17920 14368 18245 14396
rect 17920 14356 17926 14368
rect 18233 14365 18245 14368
rect 18279 14365 18291 14399
rect 18233 14359 18291 14365
rect 17954 14328 17960 14340
rect 15896 14300 16988 14328
rect 17788 14300 17960 14328
rect 15896 14288 15902 14300
rect 15930 14260 15936 14272
rect 15580 14232 15936 14260
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16114 14220 16120 14272
rect 16172 14260 16178 14272
rect 16960 14269 16988 14300
rect 17954 14288 17960 14300
rect 18012 14288 18018 14340
rect 18506 14288 18512 14340
rect 18564 14288 18570 14340
rect 18800 14337 18828 14424
rect 18601 14331 18659 14337
rect 18601 14297 18613 14331
rect 18647 14297 18659 14331
rect 18601 14291 18659 14297
rect 18785 14331 18843 14337
rect 18785 14297 18797 14331
rect 18831 14297 18843 14331
rect 18785 14291 18843 14297
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 16172 14232 16313 14260
rect 16172 14220 16178 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 16945 14263 17003 14269
rect 16945 14229 16957 14263
rect 16991 14229 17003 14263
rect 16945 14223 17003 14229
rect 18230 14220 18236 14272
rect 18288 14260 18294 14272
rect 18616 14260 18644 14291
rect 19242 14288 19248 14340
rect 19300 14288 19306 14340
rect 19628 14337 19656 14436
rect 19904 14436 20904 14464
rect 19904 14405 19932 14436
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 19622 14331 19680 14337
rect 19622 14297 19634 14331
rect 19668 14328 19680 14331
rect 19996 14328 20024 14359
rect 20162 14356 20168 14408
rect 20220 14356 20226 14408
rect 20438 14356 20444 14408
rect 20496 14356 20502 14408
rect 20732 14405 20760 14436
rect 20898 14424 20904 14436
rect 20956 14424 20962 14476
rect 21174 14424 21180 14476
rect 21232 14424 21238 14476
rect 21821 14467 21879 14473
rect 21821 14433 21833 14467
rect 21867 14464 21879 14467
rect 21867 14436 22140 14464
rect 21867 14433 21879 14436
rect 21821 14427 21879 14433
rect 22112 14405 22140 14436
rect 24946 14424 24952 14476
rect 25004 14464 25010 14476
rect 27816 14464 27844 14504
rect 28966 14464 28994 14572
rect 30650 14532 30656 14544
rect 25004 14436 27660 14464
rect 25004 14424 25010 14436
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14365 20775 14399
rect 20717 14359 20775 14365
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22462 14396 22468 14408
rect 22143 14368 22468 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 19668 14300 20024 14328
rect 20180 14328 20208 14356
rect 21468 14328 21496 14359
rect 20180 14300 21496 14328
rect 22020 14328 22048 14359
rect 22462 14356 22468 14368
rect 22520 14356 22526 14408
rect 23293 14399 23351 14405
rect 23293 14365 23305 14399
rect 23339 14365 23351 14399
rect 23293 14359 23351 14365
rect 22186 14328 22192 14340
rect 22020 14300 22192 14328
rect 19668 14297 19680 14300
rect 19622 14291 19680 14297
rect 22186 14288 22192 14300
rect 22244 14328 22250 14340
rect 23308 14328 23336 14359
rect 24210 14356 24216 14408
rect 24268 14396 24274 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24268 14368 24593 14396
rect 24268 14356 24274 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 24762 14356 24768 14408
rect 24820 14356 24826 14408
rect 25038 14356 25044 14408
rect 25096 14396 25102 14408
rect 27525 14399 27583 14405
rect 27525 14396 27537 14399
rect 25096 14368 27537 14396
rect 25096 14356 25102 14368
rect 27525 14365 27537 14368
rect 27571 14365 27583 14399
rect 27525 14359 27583 14365
rect 22244 14300 23336 14328
rect 24949 14331 25007 14337
rect 22244 14288 22250 14300
rect 24949 14297 24961 14331
rect 24995 14297 25007 14331
rect 27632 14328 27660 14436
rect 27724 14436 27844 14464
rect 28184 14436 28994 14464
rect 30484 14504 30656 14532
rect 27724 14405 27752 14436
rect 27709 14399 27767 14405
rect 27709 14365 27721 14399
rect 27755 14365 27767 14399
rect 27709 14359 27767 14365
rect 27801 14399 27859 14405
rect 27801 14365 27813 14399
rect 27847 14365 27859 14399
rect 27801 14359 27859 14365
rect 27816 14328 27844 14359
rect 28184 14340 28212 14436
rect 28552 14405 28580 14436
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28537 14399 28595 14405
rect 28537 14365 28549 14399
rect 28583 14365 28595 14399
rect 28537 14359 28595 14365
rect 28629 14399 28687 14405
rect 28629 14365 28641 14399
rect 28675 14396 28687 14399
rect 28718 14396 28724 14408
rect 28675 14368 28724 14396
rect 28675 14365 28687 14368
rect 28629 14359 28687 14365
rect 27982 14328 27988 14340
rect 27632 14300 27988 14328
rect 24949 14291 25007 14297
rect 18288 14232 18644 14260
rect 18288 14220 18294 14232
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23474 14260 23480 14272
rect 22796 14232 23480 14260
rect 22796 14220 22802 14232
rect 23474 14220 23480 14232
rect 23532 14220 23538 14272
rect 24964 14260 24992 14291
rect 27982 14288 27988 14300
rect 28040 14288 28046 14340
rect 28166 14288 28172 14340
rect 28224 14288 28230 14340
rect 28368 14328 28396 14359
rect 28718 14356 28724 14368
rect 28776 14356 28782 14408
rect 30484 14405 30512 14504
rect 30650 14492 30656 14504
rect 30708 14532 30714 14544
rect 31113 14535 31171 14541
rect 31113 14532 31125 14535
rect 30708 14504 31125 14532
rect 30708 14492 30714 14504
rect 31113 14501 31125 14504
rect 31159 14501 31171 14535
rect 31113 14495 31171 14501
rect 30561 14467 30619 14473
rect 30561 14433 30573 14467
rect 30607 14464 30619 14467
rect 30607 14436 31248 14464
rect 30607 14433 30619 14436
rect 30561 14427 30619 14433
rect 30469 14399 30527 14405
rect 30469 14365 30481 14399
rect 30515 14365 30527 14399
rect 30469 14359 30527 14365
rect 30653 14399 30711 14405
rect 30653 14365 30665 14399
rect 30699 14396 30711 14399
rect 30834 14396 30840 14408
rect 30699 14368 30840 14396
rect 30699 14365 30711 14368
rect 30653 14359 30711 14365
rect 30834 14356 30840 14368
rect 30892 14356 30898 14408
rect 31220 14405 31248 14436
rect 31205 14399 31263 14405
rect 31205 14365 31217 14399
rect 31251 14365 31263 14399
rect 31389 14399 31447 14405
rect 31389 14396 31401 14399
rect 31205 14359 31263 14365
rect 31312 14368 31401 14396
rect 31312 14340 31340 14368
rect 31389 14365 31401 14368
rect 31435 14365 31447 14399
rect 31389 14359 31447 14365
rect 31478 14356 31484 14408
rect 31536 14356 31542 14408
rect 31570 14356 31576 14408
rect 31628 14396 31634 14408
rect 31772 14405 31800 14572
rect 31941 14569 31953 14603
rect 31987 14600 31999 14603
rect 32030 14600 32036 14612
rect 31987 14572 32036 14600
rect 31987 14569 31999 14572
rect 31941 14563 31999 14569
rect 32030 14560 32036 14572
rect 32088 14560 32094 14612
rect 33042 14560 33048 14612
rect 33100 14560 33106 14612
rect 33318 14560 33324 14612
rect 33376 14560 33382 14612
rect 33060 14532 33088 14560
rect 33505 14535 33563 14541
rect 33505 14532 33517 14535
rect 33060 14504 33517 14532
rect 33505 14501 33517 14504
rect 33551 14501 33563 14535
rect 33505 14495 33563 14501
rect 32950 14424 32956 14476
rect 33008 14464 33014 14476
rect 33229 14467 33287 14473
rect 33229 14464 33241 14467
rect 33008 14436 33241 14464
rect 33008 14424 33014 14436
rect 33229 14433 33241 14436
rect 33275 14433 33287 14467
rect 33229 14427 33287 14433
rect 33594 14424 33600 14476
rect 33652 14424 33658 14476
rect 31757 14399 31815 14405
rect 31628 14368 31708 14396
rect 31628 14356 31634 14368
rect 28368 14300 30696 14328
rect 30466 14260 30472 14272
rect 24964 14232 30472 14260
rect 30466 14220 30472 14232
rect 30524 14220 30530 14272
rect 30668 14260 30696 14300
rect 30742 14288 30748 14340
rect 30800 14288 30806 14340
rect 30926 14288 30932 14340
rect 30984 14288 30990 14340
rect 31294 14288 31300 14340
rect 31352 14288 31358 14340
rect 31680 14328 31708 14368
rect 31757 14365 31769 14399
rect 31803 14365 31815 14399
rect 31757 14359 31815 14365
rect 33137 14399 33195 14405
rect 33137 14365 33149 14399
rect 33183 14396 33195 14399
rect 33612 14396 33640 14424
rect 33183 14368 33640 14396
rect 33183 14365 33195 14368
rect 33137 14359 33195 14365
rect 34054 14356 34060 14408
rect 34112 14356 34118 14408
rect 32674 14328 32680 14340
rect 31680 14300 32680 14328
rect 32674 14288 32680 14300
rect 32732 14328 32738 14340
rect 34072 14328 34100 14356
rect 32732 14300 34100 14328
rect 32732 14288 32738 14300
rect 30944 14260 30972 14288
rect 30668 14232 30972 14260
rect 1104 14170 38272 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38272 14170
rect 1104 14096 38272 14118
rect 3970 14016 3976 14068
rect 4028 14056 4034 14068
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 4028 14028 4077 14056
rect 4028 14016 4034 14028
rect 4065 14025 4077 14028
rect 4111 14025 4123 14059
rect 4065 14019 4123 14025
rect 4614 14016 4620 14068
rect 4672 14065 4678 14068
rect 4672 14059 4691 14065
rect 4679 14025 4691 14059
rect 4672 14019 4691 14025
rect 4672 14016 4678 14019
rect 4798 14016 4804 14068
rect 4856 14016 4862 14068
rect 4890 14016 4896 14068
rect 4948 14056 4954 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 4948 14028 5273 14056
rect 4948 14016 4954 14028
rect 5261 14025 5273 14028
rect 5307 14025 5319 14059
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 5261 14019 5319 14025
rect 5460 14028 6377 14056
rect 3878 13948 3884 14000
rect 3936 13988 3942 14000
rect 4433 13991 4491 13997
rect 4433 13988 4445 13991
rect 3936 13960 4445 13988
rect 3936 13948 3942 13960
rect 4433 13957 4445 13960
rect 4479 13957 4491 13991
rect 4433 13951 4491 13957
rect 2774 13880 2780 13932
rect 2832 13880 2838 13932
rect 5460 13929 5488 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 11146 14056 11152 14068
rect 6365 14019 6423 14025
rect 6656 14028 11152 14056
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13920 4031 13923
rect 5445 13923 5503 13929
rect 4019 13892 5396 13920
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 1394 13812 1400 13864
rect 1452 13812 1458 13864
rect 1670 13812 1676 13864
rect 1728 13812 1734 13864
rect 2792 13852 2820 13880
rect 4062 13852 4068 13864
rect 2792 13824 4068 13852
rect 2884 13728 2912 13824
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 4522 13852 4528 13864
rect 4295 13824 4528 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4522 13812 4528 13824
rect 4580 13852 4586 13864
rect 4798 13852 4804 13864
rect 4580 13824 4804 13852
rect 4580 13812 4586 13824
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5368 13852 5396 13892
rect 5445 13889 5457 13923
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 6656 13852 6684 14028
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11609 14059 11667 14065
rect 11609 14025 11621 14059
rect 11655 14056 11667 14059
rect 11698 14056 11704 14068
rect 11655 14028 11704 14056
rect 11655 14025 11667 14028
rect 11609 14019 11667 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 11848 14028 12449 14056
rect 11848 14016 11854 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 12437 14019 12495 14025
rect 12526 14016 12532 14068
rect 12584 14016 12590 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 14185 14059 14243 14065
rect 14185 14056 14197 14059
rect 13412 14028 14197 14056
rect 13412 14016 13418 14028
rect 14185 14025 14197 14028
rect 14231 14025 14243 14059
rect 14185 14019 14243 14025
rect 14826 14016 14832 14068
rect 14884 14016 14890 14068
rect 14918 14016 14924 14068
rect 14976 14065 14982 14068
rect 14976 14056 14985 14065
rect 14976 14028 15021 14056
rect 14976 14019 14985 14028
rect 14976 14016 14982 14019
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 15344 14028 15485 14056
rect 15344 14016 15350 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 15838 14016 15844 14068
rect 15896 14016 15902 14068
rect 15930 14016 15936 14068
rect 15988 14056 15994 14068
rect 16209 14059 16267 14065
rect 16209 14056 16221 14059
rect 15988 14028 16221 14056
rect 15988 14016 15994 14028
rect 16209 14025 16221 14028
rect 16255 14056 16267 14059
rect 16255 14028 17632 14056
rect 16255 14025 16267 14028
rect 16209 14019 16267 14025
rect 6822 13948 6828 14000
rect 6880 13948 6886 14000
rect 9306 13988 9312 14000
rect 6932 13960 7788 13988
rect 9246 13960 9312 13988
rect 6730 13880 6736 13932
rect 6788 13880 6794 13932
rect 5368 13824 6684 13852
rect 2958 13744 2964 13796
rect 3016 13784 3022 13796
rect 3605 13787 3663 13793
rect 3605 13784 3617 13787
rect 3016 13756 3617 13784
rect 3016 13744 3022 13756
rect 3605 13753 3617 13756
rect 3651 13753 3663 13787
rect 3605 13747 3663 13753
rect 6362 13744 6368 13796
rect 6420 13784 6426 13796
rect 6932 13784 6960 13960
rect 7760 13929 7788 13960
rect 9306 13948 9312 13960
rect 9364 13948 9370 14000
rect 9766 13948 9772 14000
rect 9824 13948 9830 14000
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10134 13988 10140 14000
rect 10008 13960 10140 13988
rect 10008 13948 10014 13960
rect 10134 13948 10140 13960
rect 10192 13988 10198 14000
rect 10229 13991 10287 13997
rect 10229 13988 10241 13991
rect 10192 13960 10241 13988
rect 10192 13948 10198 13960
rect 10229 13957 10241 13960
rect 10275 13957 10287 13991
rect 10229 13951 10287 13957
rect 12069 13991 12127 13997
rect 12069 13957 12081 13991
rect 12115 13988 12127 13991
rect 12544 13988 12572 14016
rect 12115 13960 12572 13988
rect 14093 13991 14151 13997
rect 12115 13957 12127 13960
rect 12069 13951 12127 13957
rect 14093 13957 14105 13991
rect 14139 13988 14151 13991
rect 14844 13988 14872 14016
rect 15856 13988 15884 14016
rect 14139 13960 14872 13988
rect 15120 13960 15884 13988
rect 14139 13957 14151 13960
rect 14093 13951 14151 13957
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13889 7803 13923
rect 9784 13920 9812 13948
rect 10042 13920 10048 13932
rect 9784 13892 10048 13920
rect 7745 13883 7803 13889
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 11882 13920 11888 13932
rect 10888 13892 11888 13920
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 7558 13852 7564 13864
rect 7064 13824 7564 13852
rect 7064 13812 7070 13824
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 9030 13812 9036 13864
rect 9088 13852 9094 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9088 13824 9873 13852
rect 9088 13812 9094 13824
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 10888 13784 10916 13892
rect 11882 13880 11888 13892
rect 11940 13920 11946 13932
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11940 13892 11989 13920
rect 11940 13880 11946 13892
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 12492 13892 12633 13920
rect 12492 13880 12498 13892
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 14829 13923 14887 13929
rect 14829 13920 14841 13923
rect 14792 13892 14841 13920
rect 14792 13880 14798 13892
rect 14829 13889 14841 13892
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 15010 13880 15016 13932
rect 15068 13880 15074 13932
rect 15120 13929 15148 13960
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13889 15163 13923
rect 15105 13883 15163 13889
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13889 15439 13923
rect 15381 13883 15439 13889
rect 11330 13812 11336 13864
rect 11388 13812 11394 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 15396 13852 15424 13883
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 15528 13892 15577 13920
rect 15528 13880 15534 13892
rect 15565 13889 15577 13892
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 16114 13880 16120 13932
rect 16172 13880 16178 13932
rect 16298 13880 16304 13932
rect 16356 13880 16362 13932
rect 17604 13929 17632 14028
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18012 14028 18552 14056
rect 18012 14016 18018 14028
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 17678 13880 17684 13932
rect 17736 13880 17742 13932
rect 17770 13880 17776 13932
rect 17828 13880 17834 13932
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 16574 13852 16580 13864
rect 15396 13824 15608 13852
rect 12161 13815 12219 13821
rect 6420 13756 6960 13784
rect 9048 13756 10916 13784
rect 11348 13784 11376 13812
rect 12176 13784 12204 13815
rect 11348 13756 12204 13784
rect 15580 13784 15608 13824
rect 16500 13824 16580 13852
rect 16500 13784 16528 13824
rect 16574 13812 16580 13824
rect 16632 13812 16638 13864
rect 17221 13855 17279 13861
rect 17221 13821 17233 13855
rect 17267 13852 17279 13855
rect 17696 13852 17724 13880
rect 17267 13824 17724 13852
rect 18248 13852 18276 13883
rect 18322 13880 18328 13932
rect 18380 13880 18386 13932
rect 18524 13929 18552 14028
rect 18782 14016 18788 14068
rect 18840 14056 18846 14068
rect 19242 14056 19248 14068
rect 18840 14028 19248 14056
rect 18840 14016 18846 14028
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 20530 14016 20536 14068
rect 20588 14016 20594 14068
rect 20625 14059 20683 14065
rect 20625 14025 20637 14059
rect 20671 14056 20683 14059
rect 22186 14056 22192 14068
rect 20671 14028 22192 14056
rect 20671 14025 20683 14028
rect 20625 14019 20683 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 23014 14016 23020 14068
rect 23072 14056 23078 14068
rect 23293 14059 23351 14065
rect 23293 14056 23305 14059
rect 23072 14028 23305 14056
rect 23072 14016 23078 14028
rect 23293 14025 23305 14028
rect 23339 14056 23351 14059
rect 24946 14056 24952 14068
rect 23339 14028 24952 14056
rect 23339 14025 23351 14028
rect 23293 14019 23351 14025
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 25038 14016 25044 14068
rect 25096 14016 25102 14068
rect 25314 14016 25320 14068
rect 25372 14016 25378 14068
rect 25866 14016 25872 14068
rect 25924 14016 25930 14068
rect 28258 14016 28264 14068
rect 28316 14056 28322 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 28316 14028 28549 14056
rect 28316 14016 28322 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 28537 14019 28595 14025
rect 28626 14016 28632 14068
rect 28684 14056 28690 14068
rect 28684 14028 28994 14056
rect 28684 14016 28690 14028
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18598 13880 18604 13932
rect 18656 13880 18662 13932
rect 20548 13929 20576 14016
rect 20732 13960 21128 13988
rect 18693 13923 18751 13929
rect 18693 13889 18705 13923
rect 18739 13920 18751 13923
rect 18877 13923 18935 13929
rect 18739 13892 18828 13920
rect 18739 13889 18751 13892
rect 18693 13883 18751 13889
rect 18616 13852 18644 13880
rect 18800 13864 18828 13892
rect 18877 13889 18889 13923
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13889 20591 13923
rect 20533 13883 20591 13889
rect 18248 13824 18644 13852
rect 17267 13821 17279 13824
rect 17221 13815 17279 13821
rect 18782 13812 18788 13864
rect 18840 13812 18846 13864
rect 18892 13852 18920 13883
rect 18966 13852 18972 13864
rect 18892 13824 18972 13852
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 15580 13756 16528 13784
rect 6420 13744 6426 13756
rect 2866 13676 2872 13728
rect 2924 13676 2930 13728
rect 3145 13719 3203 13725
rect 3145 13685 3157 13719
rect 3191 13716 3203 13719
rect 4617 13719 4675 13725
rect 4617 13716 4629 13719
rect 3191 13688 4629 13716
rect 3191 13685 3203 13688
rect 3145 13679 3203 13685
rect 4617 13685 4629 13688
rect 4663 13716 4675 13719
rect 4706 13716 4712 13728
rect 4663 13688 4712 13716
rect 4663 13685 4675 13688
rect 4617 13679 4675 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 8008 13719 8066 13725
rect 8008 13685 8020 13719
rect 8054 13716 8066 13719
rect 8202 13716 8208 13728
rect 8054 13688 8208 13716
rect 8054 13685 8066 13688
rect 8008 13679 8066 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8570 13676 8576 13728
rect 8628 13716 8634 13728
rect 9048 13716 9076 13756
rect 17862 13744 17868 13796
rect 17920 13784 17926 13796
rect 19426 13784 19432 13796
rect 17920 13756 19432 13784
rect 17920 13744 17926 13756
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 8628 13688 9076 13716
rect 8628 13676 8634 13688
rect 9490 13676 9496 13728
rect 9548 13676 9554 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 12066 13716 12072 13728
rect 9640 13688 12072 13716
rect 9640 13676 9646 13688
rect 12066 13676 12072 13688
rect 12124 13676 12130 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 20732 13716 20760 13960
rect 21100 13932 21128 13960
rect 22002 13948 22008 14000
rect 22060 13988 22066 14000
rect 22060 13960 22784 13988
rect 22060 13948 22066 13960
rect 20898 13880 20904 13932
rect 20956 13880 20962 13932
rect 21082 13880 21088 13932
rect 21140 13880 21146 13932
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 22572 13892 22661 13920
rect 20916 13852 20944 13880
rect 22572 13864 22600 13892
rect 22649 13889 22661 13892
rect 22695 13889 22707 13923
rect 22756 13920 22784 13960
rect 22830 13948 22836 14000
rect 22888 13988 22894 14000
rect 25332 13988 25360 14016
rect 22888 13960 25268 13988
rect 25332 13960 25636 13988
rect 22888 13948 22894 13960
rect 23477 13923 23535 13929
rect 23477 13920 23489 13923
rect 22756 13892 23489 13920
rect 22649 13883 22707 13889
rect 23477 13889 23489 13892
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 21361 13855 21419 13861
rect 21361 13852 21373 13855
rect 20916 13824 21373 13852
rect 21361 13821 21373 13824
rect 21407 13821 21419 13855
rect 21361 13815 21419 13821
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 22480 13784 22508 13815
rect 22554 13812 22560 13864
rect 22612 13852 22618 13864
rect 22612 13824 23337 13852
rect 22612 13812 22618 13824
rect 22480 13756 22784 13784
rect 22756 13728 22784 13756
rect 16080 13688 20760 13716
rect 16080 13676 16086 13688
rect 22738 13676 22744 13728
rect 22796 13676 22802 13728
rect 23309 13716 23337 13824
rect 23382 13744 23388 13796
rect 23440 13784 23446 13796
rect 23492 13784 23520 13883
rect 23658 13880 23664 13932
rect 23716 13920 23722 13932
rect 24210 13920 24216 13932
rect 23716 13892 24216 13920
rect 23716 13880 23722 13892
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24765 13923 24823 13929
rect 24765 13889 24777 13923
rect 24811 13918 24823 13923
rect 24854 13918 24860 13932
rect 24811 13890 24860 13918
rect 24811 13889 24823 13890
rect 24765 13883 24823 13889
rect 24854 13880 24860 13890
rect 24912 13880 24918 13932
rect 25130 13880 25136 13932
rect 25188 13880 25194 13932
rect 25240 13929 25268 13960
rect 25225 13923 25283 13929
rect 25225 13889 25237 13923
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 25317 13923 25375 13929
rect 25317 13889 25329 13923
rect 25363 13889 25375 13923
rect 25317 13883 25375 13889
rect 23753 13855 23811 13861
rect 23753 13821 23765 13855
rect 23799 13852 23811 13855
rect 24029 13855 24087 13861
rect 24029 13852 24041 13855
rect 23799 13824 24041 13852
rect 23799 13821 23811 13824
rect 23753 13815 23811 13821
rect 24029 13821 24041 13824
rect 24075 13852 24087 13855
rect 24118 13852 24124 13864
rect 24075 13824 24124 13852
rect 24075 13821 24087 13824
rect 24029 13815 24087 13821
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 24872 13852 24900 13880
rect 24228 13824 24900 13852
rect 25148 13852 25176 13880
rect 25332 13852 25360 13883
rect 25498 13880 25504 13932
rect 25556 13880 25562 13932
rect 25608 13929 25636 13960
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 25682 13880 25688 13932
rect 25740 13880 25746 13932
rect 25884 13929 25912 14016
rect 28966 13988 28994 14028
rect 30742 14016 30748 14068
rect 30800 14056 30806 14068
rect 31205 14059 31263 14065
rect 31205 14056 31217 14059
rect 30800 14028 31217 14056
rect 30800 14016 30806 14028
rect 31205 14025 31217 14028
rect 31251 14025 31263 14059
rect 31205 14019 31263 14025
rect 31570 14016 31576 14068
rect 31628 14016 31634 14068
rect 33318 14016 33324 14068
rect 33376 14056 33382 14068
rect 33597 14059 33655 14065
rect 33597 14056 33609 14059
rect 33376 14028 33609 14056
rect 33376 14016 33382 14028
rect 33597 14025 33609 14028
rect 33643 14056 33655 14059
rect 33643 14028 34008 14056
rect 33643 14025 33655 14028
rect 33597 14019 33655 14025
rect 31588 13988 31616 14016
rect 33870 13988 33876 14000
rect 26252 13960 26924 13988
rect 28966 13960 31616 13988
rect 31864 13960 33876 13988
rect 26252 13929 26280 13960
rect 26896 13932 26924 13960
rect 31864 13932 31892 13960
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13889 25927 13923
rect 25869 13883 25927 13889
rect 26237 13923 26295 13929
rect 26237 13889 26249 13923
rect 26283 13889 26295 13923
rect 26237 13883 26295 13889
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13920 26479 13923
rect 26694 13920 26700 13932
rect 26467 13892 26700 13920
rect 26467 13889 26479 13892
rect 26421 13883 26479 13889
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 26878 13880 26884 13932
rect 26936 13920 26942 13932
rect 26973 13923 27031 13929
rect 26973 13920 26985 13923
rect 26936 13892 26985 13920
rect 26936 13880 26942 13892
rect 26973 13889 26985 13892
rect 27019 13889 27031 13923
rect 26973 13883 27031 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 28166 13920 28172 13932
rect 27203 13892 28172 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 25148 13824 25360 13852
rect 26712 13852 26740 13880
rect 27172 13852 27200 13883
rect 28166 13880 28172 13892
rect 28224 13880 28230 13932
rect 28445 13923 28503 13929
rect 28445 13889 28457 13923
rect 28491 13889 28503 13923
rect 28445 13883 28503 13889
rect 26712 13824 27200 13852
rect 24228 13784 24256 13824
rect 23440 13756 24256 13784
rect 24673 13787 24731 13793
rect 23440 13744 23446 13756
rect 24673 13753 24685 13787
rect 24719 13753 24731 13787
rect 24673 13747 24731 13753
rect 23658 13716 23664 13728
rect 23309 13688 23664 13716
rect 23658 13676 23664 13688
rect 23716 13676 23722 13728
rect 24026 13676 24032 13728
rect 24084 13716 24090 13728
rect 24688 13716 24716 13747
rect 25866 13744 25872 13796
rect 25924 13784 25930 13796
rect 28460 13784 28488 13883
rect 28626 13880 28632 13932
rect 28684 13880 28690 13932
rect 31021 13923 31079 13929
rect 31021 13889 31033 13923
rect 31067 13920 31079 13923
rect 31067 13892 31754 13920
rect 31067 13889 31079 13892
rect 31021 13883 31079 13889
rect 31726 13864 31754 13892
rect 31846 13880 31852 13932
rect 31904 13880 31910 13932
rect 33134 13880 33140 13932
rect 33192 13880 33198 13932
rect 33226 13880 33232 13932
rect 33284 13880 33290 13932
rect 33704 13929 33732 13960
rect 33870 13948 33876 13960
rect 33928 13948 33934 14000
rect 33980 13932 34008 14028
rect 33505 13923 33563 13929
rect 33505 13889 33517 13923
rect 33551 13889 33563 13923
rect 33505 13883 33563 13889
rect 33689 13923 33747 13929
rect 33689 13889 33701 13923
rect 33735 13889 33747 13923
rect 33689 13883 33747 13889
rect 30558 13812 30564 13864
rect 30616 13852 30622 13864
rect 30837 13855 30895 13861
rect 30837 13852 30849 13855
rect 30616 13824 30849 13852
rect 30616 13812 30622 13824
rect 30837 13821 30849 13824
rect 30883 13821 30895 13855
rect 31726 13824 31760 13864
rect 30837 13815 30895 13821
rect 31754 13812 31760 13824
rect 31812 13852 31818 13864
rect 32582 13852 32588 13864
rect 31812 13824 32588 13852
rect 31812 13812 31818 13824
rect 32582 13812 32588 13824
rect 32640 13812 32646 13864
rect 33244 13852 33272 13880
rect 33413 13855 33471 13861
rect 33413 13852 33425 13855
rect 33244 13824 33425 13852
rect 33413 13821 33425 13824
rect 33459 13821 33471 13855
rect 33520 13852 33548 13883
rect 33778 13880 33784 13932
rect 33836 13880 33842 13932
rect 33962 13880 33968 13932
rect 34020 13880 34026 13932
rect 33796 13852 33824 13880
rect 33520 13824 33824 13852
rect 33413 13815 33471 13821
rect 25924 13756 28488 13784
rect 25924 13744 25930 13756
rect 24084 13688 24716 13716
rect 25777 13719 25835 13725
rect 24084 13676 24090 13688
rect 25777 13685 25789 13719
rect 25823 13716 25835 13719
rect 25958 13716 25964 13728
rect 25823 13688 25964 13716
rect 25823 13685 25835 13688
rect 25777 13679 25835 13685
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 26234 13676 26240 13728
rect 26292 13676 26298 13728
rect 27065 13719 27123 13725
rect 27065 13685 27077 13719
rect 27111 13716 27123 13719
rect 27246 13716 27252 13728
rect 27111 13688 27252 13716
rect 27111 13685 27123 13688
rect 27065 13679 27123 13685
rect 27246 13676 27252 13688
rect 27304 13676 27310 13728
rect 28460 13716 28488 13756
rect 28534 13744 28540 13796
rect 28592 13784 28598 13796
rect 29914 13784 29920 13796
rect 28592 13756 29920 13784
rect 28592 13744 28598 13756
rect 29914 13744 29920 13756
rect 29972 13744 29978 13796
rect 33229 13787 33287 13793
rect 33229 13753 33241 13787
rect 33275 13784 33287 13787
rect 33275 13756 33640 13784
rect 33275 13753 33287 13756
rect 33229 13747 33287 13753
rect 33612 13728 33640 13756
rect 31662 13716 31668 13728
rect 28460 13688 31668 13716
rect 31662 13676 31668 13688
rect 31720 13676 31726 13728
rect 32950 13676 32956 13728
rect 33008 13716 33014 13728
rect 33321 13719 33379 13725
rect 33321 13716 33333 13719
rect 33008 13688 33333 13716
rect 33008 13676 33014 13688
rect 33321 13685 33333 13688
rect 33367 13685 33379 13719
rect 33321 13679 33379 13685
rect 33594 13676 33600 13728
rect 33652 13676 33658 13728
rect 1104 13626 38272 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38272 13626
rect 1104 13552 38272 13574
rect 934 13472 940 13524
rect 992 13512 998 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 992 13484 1593 13512
rect 992 13472 998 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1949 13515 2007 13521
rect 1949 13512 1961 13515
rect 1728 13484 1961 13512
rect 1728 13472 1734 13484
rect 1949 13481 1961 13484
rect 1995 13481 2007 13515
rect 1949 13475 2007 13481
rect 3786 13472 3792 13524
rect 3844 13472 3850 13524
rect 6362 13472 6368 13524
rect 6420 13512 6426 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 6420 13484 6561 13512
rect 6420 13472 6426 13484
rect 6549 13481 6561 13484
rect 6595 13512 6607 13515
rect 6822 13512 6828 13524
rect 6595 13484 6828 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 8202 13472 8208 13524
rect 8260 13472 8266 13524
rect 9582 13472 9588 13524
rect 9640 13472 9646 13524
rect 10318 13512 10324 13524
rect 9784 13484 10324 13512
rect 2501 13447 2559 13453
rect 2501 13413 2513 13447
rect 2547 13413 2559 13447
rect 2501 13407 2559 13413
rect 8941 13447 8999 13453
rect 8941 13413 8953 13447
rect 8987 13413 8999 13447
rect 8941 13407 8999 13413
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 2516 13308 2544 13407
rect 2958 13336 2964 13388
rect 3016 13336 3022 13388
rect 3050 13336 3056 13388
rect 3108 13336 3114 13388
rect 3804 13348 4752 13376
rect 3804 13317 3832 13348
rect 4724 13320 4752 13348
rect 2179 13280 2544 13308
rect 2869 13311 2927 13317
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 2915 13280 3801 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 3878 13268 3884 13320
rect 3936 13268 3942 13320
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13308 4123 13311
rect 4111 13280 4660 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 1489 13243 1547 13249
rect 1489 13209 1501 13243
rect 1535 13209 1547 13243
rect 3896 13240 3924 13268
rect 3973 13243 4031 13249
rect 3973 13240 3985 13243
rect 1489 13203 1547 13209
rect 2746 13212 3096 13240
rect 3896 13212 3985 13240
rect 1504 13172 1532 13203
rect 2746 13172 2774 13212
rect 3068 13184 3096 13212
rect 3973 13209 3985 13212
rect 4019 13209 4031 13243
rect 3973 13203 4031 13209
rect 4632 13184 4660 13280
rect 4706 13268 4712 13320
rect 4764 13268 4770 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8956 13308 8984 13407
rect 9600 13385 9628 13472
rect 9784 13385 9812 13484
rect 10318 13472 10324 13484
rect 10376 13472 10382 13524
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 12437 13515 12495 13521
rect 12437 13512 12449 13515
rect 11204 13484 12449 13512
rect 11204 13472 11210 13484
rect 12437 13481 12449 13484
rect 12483 13481 12495 13515
rect 12437 13475 12495 13481
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 14550 13512 14556 13524
rect 12584 13484 14556 13512
rect 12584 13472 12590 13484
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 14921 13515 14979 13521
rect 14921 13481 14933 13515
rect 14967 13512 14979 13515
rect 15010 13512 15016 13524
rect 14967 13484 15016 13512
rect 14967 13481 14979 13484
rect 14921 13475 14979 13481
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 17405 13515 17463 13521
rect 17405 13481 17417 13515
rect 17451 13512 17463 13515
rect 18322 13512 18328 13524
rect 17451 13484 18328 13512
rect 17451 13481 17463 13484
rect 17405 13475 17463 13481
rect 18322 13472 18328 13484
rect 18380 13472 18386 13524
rect 20438 13472 20444 13524
rect 20496 13512 20502 13524
rect 20714 13512 20720 13524
rect 20496 13484 20720 13512
rect 20496 13472 20502 13484
rect 20714 13472 20720 13484
rect 20772 13512 20778 13524
rect 21177 13515 21235 13521
rect 21177 13512 21189 13515
rect 20772 13484 21189 13512
rect 20772 13472 20778 13484
rect 21177 13481 21189 13484
rect 21223 13481 21235 13515
rect 21177 13475 21235 13481
rect 22189 13515 22247 13521
rect 22189 13481 22201 13515
rect 22235 13512 22247 13515
rect 22554 13512 22560 13524
rect 22235 13484 22560 13512
rect 22235 13481 22247 13484
rect 22189 13475 22247 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 23198 13472 23204 13524
rect 23256 13512 23262 13524
rect 24673 13515 24731 13521
rect 23256 13484 23612 13512
rect 23256 13472 23262 13484
rect 15470 13444 15476 13456
rect 12820 13416 13124 13444
rect 12820 13388 12848 13416
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13345 9643 13379
rect 9585 13339 9643 13345
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 9858 13376 9864 13388
rect 9815 13348 9864 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10042 13336 10048 13388
rect 10100 13336 10106 13388
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 10468 13348 12756 13376
rect 10468 13336 10474 13348
rect 8435 13280 8984 13308
rect 9953 13311 10011 13317
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 9953 13277 9965 13311
rect 9999 13308 10011 13311
rect 10060 13308 10088 13336
rect 9999 13280 10088 13308
rect 12728 13308 12756 13348
rect 12802 13336 12808 13388
rect 12860 13336 12866 13388
rect 13096 13385 13124 13416
rect 15120 13416 15476 13444
rect 12897 13379 12955 13385
rect 12897 13345 12909 13379
rect 12943 13376 12955 13379
rect 13081 13379 13139 13385
rect 12943 13348 13032 13376
rect 12943 13345 12955 13348
rect 12897 13339 12955 13345
rect 13004 13308 13032 13348
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13354 13376 13360 13388
rect 13127 13348 13360 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 13170 13308 13176 13320
rect 12728 13280 12940 13308
rect 13004 13280 13176 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 5261 13243 5319 13249
rect 5261 13209 5273 13243
rect 5307 13240 5319 13243
rect 7834 13240 7840 13252
rect 5307 13212 7840 13240
rect 5307 13209 5319 13212
rect 5261 13203 5319 13209
rect 7834 13200 7840 13212
rect 7892 13240 7898 13252
rect 9122 13240 9128 13252
rect 7892 13212 9128 13240
rect 7892 13200 7898 13212
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9401 13243 9459 13249
rect 9401 13209 9413 13243
rect 9447 13240 9459 13243
rect 9490 13240 9496 13252
rect 9447 13212 9496 13240
rect 9447 13209 9459 13212
rect 9401 13203 9459 13209
rect 9490 13200 9496 13212
rect 9548 13240 9554 13252
rect 12526 13240 12532 13252
rect 9548 13212 12532 13240
rect 9548 13200 9554 13212
rect 12526 13200 12532 13212
rect 12584 13200 12590 13252
rect 1504 13144 2774 13172
rect 3050 13132 3056 13184
rect 3108 13132 3114 13184
rect 4614 13132 4620 13184
rect 4672 13132 4678 13184
rect 6730 13132 6736 13184
rect 6788 13172 6794 13184
rect 8662 13172 8668 13184
rect 6788 13144 8668 13172
rect 6788 13132 6794 13144
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 9306 13132 9312 13184
rect 9364 13132 9370 13184
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 10137 13175 10195 13181
rect 10137 13172 10149 13175
rect 9640 13144 10149 13172
rect 9640 13132 9646 13144
rect 10137 13141 10149 13144
rect 10183 13141 10195 13175
rect 10137 13135 10195 13141
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12805 13175 12863 13181
rect 12805 13172 12817 13175
rect 12492 13144 12817 13172
rect 12492 13132 12498 13144
rect 12805 13141 12817 13144
rect 12851 13141 12863 13175
rect 12912 13172 12940 13280
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 15010 13268 15016 13320
rect 15068 13308 15074 13320
rect 15120 13317 15148 13416
rect 15470 13404 15476 13416
rect 15528 13444 15534 13456
rect 16666 13444 16672 13456
rect 15528 13416 16672 13444
rect 15528 13404 15534 13416
rect 16666 13404 16672 13416
rect 16724 13404 16730 13456
rect 22094 13444 22100 13456
rect 18616 13416 22100 13444
rect 15396 13348 15700 13376
rect 15105 13311 15163 13317
rect 15105 13308 15117 13311
rect 15068 13280 15117 13308
rect 15068 13268 15074 13280
rect 15105 13277 15117 13280
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 15396 13317 15424 13348
rect 15672 13320 15700 13348
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 16816 13280 17417 13308
rect 16816 13268 16822 13280
rect 17405 13277 17417 13280
rect 17451 13277 17463 13311
rect 17405 13271 17463 13277
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17552 13280 17601 13308
rect 17552 13268 17558 13280
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 14568 13240 14596 13268
rect 18616 13249 18644 13416
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 23584 13444 23612 13484
rect 24673 13481 24685 13515
rect 24719 13512 24731 13515
rect 25498 13512 25504 13524
rect 24719 13484 25504 13512
rect 24719 13481 24731 13484
rect 24673 13475 24731 13481
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 27246 13472 27252 13524
rect 27304 13512 27310 13524
rect 27304 13484 27660 13512
rect 27304 13472 27310 13484
rect 24854 13444 24860 13456
rect 23584 13416 24860 13444
rect 24854 13404 24860 13416
rect 24912 13404 24918 13456
rect 27632 13444 27660 13484
rect 27890 13472 27896 13524
rect 27948 13512 27954 13524
rect 28261 13515 28319 13521
rect 28261 13512 28273 13515
rect 27948 13484 28273 13512
rect 27948 13472 27954 13484
rect 28261 13481 28273 13484
rect 28307 13481 28319 13515
rect 29181 13515 29239 13521
rect 28261 13475 28319 13481
rect 28368 13484 28994 13512
rect 28368 13444 28396 13484
rect 25792 13416 27568 13444
rect 27632 13416 28396 13444
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 18785 13379 18843 13385
rect 18785 13376 18797 13379
rect 18748 13348 18797 13376
rect 18748 13336 18754 13348
rect 18785 13345 18797 13348
rect 18831 13345 18843 13379
rect 18785 13339 18843 13345
rect 20162 13336 20168 13388
rect 20220 13336 20226 13388
rect 20806 13376 20812 13388
rect 20548 13348 20812 13376
rect 20180 13308 20208 13336
rect 20548 13317 20576 13348
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 23109 13379 23167 13385
rect 21836 13348 22140 13376
rect 20257 13311 20315 13317
rect 20257 13308 20269 13311
rect 20180 13280 20269 13308
rect 20257 13277 20269 13280
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 20533 13311 20591 13317
rect 20533 13277 20545 13311
rect 20579 13277 20591 13311
rect 20533 13271 20591 13277
rect 20626 13311 20684 13317
rect 20626 13277 20638 13311
rect 20672 13308 20684 13311
rect 20714 13308 20720 13320
rect 20672 13280 20720 13308
rect 20672 13277 20684 13280
rect 20626 13271 20684 13277
rect 18601 13243 18659 13249
rect 18601 13240 18613 13243
rect 14568 13212 18613 13240
rect 18601 13209 18613 13212
rect 18647 13209 18659 13243
rect 18601 13203 18659 13209
rect 18693 13243 18751 13249
rect 18693 13209 18705 13243
rect 18739 13240 18751 13243
rect 20346 13240 20352 13252
rect 18739 13212 20352 13240
rect 18739 13209 18751 13212
rect 18693 13203 18751 13209
rect 20346 13200 20352 13212
rect 20404 13200 20410 13252
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 12912 13144 18245 13172
rect 12805 13135 12863 13141
rect 18233 13141 18245 13144
rect 18279 13141 18291 13175
rect 20456 13172 20484 13271
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 21836 13317 21864 13348
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13308 20959 13311
rect 21821 13311 21879 13317
rect 21821 13308 21833 13311
rect 20947 13280 21833 13308
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 21821 13277 21833 13280
rect 21867 13277 21879 13311
rect 21821 13271 21879 13277
rect 22005 13311 22063 13317
rect 22005 13277 22017 13311
rect 22051 13277 22063 13311
rect 22005 13271 22063 13277
rect 20990 13200 20996 13252
rect 21048 13200 21054 13252
rect 21174 13200 21180 13252
rect 21232 13249 21238 13252
rect 21232 13243 21251 13249
rect 21239 13209 21251 13243
rect 22020 13240 22048 13271
rect 21232 13203 21251 13209
rect 21744 13212 22048 13240
rect 22112 13240 22140 13348
rect 22204 13348 22600 13376
rect 22204 13320 22232 13348
rect 22186 13268 22192 13320
rect 22244 13268 22250 13320
rect 22370 13268 22376 13320
rect 22428 13268 22434 13320
rect 22572 13317 22600 13348
rect 23109 13345 23121 13379
rect 23155 13376 23167 13379
rect 25685 13379 25743 13385
rect 25685 13376 25697 13379
rect 23155 13348 25176 13376
rect 23155 13345 23167 13348
rect 23109 13339 23167 13345
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13277 22615 13311
rect 22557 13271 22615 13277
rect 23294 13311 23352 13317
rect 23294 13277 23306 13311
rect 23340 13277 23352 13311
rect 23294 13271 23352 13277
rect 22388 13240 22416 13268
rect 22112 13212 22416 13240
rect 22741 13243 22799 13249
rect 21232 13200 21238 13203
rect 21192 13172 21220 13200
rect 21744 13184 21772 13212
rect 22741 13209 22753 13243
rect 22787 13240 22799 13243
rect 23106 13240 23112 13252
rect 22787 13212 23112 13240
rect 22787 13209 22799 13212
rect 22741 13203 22799 13209
rect 20456 13144 21220 13172
rect 21361 13175 21419 13181
rect 18233 13135 18291 13141
rect 21361 13141 21373 13175
rect 21407 13172 21419 13175
rect 21726 13172 21732 13184
rect 21407 13144 21732 13172
rect 21407 13141 21419 13144
rect 21361 13135 21419 13141
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 21818 13132 21824 13184
rect 21876 13172 21882 13184
rect 22756 13172 22784 13203
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 23308 13240 23336 13271
rect 23382 13268 23388 13320
rect 23440 13268 23446 13320
rect 23474 13268 23480 13320
rect 23532 13268 23538 13320
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13308 23627 13311
rect 23658 13308 23664 13320
rect 23615 13280 23664 13308
rect 23615 13277 23627 13280
rect 23569 13271 23627 13277
rect 23658 13268 23664 13280
rect 23716 13268 23722 13320
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 23750 13240 23756 13252
rect 23308 13212 23756 13240
rect 23750 13200 23756 13212
rect 23808 13200 23814 13252
rect 21876 13144 22784 13172
rect 21876 13132 21882 13144
rect 23382 13132 23388 13184
rect 23440 13172 23446 13184
rect 24872 13172 24900 13271
rect 23440 13144 24900 13172
rect 24964 13172 24992 13271
rect 25038 13268 25044 13320
rect 25096 13268 25102 13320
rect 25148 13317 25176 13348
rect 25240 13348 25697 13376
rect 25240 13317 25268 13348
rect 25685 13345 25697 13348
rect 25731 13345 25743 13379
rect 25685 13339 25743 13345
rect 25792 13320 25820 13416
rect 26160 13348 27476 13376
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13277 25191 13311
rect 25133 13271 25191 13277
rect 25225 13311 25283 13317
rect 25225 13277 25237 13311
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 25593 13311 25651 13317
rect 25593 13277 25605 13311
rect 25639 13277 25651 13311
rect 25593 13271 25651 13277
rect 25056 13240 25084 13268
rect 25608 13240 25636 13271
rect 25774 13268 25780 13320
rect 25832 13268 25838 13320
rect 25958 13268 25964 13320
rect 26016 13308 26022 13320
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 26016 13280 26065 13308
rect 26016 13268 26022 13280
rect 26053 13277 26065 13280
rect 26099 13277 26111 13311
rect 26160 13308 26188 13348
rect 26234 13308 26240 13320
rect 26160 13280 26240 13308
rect 26053 13271 26111 13277
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 26329 13311 26387 13317
rect 26329 13277 26341 13311
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 26344 13240 26372 13271
rect 26418 13268 26424 13320
rect 26476 13268 26482 13320
rect 26510 13268 26516 13320
rect 26568 13308 26574 13320
rect 26605 13311 26663 13317
rect 26605 13308 26617 13311
rect 26568 13280 26617 13308
rect 26568 13268 26574 13280
rect 26605 13277 26617 13280
rect 26651 13277 26663 13311
rect 26970 13308 26976 13320
rect 26605 13271 26663 13277
rect 26712 13280 26976 13308
rect 26712 13240 26740 13280
rect 26970 13268 26976 13280
rect 27028 13268 27034 13320
rect 27065 13311 27123 13317
rect 27065 13277 27077 13311
rect 27111 13277 27123 13311
rect 27065 13271 27123 13277
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13308 27215 13311
rect 27246 13308 27252 13320
rect 27203 13280 27252 13308
rect 27203 13277 27215 13280
rect 27157 13271 27215 13277
rect 25056 13212 26740 13240
rect 26786 13200 26792 13252
rect 26844 13200 26850 13252
rect 25866 13172 25872 13184
rect 24964 13144 25872 13172
rect 23440 13132 23446 13144
rect 25866 13132 25872 13144
rect 25924 13132 25930 13184
rect 26326 13132 26332 13184
rect 26384 13172 26390 13184
rect 26881 13175 26939 13181
rect 26881 13172 26893 13175
rect 26384 13144 26893 13172
rect 26384 13132 26390 13144
rect 26881 13141 26893 13144
rect 26927 13141 26939 13175
rect 27080 13172 27108 13271
rect 27246 13268 27252 13280
rect 27304 13268 27310 13320
rect 27448 13317 27476 13348
rect 27341 13311 27399 13317
rect 27341 13277 27353 13311
rect 27387 13277 27399 13311
rect 27341 13271 27399 13277
rect 27433 13311 27491 13317
rect 27433 13277 27445 13311
rect 27479 13277 27491 13311
rect 27433 13271 27491 13277
rect 27356 13240 27384 13271
rect 27540 13240 27568 13416
rect 28626 13404 28632 13456
rect 28684 13404 28690 13456
rect 28966 13444 28994 13484
rect 29181 13481 29193 13515
rect 29227 13512 29239 13515
rect 29227 13484 29316 13512
rect 29227 13481 29239 13484
rect 29181 13475 29239 13481
rect 29288 13444 29316 13484
rect 30098 13472 30104 13524
rect 30156 13472 30162 13524
rect 31938 13472 31944 13524
rect 31996 13472 32002 13524
rect 32122 13472 32128 13524
rect 32180 13472 32186 13524
rect 33686 13472 33692 13524
rect 33744 13512 33750 13524
rect 33781 13515 33839 13521
rect 33781 13512 33793 13515
rect 33744 13484 33793 13512
rect 33744 13472 33750 13484
rect 33781 13481 33793 13484
rect 33827 13481 33839 13515
rect 33781 13475 33839 13481
rect 29822 13444 29828 13456
rect 28966 13416 29158 13444
rect 29288 13416 29828 13444
rect 28644 13376 28672 13404
rect 29130 13384 29158 13416
rect 29822 13404 29828 13416
rect 29880 13404 29886 13456
rect 29130 13376 29316 13384
rect 29365 13379 29423 13385
rect 29365 13376 29377 13379
rect 28644 13348 28764 13376
rect 29130 13356 29377 13376
rect 29288 13348 29377 13356
rect 28442 13268 28448 13320
rect 28500 13268 28506 13320
rect 28534 13268 28540 13320
rect 28592 13268 28598 13320
rect 28736 13317 28764 13348
rect 29365 13345 29377 13348
rect 29411 13345 29423 13379
rect 30116 13376 30144 13472
rect 32677 13447 32735 13453
rect 32677 13444 32689 13447
rect 31864 13416 32689 13444
rect 31754 13376 31760 13388
rect 30116 13348 31760 13376
rect 29365 13339 29423 13345
rect 28629 13311 28687 13317
rect 28629 13277 28641 13311
rect 28675 13277 28687 13311
rect 28629 13271 28687 13277
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13277 28779 13311
rect 28994 13286 29000 13320
rect 28721 13271 28779 13277
rect 27356 13212 27568 13240
rect 28644 13240 28672 13271
rect 28966 13268 29000 13286
rect 29052 13268 29058 13320
rect 29089 13311 29147 13317
rect 29089 13277 29101 13311
rect 29135 13306 29147 13311
rect 30469 13311 30527 13317
rect 30469 13308 30481 13311
rect 29135 13278 29224 13306
rect 29135 13277 29147 13278
rect 29089 13271 29147 13277
rect 28966 13258 29040 13268
rect 28966 13240 28994 13258
rect 28644 13212 28994 13240
rect 29196 13240 29224 13278
rect 30024 13280 30481 13308
rect 29196 13212 29500 13240
rect 27522 13172 27528 13184
rect 27080 13144 27528 13172
rect 26881 13135 26939 13141
rect 27522 13132 27528 13144
rect 27580 13132 27586 13184
rect 28813 13175 28871 13181
rect 28813 13141 28825 13175
rect 28859 13172 28871 13175
rect 28994 13172 29000 13184
rect 28859 13144 29000 13172
rect 28859 13141 28871 13144
rect 28813 13135 28871 13141
rect 28994 13132 29000 13144
rect 29052 13132 29058 13184
rect 29362 13132 29368 13184
rect 29420 13132 29426 13184
rect 29472 13172 29500 13212
rect 29638 13200 29644 13252
rect 29696 13240 29702 13252
rect 30024 13240 30052 13280
rect 30469 13277 30481 13280
rect 30515 13277 30527 13311
rect 30469 13271 30527 13277
rect 30650 13268 30656 13320
rect 30708 13268 30714 13320
rect 31036 13317 31064 13348
rect 31754 13336 31760 13348
rect 31812 13336 31818 13388
rect 31864 13385 31892 13416
rect 32677 13413 32689 13416
rect 32723 13413 32735 13447
rect 32677 13407 32735 13413
rect 31849 13379 31907 13385
rect 31849 13345 31861 13379
rect 31895 13345 31907 13379
rect 31849 13339 31907 13345
rect 32861 13379 32919 13385
rect 32861 13345 32873 13379
rect 32907 13376 32919 13379
rect 33704 13376 33732 13472
rect 32907 13348 33732 13376
rect 33796 13348 34100 13376
rect 32907 13345 32919 13348
rect 32861 13339 32919 13345
rect 33796 13320 33824 13348
rect 30745 13311 30803 13317
rect 30745 13277 30757 13311
rect 30791 13277 30803 13311
rect 30745 13271 30803 13277
rect 30837 13311 30895 13317
rect 30837 13277 30849 13311
rect 30883 13277 30895 13311
rect 30837 13271 30895 13277
rect 31021 13311 31079 13317
rect 31021 13277 31033 13311
rect 31067 13277 31079 13311
rect 31021 13271 31079 13277
rect 31205 13311 31263 13317
rect 31205 13277 31217 13311
rect 31251 13308 31263 13311
rect 31573 13311 31631 13317
rect 31573 13308 31585 13311
rect 31251 13280 31585 13308
rect 31251 13277 31263 13280
rect 31205 13271 31263 13277
rect 31573 13277 31585 13280
rect 31619 13277 31631 13311
rect 31573 13271 31631 13277
rect 29696 13212 30052 13240
rect 29696 13200 29702 13212
rect 30098 13200 30104 13252
rect 30156 13200 30162 13252
rect 30374 13200 30380 13252
rect 30432 13240 30438 13252
rect 30760 13240 30788 13271
rect 30432 13212 30788 13240
rect 30432 13200 30438 13212
rect 30116 13172 30144 13200
rect 30852 13184 30880 13271
rect 31662 13268 31668 13320
rect 31720 13308 31726 13320
rect 31720 13280 32812 13308
rect 31720 13268 31726 13280
rect 32784 13240 32812 13280
rect 32950 13268 32956 13320
rect 33008 13268 33014 13320
rect 33502 13268 33508 13320
rect 33560 13268 33566 13320
rect 33597 13311 33655 13317
rect 33597 13277 33609 13311
rect 33643 13277 33655 13311
rect 33597 13271 33655 13277
rect 33042 13240 33048 13252
rect 32784 13212 33048 13240
rect 33042 13200 33048 13212
rect 33100 13240 33106 13252
rect 33229 13243 33287 13249
rect 33229 13240 33241 13243
rect 33100 13212 33241 13240
rect 33100 13200 33106 13212
rect 33229 13209 33241 13212
rect 33275 13209 33287 13243
rect 33229 13203 33287 13209
rect 33318 13200 33324 13252
rect 33376 13200 33382 13252
rect 33612 13184 33640 13271
rect 33778 13268 33784 13320
rect 33836 13268 33842 13320
rect 33870 13268 33876 13320
rect 33928 13268 33934 13320
rect 34072 13317 34100 13348
rect 34057 13311 34115 13317
rect 34057 13277 34069 13311
rect 34103 13277 34115 13311
rect 34057 13271 34115 13277
rect 29472 13144 30144 13172
rect 30466 13132 30472 13184
rect 30524 13172 30530 13184
rect 30834 13172 30840 13184
rect 30524 13144 30840 13172
rect 30524 13132 30530 13144
rect 30834 13132 30840 13144
rect 30892 13132 30898 13184
rect 33594 13132 33600 13184
rect 33652 13132 33658 13184
rect 34238 13132 34244 13184
rect 34296 13132 34302 13184
rect 1104 13082 38272 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38272 13082
rect 1104 13008 38272 13030
rect 2866 12968 2872 12980
rect 2746 12940 2872 12968
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 2746 12832 2774 12940
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 4249 12971 4307 12977
rect 4249 12937 4261 12971
rect 4295 12968 4307 12971
rect 6365 12971 6423 12977
rect 4295 12940 5856 12968
rect 4295 12937 4307 12940
rect 4249 12931 4307 12937
rect 4798 12900 4804 12912
rect 4448 12872 4804 12900
rect 2271 12804 2774 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 3878 12832 3884 12844
rect 3476 12804 3884 12832
rect 3476 12792 3482 12804
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 2866 12724 2872 12776
rect 2924 12724 2930 12776
rect 4448 12773 4476 12872
rect 4798 12860 4804 12872
rect 4856 12900 4862 12912
rect 5166 12900 5172 12912
rect 4856 12872 5172 12900
rect 4856 12860 4862 12872
rect 5166 12860 5172 12872
rect 5224 12860 5230 12912
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12733 3571 12767
rect 3513 12727 3571 12733
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 3835 12736 4353 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 4433 12767 4491 12773
rect 4433 12733 4445 12767
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 3528 12696 3556 12727
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 4632 12696 4660 12724
rect 3528 12668 4660 12696
rect 5828 12696 5856 12940
rect 6365 12937 6377 12971
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12832 5963 12835
rect 6380 12832 6408 12931
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6604 12940 6837 12968
rect 6604 12928 6610 12940
rect 6825 12937 6837 12940
rect 6871 12968 6883 12971
rect 7190 12968 7196 12980
rect 6871 12940 7196 12968
rect 6871 12937 6883 12940
rect 6825 12931 6883 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 9272 12940 9321 12968
rect 9272 12928 9278 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 10597 12971 10655 12977
rect 10597 12937 10609 12971
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 8754 12860 8760 12912
rect 8812 12860 8818 12912
rect 5951 12804 6408 12832
rect 6733 12835 6791 12841
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 6733 12801 6745 12835
rect 6779 12832 6791 12835
rect 8202 12832 8208 12844
rect 6779 12804 8208 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 10410 12832 10416 12844
rect 8312 12804 10416 12832
rect 7006 12724 7012 12776
rect 7064 12724 7070 12776
rect 8312 12696 8340 12804
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10612 12832 10640 12931
rect 10870 12928 10876 12980
rect 10928 12928 10934 12980
rect 11057 12971 11115 12977
rect 11057 12937 11069 12971
rect 11103 12968 11115 12971
rect 11974 12968 11980 12980
rect 11103 12940 11980 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 11974 12928 11980 12940
rect 12032 12968 12038 12980
rect 12250 12968 12256 12980
rect 12032 12940 12256 12968
rect 12032 12928 12038 12940
rect 12250 12928 12256 12940
rect 12308 12968 12314 12980
rect 15010 12968 15016 12980
rect 12308 12940 15016 12968
rect 12308 12928 12314 12940
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 16172 12940 16221 12968
rect 16172 12928 16178 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 16209 12931 16267 12937
rect 18138 12928 18144 12980
rect 18196 12928 18202 12980
rect 20441 12971 20499 12977
rect 20441 12937 20453 12971
rect 20487 12968 20499 12971
rect 20487 12940 22094 12968
rect 20487 12937 20499 12940
rect 20441 12931 20499 12937
rect 10551 12804 10640 12832
rect 10888 12832 10916 12928
rect 14090 12900 14096 12912
rect 11072 12872 14096 12900
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10888 12804 10977 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8720 12736 9229 12764
rect 8720 12724 8726 12736
rect 9217 12733 9229 12736
rect 9263 12764 9275 12767
rect 9306 12764 9312 12776
rect 9263 12736 9312 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 9306 12724 9312 12736
rect 9364 12764 9370 12776
rect 9582 12764 9588 12776
rect 9364 12736 9588 12764
rect 9364 12724 9370 12736
rect 9582 12724 9588 12736
rect 9640 12764 9646 12776
rect 11072 12764 11100 12872
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 16022 12860 16028 12912
rect 16080 12860 16086 12912
rect 11330 12832 11336 12844
rect 11256 12804 11336 12832
rect 11256 12773 11284 12804
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12400 12804 13185 12832
rect 12400 12792 12406 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 14918 12832 14924 12844
rect 13311 12804 14924 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 14918 12792 14924 12804
rect 14976 12832 14982 12844
rect 16850 12832 16856 12844
rect 14976 12804 16856 12832
rect 14976 12792 14982 12804
rect 16850 12792 16856 12804
rect 16908 12832 16914 12844
rect 17494 12832 17500 12844
rect 16908 12804 17500 12832
rect 16908 12792 16914 12804
rect 17494 12792 17500 12804
rect 17552 12832 17558 12844
rect 18156 12832 18184 12928
rect 18598 12860 18604 12912
rect 18656 12900 18662 12912
rect 20901 12903 20959 12909
rect 18656 12872 18814 12900
rect 18656 12860 18662 12872
rect 20901 12869 20913 12903
rect 20947 12900 20959 12903
rect 20990 12900 20996 12912
rect 20947 12872 20996 12900
rect 20947 12869 20959 12872
rect 20901 12863 20959 12869
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 17552 12804 17908 12832
rect 18156 12804 18245 12832
rect 17552 12792 17558 12804
rect 9640 12736 11100 12764
rect 11241 12767 11299 12773
rect 9640 12724 9646 12736
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 11287 12736 13369 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 13357 12733 13369 12736
rect 13403 12764 13415 12767
rect 13630 12764 13636 12776
rect 13403 12736 13636 12764
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 13630 12724 13636 12736
rect 13688 12764 13694 12776
rect 15378 12764 15384 12776
rect 13688 12736 15384 12764
rect 13688 12724 13694 12736
rect 15378 12724 15384 12736
rect 15436 12764 15442 12776
rect 15562 12764 15568 12776
rect 15436 12736 15568 12764
rect 15436 12724 15442 12736
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 17770 12764 17776 12776
rect 15672 12736 17776 12764
rect 5828 12668 8340 12696
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12696 8815 12699
rect 9030 12696 9036 12708
rect 8803 12668 9036 12696
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 12250 12656 12256 12708
rect 12308 12696 12314 12708
rect 12308 12668 12940 12696
rect 12308 12656 12314 12668
rect 3878 12588 3884 12640
rect 3936 12588 3942 12640
rect 5718 12588 5724 12640
rect 5776 12588 5782 12640
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 8444 12600 9505 12628
rect 8444 12588 8450 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9493 12591 9551 12597
rect 10321 12631 10379 12637
rect 10321 12597 10333 12631
rect 10367 12628 10379 12631
rect 10410 12628 10416 12640
rect 10367 12600 10416 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 12802 12588 12808 12640
rect 12860 12588 12866 12640
rect 12912 12628 12940 12668
rect 15672 12628 15700 12736
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 17880 12696 17908 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 18380 12804 18429 12832
rect 18380 12792 18386 12804
rect 18417 12801 18429 12804
rect 18463 12832 18475 12835
rect 19058 12832 19064 12844
rect 18463 12804 19064 12832
rect 18463 12801 18475 12804
rect 18417 12795 18475 12801
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12832 20315 12835
rect 20806 12832 20812 12844
rect 20303 12804 20812 12832
rect 20303 12801 20315 12804
rect 20257 12795 20315 12801
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 20625 12767 20683 12773
rect 20625 12733 20637 12767
rect 20671 12764 20683 12767
rect 20916 12764 20944 12863
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 21101 12903 21159 12909
rect 21101 12900 21113 12903
rect 21100 12869 21113 12900
rect 21147 12869 21159 12903
rect 22066 12900 22094 12940
rect 23014 12928 23020 12980
rect 23072 12968 23078 12980
rect 23382 12968 23388 12980
rect 23072 12940 23388 12968
rect 23072 12928 23078 12940
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 25130 12928 25136 12980
rect 25188 12968 25194 12980
rect 25590 12968 25596 12980
rect 25188 12940 25596 12968
rect 25188 12928 25194 12940
rect 25590 12928 25596 12940
rect 25648 12968 25654 12980
rect 25648 12940 26556 12968
rect 25648 12928 25654 12940
rect 23569 12903 23627 12909
rect 23569 12900 23581 12903
rect 22066 12872 23581 12900
rect 21100 12863 21159 12869
rect 20671 12736 20944 12764
rect 20671 12733 20683 12736
rect 20625 12727 20683 12733
rect 20640 12696 20668 12727
rect 15804 12668 16436 12696
rect 17880 12668 20668 12696
rect 15804 12656 15810 12668
rect 16408 12637 16436 12668
rect 20898 12656 20904 12708
rect 20956 12696 20962 12708
rect 21100 12696 21128 12863
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 22848 12841 22876 12872
rect 23308 12841 23336 12872
rect 23569 12869 23581 12872
rect 23615 12869 23627 12903
rect 24578 12900 24584 12912
rect 23569 12863 23627 12869
rect 23860 12872 24584 12900
rect 22649 12835 22707 12841
rect 22649 12832 22661 12835
rect 22520 12804 22661 12832
rect 22520 12792 22526 12804
rect 22649 12801 22661 12804
rect 22695 12801 22707 12835
rect 22649 12795 22707 12801
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12801 22891 12835
rect 22833 12795 22891 12801
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 23753 12835 23811 12841
rect 23753 12801 23765 12835
rect 23799 12801 23811 12835
rect 23753 12795 23811 12801
rect 21726 12724 21732 12776
rect 21784 12764 21790 12776
rect 21821 12767 21879 12773
rect 21821 12764 21833 12767
rect 21784 12736 21833 12764
rect 21784 12724 21790 12736
rect 21821 12733 21833 12736
rect 21867 12733 21879 12767
rect 21821 12727 21879 12733
rect 22094 12724 22100 12776
rect 22152 12724 22158 12776
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 22370 12724 22376 12776
rect 22428 12764 22434 12776
rect 23216 12764 23244 12795
rect 23768 12764 23796 12795
rect 22428 12736 23796 12764
rect 22428 12724 22434 12736
rect 20956 12668 21128 12696
rect 22296 12696 22324 12724
rect 22738 12696 22744 12708
rect 22296 12668 22744 12696
rect 20956 12656 20962 12668
rect 22738 12656 22744 12668
rect 22796 12656 22802 12708
rect 22925 12699 22983 12705
rect 22925 12665 22937 12699
rect 22971 12696 22983 12699
rect 23750 12696 23756 12708
rect 22971 12668 23756 12696
rect 22971 12665 22983 12668
rect 22925 12659 22983 12665
rect 23750 12656 23756 12668
rect 23808 12696 23814 12708
rect 23860 12696 23888 12872
rect 24578 12860 24584 12872
rect 24636 12900 24642 12912
rect 25682 12900 25688 12912
rect 24636 12872 25688 12900
rect 24636 12860 24642 12872
rect 25682 12860 25688 12872
rect 25740 12860 25746 12912
rect 24394 12792 24400 12844
rect 24452 12832 24458 12844
rect 25314 12832 25320 12844
rect 24452 12804 25320 12832
rect 24452 12792 24458 12804
rect 25314 12792 25320 12804
rect 25372 12792 25378 12844
rect 26326 12792 26332 12844
rect 26384 12792 26390 12844
rect 26528 12841 26556 12940
rect 26786 12928 26792 12980
rect 26844 12928 26850 12980
rect 28626 12928 28632 12980
rect 28684 12968 28690 12980
rect 29181 12971 29239 12977
rect 28684 12940 29040 12968
rect 28684 12928 28690 12940
rect 26804 12900 26832 12928
rect 26804 12872 27476 12900
rect 26513 12835 26571 12841
rect 26513 12801 26525 12835
rect 26559 12801 26571 12835
rect 26513 12795 26571 12801
rect 26602 12792 26608 12844
rect 26660 12832 26666 12844
rect 26970 12832 26976 12844
rect 26660 12804 26976 12832
rect 26660 12792 26666 12804
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27246 12792 27252 12844
rect 27304 12792 27310 12844
rect 27448 12841 27476 12872
rect 28902 12860 28908 12912
rect 28960 12860 28966 12912
rect 29012 12900 29040 12940
rect 29181 12937 29193 12971
rect 29227 12937 29239 12971
rect 29181 12931 29239 12937
rect 31113 12971 31171 12977
rect 31113 12937 31125 12971
rect 31159 12968 31171 12971
rect 31478 12968 31484 12980
rect 31159 12940 31484 12968
rect 31159 12937 31171 12940
rect 31113 12931 31171 12937
rect 29196 12900 29224 12931
rect 31478 12928 31484 12940
rect 31536 12928 31542 12980
rect 32493 12971 32551 12977
rect 32493 12968 32505 12971
rect 31804 12940 32505 12968
rect 31804 12909 31832 12940
rect 32493 12937 32505 12940
rect 32539 12937 32551 12971
rect 32493 12931 32551 12937
rect 33042 12928 33048 12980
rect 33100 12928 33106 12980
rect 33134 12928 33140 12980
rect 33192 12968 33198 12980
rect 33502 12968 33508 12980
rect 33192 12940 33508 12968
rect 33192 12928 33198 12940
rect 33502 12928 33508 12940
rect 33560 12968 33566 12980
rect 33873 12971 33931 12977
rect 33873 12968 33885 12971
rect 33560 12940 33885 12968
rect 33560 12928 33566 12940
rect 33873 12937 33885 12940
rect 33919 12937 33931 12971
rect 33873 12931 33931 12937
rect 34238 12928 34244 12980
rect 34296 12928 34302 12980
rect 31389 12903 31447 12909
rect 31389 12900 31401 12903
rect 29012 12872 29592 12900
rect 27341 12835 27399 12841
rect 27341 12801 27353 12835
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12801 27491 12835
rect 27433 12795 27491 12801
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 25038 12764 25044 12776
rect 24912 12736 25044 12764
rect 24912 12724 24918 12736
rect 25038 12724 25044 12736
rect 25096 12724 25102 12776
rect 23808 12668 23888 12696
rect 23808 12656 23814 12668
rect 26326 12656 26332 12708
rect 26384 12696 26390 12708
rect 26421 12699 26479 12705
rect 26421 12696 26433 12699
rect 26384 12668 26433 12696
rect 26384 12656 26390 12668
rect 26421 12665 26433 12668
rect 26467 12665 26479 12699
rect 27356 12696 27384 12795
rect 27614 12792 27620 12844
rect 27672 12792 27678 12844
rect 28813 12835 28871 12841
rect 28813 12801 28825 12835
rect 28859 12832 28871 12835
rect 28920 12832 28948 12860
rect 28859 12804 28948 12832
rect 28859 12801 28871 12804
rect 28813 12795 28871 12801
rect 29086 12792 29092 12844
rect 29144 12792 29150 12844
rect 29270 12792 29276 12844
rect 29328 12792 29334 12844
rect 29457 12835 29515 12841
rect 29457 12801 29469 12835
rect 29503 12832 29515 12835
rect 29564 12832 29592 12872
rect 29503 12804 29592 12832
rect 30300 12872 31401 12900
rect 29503 12801 29515 12804
rect 29457 12795 29515 12801
rect 28905 12767 28963 12773
rect 28905 12733 28917 12767
rect 28951 12764 28963 12767
rect 28994 12764 29000 12776
rect 28951 12736 29000 12764
rect 28951 12733 28963 12736
rect 28905 12727 28963 12733
rect 28994 12724 29000 12736
rect 29052 12724 29058 12776
rect 26421 12659 26479 12665
rect 26896 12668 27384 12696
rect 29104 12696 29132 12792
rect 29288 12764 29316 12792
rect 30300 12764 30328 12872
rect 31389 12869 31401 12872
rect 31435 12900 31447 12903
rect 31573 12903 31631 12909
rect 31573 12900 31585 12903
rect 31435 12872 31585 12900
rect 31435 12869 31447 12872
rect 31389 12863 31447 12869
rect 31573 12869 31585 12872
rect 31619 12869 31631 12903
rect 31573 12863 31631 12869
rect 31789 12903 31847 12909
rect 31789 12869 31801 12903
rect 31835 12869 31847 12903
rect 32309 12903 32367 12909
rect 32309 12900 32321 12903
rect 31789 12863 31847 12869
rect 31956 12872 32321 12900
rect 30558 12792 30564 12844
rect 30616 12832 30622 12844
rect 30745 12835 30803 12841
rect 30745 12832 30757 12835
rect 30616 12804 30757 12832
rect 30616 12792 30622 12804
rect 30745 12801 30757 12804
rect 30791 12801 30803 12835
rect 30745 12795 30803 12801
rect 31297 12835 31355 12841
rect 31297 12801 31309 12835
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 30653 12767 30711 12773
rect 30653 12764 30665 12767
rect 29288 12736 30328 12764
rect 30392 12736 30665 12764
rect 29273 12699 29331 12705
rect 29273 12696 29285 12699
rect 29104 12668 29285 12696
rect 16209 12631 16267 12637
rect 16209 12628 16221 12631
rect 12912 12600 16221 12628
rect 16209 12597 16221 12600
rect 16255 12597 16267 12631
rect 16209 12591 16267 12597
rect 16393 12631 16451 12637
rect 16393 12597 16405 12631
rect 16439 12597 16451 12631
rect 16393 12591 16451 12597
rect 20714 12588 20720 12640
rect 20772 12588 20778 12640
rect 21082 12588 21088 12640
rect 21140 12588 21146 12640
rect 21269 12631 21327 12637
rect 21269 12597 21281 12631
rect 21315 12628 21327 12631
rect 22646 12628 22652 12640
rect 21315 12600 22652 12628
rect 21315 12597 21327 12600
rect 21269 12591 21327 12597
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 23845 12631 23903 12637
rect 23845 12597 23857 12631
rect 23891 12628 23903 12631
rect 24486 12628 24492 12640
rect 23891 12600 24492 12628
rect 23891 12597 23903 12600
rect 23845 12591 23903 12597
rect 24486 12588 24492 12600
rect 24544 12588 24550 12640
rect 25682 12588 25688 12640
rect 25740 12628 25746 12640
rect 26602 12628 26608 12640
rect 25740 12600 26608 12628
rect 25740 12588 25746 12600
rect 26602 12588 26608 12600
rect 26660 12628 26666 12640
rect 26896 12628 26924 12668
rect 29273 12665 29285 12668
rect 29319 12665 29331 12699
rect 29638 12696 29644 12708
rect 29273 12659 29331 12665
rect 29380 12668 29644 12696
rect 26660 12600 26924 12628
rect 26973 12631 27031 12637
rect 26660 12588 26666 12600
rect 26973 12597 26985 12631
rect 27019 12628 27031 12631
rect 29380 12628 29408 12668
rect 29638 12656 29644 12668
rect 29696 12656 29702 12708
rect 29822 12656 29828 12708
rect 29880 12696 29886 12708
rect 30392 12696 30420 12736
rect 30653 12733 30665 12736
rect 30699 12733 30711 12767
rect 31312 12764 31340 12795
rect 31478 12792 31484 12844
rect 31536 12832 31542 12844
rect 31956 12832 31984 12872
rect 32309 12869 32321 12872
rect 32355 12900 32367 12903
rect 33318 12900 33324 12912
rect 32355 12872 33324 12900
rect 32355 12869 32367 12872
rect 32309 12863 32367 12869
rect 33318 12860 33324 12872
rect 33376 12860 33382 12912
rect 34256 12900 34284 12928
rect 33796 12872 34284 12900
rect 31536 12804 31984 12832
rect 32125 12835 32183 12841
rect 31536 12792 31542 12804
rect 32125 12801 32137 12835
rect 32171 12830 32183 12835
rect 32171 12802 32260 12830
rect 32171 12801 32183 12802
rect 32125 12795 32183 12801
rect 31754 12764 31760 12776
rect 31312 12736 31760 12764
rect 30653 12727 30711 12733
rect 31754 12724 31760 12736
rect 31812 12764 31818 12776
rect 32232 12764 32260 12802
rect 32950 12792 32956 12844
rect 33008 12792 33014 12844
rect 33796 12841 33824 12872
rect 33413 12835 33471 12841
rect 33413 12801 33425 12835
rect 33459 12801 33471 12835
rect 33413 12795 33471 12801
rect 33781 12835 33839 12841
rect 33781 12801 33793 12835
rect 33827 12801 33839 12835
rect 33781 12795 33839 12801
rect 31812 12736 32260 12764
rect 31812 12724 31818 12736
rect 32490 12724 32496 12776
rect 32548 12764 32554 12776
rect 33428 12764 33456 12795
rect 33962 12792 33968 12844
rect 34020 12792 34026 12844
rect 32548 12736 33456 12764
rect 32548 12724 32554 12736
rect 29880 12668 30420 12696
rect 29880 12656 29886 12668
rect 30466 12656 30472 12708
rect 30524 12696 30530 12708
rect 30524 12668 31156 12696
rect 30524 12656 30530 12668
rect 27019 12600 29408 12628
rect 27019 12597 27031 12600
rect 26973 12591 27031 12597
rect 29546 12588 29552 12640
rect 29604 12628 29610 12640
rect 30374 12628 30380 12640
rect 29604 12600 30380 12628
rect 29604 12588 29610 12600
rect 30374 12588 30380 12600
rect 30432 12588 30438 12640
rect 31128 12628 31156 12668
rect 31938 12656 31944 12708
rect 31996 12656 32002 12708
rect 33428 12696 33456 12736
rect 34330 12696 34336 12708
rect 33428 12668 34336 12696
rect 34330 12656 34336 12668
rect 34388 12656 34394 12708
rect 31757 12631 31815 12637
rect 31757 12628 31769 12631
rect 31128 12600 31769 12628
rect 31757 12597 31769 12600
rect 31803 12597 31815 12631
rect 31757 12591 31815 12597
rect 1104 12538 38272 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38272 12538
rect 1104 12464 38272 12486
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 8846 12424 8852 12436
rect 8619 12396 8852 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 15102 12424 15108 12436
rect 11664 12396 15108 12424
rect 11664 12384 11670 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 19392 12396 19441 12424
rect 19392 12384 19398 12396
rect 19429 12393 19441 12396
rect 19475 12393 19487 12427
rect 19889 12427 19947 12433
rect 19889 12424 19901 12427
rect 19429 12387 19487 12393
rect 19536 12396 19901 12424
rect 1394 12316 1400 12368
rect 1452 12356 1458 12368
rect 1452 12328 5212 12356
rect 1452 12316 1458 12328
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3234 12288 3240 12300
rect 2915 12260 3240 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3234 12248 3240 12260
rect 3292 12288 3298 12300
rect 3786 12288 3792 12300
rect 3292 12260 3792 12288
rect 3292 12248 3298 12260
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 5184 12297 5212 12328
rect 8018 12316 8024 12368
rect 8076 12356 8082 12368
rect 8941 12359 8999 12365
rect 8941 12356 8953 12359
rect 8076 12328 8953 12356
rect 8076 12316 8082 12328
rect 8941 12325 8953 12328
rect 8987 12325 8999 12359
rect 8941 12319 8999 12325
rect 9309 12359 9367 12365
rect 9309 12325 9321 12359
rect 9355 12356 9367 12359
rect 9398 12356 9404 12368
rect 9355 12328 9404 12356
rect 9355 12325 9367 12328
rect 9309 12319 9367 12325
rect 9398 12316 9404 12328
rect 9456 12316 9462 12368
rect 15396 12328 16068 12356
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12288 5227 12291
rect 6086 12288 6092 12300
rect 5215 12260 6092 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 6880 12260 10241 12288
rect 6880 12248 6886 12260
rect 10229 12257 10241 12260
rect 10275 12288 10287 12291
rect 11054 12288 11060 12300
rect 10275 12260 11060 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12253 12291 12311 12297
rect 12253 12288 12265 12291
rect 12032 12260 12265 12288
rect 12032 12248 12038 12260
rect 12253 12257 12265 12260
rect 12299 12257 12311 12291
rect 13262 12288 13268 12300
rect 12253 12251 12311 12257
rect 12728 12260 13268 12288
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12220 2007 12223
rect 2685 12223 2743 12229
rect 1995 12192 2268 12220
rect 1995 12189 2007 12192
rect 1949 12183 2007 12189
rect 1762 12044 1768 12096
rect 1820 12044 1826 12096
rect 2240 12093 2268 12192
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 3878 12220 3884 12232
rect 2731 12192 3884 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 8343 12192 8708 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 2593 12155 2651 12161
rect 2593 12121 2605 12155
rect 2639 12152 2651 12155
rect 2774 12152 2780 12164
rect 2639 12124 2780 12152
rect 2639 12121 2651 12124
rect 2593 12115 2651 12121
rect 2774 12112 2780 12124
rect 2832 12152 2838 12164
rect 3418 12152 3424 12164
rect 2832 12124 3424 12152
rect 2832 12112 2838 12124
rect 3418 12112 3424 12124
rect 3476 12112 3482 12164
rect 5445 12155 5503 12161
rect 5445 12121 5457 12155
rect 5491 12152 5503 12155
rect 5718 12152 5724 12164
rect 5491 12124 5724 12152
rect 5491 12121 5503 12124
rect 5445 12115 5503 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 7374 12152 7380 12164
rect 6670 12124 7380 12152
rect 7374 12112 7380 12124
rect 7432 12112 7438 12164
rect 8680 12096 8708 12192
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 8812 12192 9137 12220
rect 8812 12180 8818 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9585 12223 9643 12229
rect 9585 12220 9597 12223
rect 9447 12192 9597 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9585 12189 9597 12192
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 12728 12220 12756 12260
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15396 12297 15424 12328
rect 15381 12291 15439 12297
rect 15381 12288 15393 12291
rect 15252 12260 15393 12288
rect 15252 12248 15258 12260
rect 15381 12257 15393 12260
rect 15427 12257 15439 12291
rect 15381 12251 15439 12257
rect 15562 12248 15568 12300
rect 15620 12248 15626 12300
rect 16040 12288 16068 12328
rect 18417 12291 18475 12297
rect 18417 12288 18429 12291
rect 16040 12260 18429 12288
rect 18417 12257 18429 12260
rect 18463 12288 18475 12291
rect 18782 12288 18788 12300
rect 18463 12260 18788 12288
rect 18463 12257 18475 12260
rect 18417 12251 18475 12257
rect 18782 12248 18788 12260
rect 18840 12248 18846 12300
rect 19444 12288 19472 12387
rect 19536 12368 19564 12396
rect 19889 12393 19901 12396
rect 19935 12393 19947 12427
rect 19889 12387 19947 12393
rect 21361 12427 21419 12433
rect 21361 12393 21373 12427
rect 21407 12424 21419 12427
rect 21821 12427 21879 12433
rect 21407 12396 21588 12424
rect 21407 12393 21419 12396
rect 21361 12387 21419 12393
rect 19518 12316 19524 12368
rect 19576 12316 19582 12368
rect 19613 12359 19671 12365
rect 19613 12325 19625 12359
rect 19659 12356 19671 12359
rect 20162 12356 20168 12368
rect 19659 12328 20168 12356
rect 19659 12325 19671 12328
rect 19613 12319 19671 12325
rect 20162 12316 20168 12328
rect 20220 12316 20226 12368
rect 21560 12356 21588 12396
rect 21821 12393 21833 12427
rect 21867 12424 21879 12427
rect 22462 12424 22468 12436
rect 21867 12396 22468 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 22462 12384 22468 12396
rect 22520 12384 22526 12436
rect 22664 12396 23612 12424
rect 22664 12368 22692 12396
rect 21560 12328 22094 12356
rect 21818 12288 21824 12300
rect 19444 12260 19564 12288
rect 11638 12192 12756 12220
rect 10045 12183 10103 12189
rect 10060 12152 10088 12183
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12860 12192 13093 12220
rect 12860 12180 12866 12192
rect 13081 12189 13093 12192
rect 13127 12189 13139 12223
rect 13081 12183 13139 12189
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18138 12220 18144 12232
rect 18003 12192 18144 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 9232 12124 10088 12152
rect 2225 12087 2283 12093
rect 2225 12053 2237 12087
rect 2271 12053 2283 12087
rect 2225 12047 2283 12053
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12084 8815 12087
rect 9232 12084 9260 12124
rect 10502 12112 10508 12164
rect 10560 12112 10566 12164
rect 15948 12152 15976 12183
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 12406 12124 15976 12152
rect 8803 12056 9260 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 9548 12056 9965 12084
rect 9548 12044 9554 12056
rect 9953 12053 9965 12056
rect 9999 12053 10011 12087
rect 9953 12047 10011 12053
rect 11514 12044 11520 12096
rect 11572 12084 11578 12096
rect 12406 12084 12434 12124
rect 16206 12112 16212 12164
rect 16264 12112 16270 12164
rect 19245 12155 19303 12161
rect 16316 12124 16698 12152
rect 11572 12056 12434 12084
rect 11572 12044 11578 12056
rect 12894 12044 12900 12096
rect 12952 12044 12958 12096
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15194 12084 15200 12096
rect 14967 12056 15200 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 15286 12044 15292 12096
rect 15344 12044 15350 12096
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 16316 12084 16344 12124
rect 19245 12121 19257 12155
rect 19291 12152 19303 12155
rect 19334 12152 19340 12164
rect 19291 12124 19340 12152
rect 19291 12121 19303 12124
rect 19245 12115 19303 12121
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 19426 12112 19432 12164
rect 19484 12161 19490 12164
rect 19484 12155 19508 12161
rect 19496 12121 19508 12155
rect 19536 12152 19564 12260
rect 21008 12260 21824 12288
rect 21008 12229 21036 12260
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 22066 12288 22094 12328
rect 22646 12316 22652 12368
rect 22704 12316 22710 12368
rect 23290 12356 23296 12368
rect 22940 12328 23296 12356
rect 22370 12288 22376 12300
rect 22066 12260 22376 12288
rect 22370 12248 22376 12260
rect 22428 12288 22434 12300
rect 22940 12297 22968 12328
rect 23290 12316 23296 12328
rect 23348 12356 23354 12368
rect 23385 12359 23443 12365
rect 23385 12356 23397 12359
rect 23348 12328 23397 12356
rect 23348 12316 23354 12328
rect 23385 12325 23397 12328
rect 23431 12325 23443 12359
rect 23385 12319 23443 12325
rect 23477 12359 23535 12365
rect 23477 12325 23489 12359
rect 23523 12325 23535 12359
rect 23477 12319 23535 12325
rect 22833 12291 22891 12297
rect 22833 12288 22845 12291
rect 22428 12260 22845 12288
rect 22428 12248 22434 12260
rect 22833 12257 22845 12260
rect 22879 12257 22891 12291
rect 22833 12251 22891 12257
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12288 23167 12291
rect 23492 12288 23520 12319
rect 23584 12300 23612 12396
rect 24026 12384 24032 12436
rect 24084 12384 24090 12436
rect 24394 12384 24400 12436
rect 24452 12384 24458 12436
rect 26237 12427 26295 12433
rect 24780 12396 26188 12424
rect 24044 12356 24072 12384
rect 24780 12356 24808 12396
rect 25225 12359 25283 12365
rect 25225 12356 25237 12359
rect 24044 12328 24808 12356
rect 24872 12328 25237 12356
rect 23155 12260 23520 12288
rect 23155 12257 23167 12260
rect 23109 12251 23167 12257
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12189 21051 12223
rect 20993 12183 21051 12189
rect 21361 12223 21419 12229
rect 21361 12189 21373 12223
rect 21407 12220 21419 12223
rect 22940 12220 22968 12251
rect 23566 12248 23572 12300
rect 23624 12248 23630 12300
rect 24872 12297 24900 12328
rect 25225 12325 25237 12328
rect 25271 12325 25283 12359
rect 26160 12356 26188 12396
rect 26237 12393 26249 12427
rect 26283 12424 26295 12427
rect 27614 12424 27620 12436
rect 26283 12396 27620 12424
rect 26283 12393 26295 12396
rect 26237 12387 26295 12393
rect 27614 12384 27620 12396
rect 27672 12384 27678 12436
rect 28629 12427 28687 12433
rect 28629 12393 28641 12427
rect 28675 12424 28687 12427
rect 28810 12424 28816 12436
rect 28675 12396 28816 12424
rect 28675 12393 28687 12396
rect 28629 12387 28687 12393
rect 28810 12384 28816 12396
rect 28868 12384 28874 12436
rect 29454 12424 29460 12436
rect 28920 12396 29460 12424
rect 28920 12356 28948 12396
rect 29454 12384 29460 12396
rect 29512 12384 29518 12436
rect 29546 12384 29552 12436
rect 29604 12424 29610 12436
rect 30190 12424 30196 12436
rect 29604 12396 30196 12424
rect 29604 12384 29610 12396
rect 30190 12384 30196 12396
rect 30248 12384 30254 12436
rect 26160 12328 28948 12356
rect 25225 12319 25283 12325
rect 28994 12316 29000 12368
rect 29052 12356 29058 12368
rect 29052 12328 29868 12356
rect 29052 12316 29058 12328
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12257 24915 12291
rect 24857 12251 24915 12257
rect 25130 12248 25136 12300
rect 25188 12248 25194 12300
rect 25314 12248 25320 12300
rect 25372 12248 25378 12300
rect 25866 12248 25872 12300
rect 25924 12288 25930 12300
rect 26694 12288 26700 12300
rect 25924 12260 26700 12288
rect 25924 12248 25930 12260
rect 26694 12248 26700 12260
rect 26752 12288 26758 12300
rect 26789 12291 26847 12297
rect 26789 12288 26801 12291
rect 26752 12260 26801 12288
rect 26752 12248 26758 12260
rect 26789 12257 26801 12260
rect 26835 12257 26847 12291
rect 26789 12251 26847 12257
rect 26878 12248 26884 12300
rect 26936 12288 26942 12300
rect 27982 12288 27988 12300
rect 26936 12260 27988 12288
rect 26936 12248 26942 12260
rect 27982 12248 27988 12260
rect 28040 12248 28046 12300
rect 29840 12297 29868 12328
rect 30006 12316 30012 12368
rect 30064 12356 30070 12368
rect 30466 12356 30472 12368
rect 30064 12328 30472 12356
rect 30064 12316 30070 12328
rect 30466 12316 30472 12328
rect 30524 12316 30530 12368
rect 29733 12291 29791 12297
rect 29733 12288 29745 12291
rect 28092 12260 29745 12288
rect 21407 12192 22968 12220
rect 23017 12223 23075 12229
rect 21407 12189 21419 12192
rect 21361 12183 21419 12189
rect 21652 12161 21680 12192
rect 23017 12189 23029 12223
rect 23063 12220 23075 12223
rect 23198 12220 23204 12232
rect 23063 12192 23204 12220
rect 23063 12189 23075 12192
rect 23017 12183 23075 12189
rect 23198 12180 23204 12192
rect 23256 12220 23262 12232
rect 23293 12223 23351 12229
rect 23293 12220 23305 12223
rect 23256 12192 23305 12220
rect 23256 12180 23262 12192
rect 23293 12189 23305 12192
rect 23339 12220 23351 12223
rect 23382 12220 23388 12232
rect 23339 12192 23388 12220
rect 23339 12189 23351 12192
rect 23293 12183 23351 12189
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 24302 12180 24308 12232
rect 24360 12220 24366 12232
rect 24578 12220 24584 12232
rect 24360 12192 24584 12220
rect 24360 12180 24366 12192
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 19705 12155 19763 12161
rect 19705 12152 19717 12155
rect 19536 12124 19717 12152
rect 19484 12115 19508 12121
rect 19705 12121 19717 12124
rect 19751 12121 19763 12155
rect 19705 12115 19763 12121
rect 21637 12155 21695 12161
rect 21637 12121 21649 12155
rect 21683 12121 21695 12155
rect 21637 12115 21695 12121
rect 19484 12112 19490 12115
rect 22462 12112 22468 12164
rect 22520 12152 22526 12164
rect 24688 12152 24716 12183
rect 24762 12180 24768 12232
rect 24820 12180 24826 12232
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12220 25099 12223
rect 25682 12220 25688 12232
rect 25087 12192 25688 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 24854 12152 24860 12164
rect 22520 12124 24624 12152
rect 24688 12124 24860 12152
rect 22520 12112 22526 12124
rect 15620 12056 16344 12084
rect 15620 12044 15626 12056
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 19905 12087 19963 12093
rect 19905 12084 19917 12087
rect 18748 12056 19917 12084
rect 18748 12044 18754 12056
rect 19905 12053 19917 12056
rect 19951 12053 19963 12087
rect 19905 12047 19963 12053
rect 20070 12044 20076 12096
rect 20128 12044 20134 12096
rect 21450 12044 21456 12096
rect 21508 12084 21514 12096
rect 21545 12087 21603 12093
rect 21545 12084 21557 12087
rect 21508 12056 21557 12084
rect 21508 12044 21514 12056
rect 21545 12053 21557 12056
rect 21591 12053 21603 12087
rect 21545 12047 21603 12053
rect 21818 12044 21824 12096
rect 21876 12093 21882 12096
rect 21876 12087 21895 12093
rect 21883 12053 21895 12087
rect 21876 12047 21895 12053
rect 22005 12087 22063 12093
rect 22005 12053 22017 12087
rect 22051 12084 22063 12087
rect 22554 12084 22560 12096
rect 22051 12056 22560 12084
rect 22051 12053 22063 12056
rect 22005 12047 22063 12053
rect 21876 12044 21882 12047
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 22649 12087 22707 12093
rect 22649 12053 22661 12087
rect 22695 12084 22707 12087
rect 22922 12084 22928 12096
rect 22695 12056 22928 12084
rect 22695 12053 22707 12056
rect 22649 12047 22707 12053
rect 22922 12044 22928 12056
rect 22980 12044 22986 12096
rect 24596 12084 24624 12124
rect 24854 12112 24860 12124
rect 24912 12112 24918 12164
rect 25056 12084 25084 12183
rect 25682 12180 25688 12192
rect 25740 12180 25746 12232
rect 26326 12180 26332 12232
rect 26384 12220 26390 12232
rect 28092 12220 28120 12260
rect 29733 12257 29745 12260
rect 29779 12257 29791 12291
rect 29733 12251 29791 12257
rect 29825 12291 29883 12297
rect 29825 12257 29837 12291
rect 29871 12288 29883 12291
rect 29871 12260 30788 12288
rect 29871 12257 29883 12260
rect 29825 12251 29883 12257
rect 26384 12192 28120 12220
rect 26384 12180 26390 12192
rect 28902 12180 28908 12232
rect 28960 12180 28966 12232
rect 29273 12223 29331 12229
rect 29273 12189 29285 12223
rect 29319 12189 29331 12223
rect 29273 12183 29331 12189
rect 29365 12223 29423 12229
rect 29365 12189 29377 12223
rect 29411 12220 29423 12223
rect 29454 12220 29460 12232
rect 29411 12192 29460 12220
rect 29411 12189 29423 12192
rect 29365 12183 29423 12189
rect 25958 12112 25964 12164
rect 26016 12152 26022 12164
rect 28997 12155 29055 12161
rect 28997 12152 29009 12155
rect 26016 12124 29009 12152
rect 26016 12112 26022 12124
rect 28997 12121 29009 12124
rect 29043 12121 29055 12155
rect 29288 12152 29316 12183
rect 29454 12180 29460 12192
rect 29512 12180 29518 12232
rect 30190 12180 30196 12232
rect 30248 12180 30254 12232
rect 30558 12180 30564 12232
rect 30616 12180 30622 12232
rect 30760 12229 30788 12260
rect 30745 12223 30803 12229
rect 30745 12189 30757 12223
rect 30791 12189 30803 12223
rect 30745 12183 30803 12189
rect 30576 12152 30604 12180
rect 29288 12124 29868 12152
rect 28997 12115 29055 12121
rect 29840 12096 29868 12124
rect 30024 12124 30604 12152
rect 24596 12056 25084 12084
rect 25774 12044 25780 12096
rect 25832 12084 25838 12096
rect 26605 12087 26663 12093
rect 26605 12084 26617 12087
rect 25832 12056 26617 12084
rect 25832 12044 25838 12056
rect 26605 12053 26617 12056
rect 26651 12053 26663 12087
rect 26605 12047 26663 12053
rect 26694 12044 26700 12096
rect 26752 12044 26758 12096
rect 29089 12087 29147 12093
rect 29089 12053 29101 12087
rect 29135 12084 29147 12087
rect 29270 12084 29276 12096
rect 29135 12056 29276 12084
rect 29135 12053 29147 12056
rect 29089 12047 29147 12053
rect 29270 12044 29276 12056
rect 29328 12044 29334 12096
rect 29822 12044 29828 12096
rect 29880 12044 29886 12096
rect 30024 12093 30052 12124
rect 30009 12087 30067 12093
rect 30009 12053 30021 12087
rect 30055 12053 30067 12087
rect 30009 12047 30067 12053
rect 30098 12044 30104 12096
rect 30156 12044 30162 12096
rect 30650 12044 30656 12096
rect 30708 12044 30714 12096
rect 1104 11994 38272 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38272 11994
rect 1104 11920 38272 11942
rect 1762 11840 1768 11892
rect 1820 11840 1826 11892
rect 3145 11883 3203 11889
rect 3145 11849 3157 11883
rect 3191 11880 3203 11883
rect 3418 11880 3424 11892
rect 3191 11852 3424 11880
rect 3191 11849 3203 11852
rect 3145 11843 3203 11849
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 5997 11883 6055 11889
rect 5997 11849 6009 11883
rect 6043 11880 6055 11883
rect 6043 11852 6684 11880
rect 6043 11849 6055 11852
rect 5997 11843 6055 11849
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 1780 11812 1808 11840
rect 6656 11821 6684 11852
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 9398 11880 9404 11892
rect 8720 11852 9404 11880
rect 8720 11840 8726 11852
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 12894 11840 12900 11892
rect 12952 11880 12958 11892
rect 15010 11880 15016 11892
rect 12952 11852 13216 11880
rect 12952 11840 12958 11852
rect 1719 11784 1808 11812
rect 6641 11815 6699 11821
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 6641 11781 6653 11815
rect 6687 11781 6699 11815
rect 6641 11775 6699 11781
rect 7374 11772 7380 11824
rect 7432 11772 7438 11824
rect 9214 11812 9220 11824
rect 8496 11784 9220 11812
rect 1394 11704 1400 11756
rect 1452 11704 1458 11756
rect 2958 11744 2964 11756
rect 2806 11716 2964 11744
rect 2958 11704 2964 11716
rect 3016 11744 3022 11756
rect 3786 11744 3792 11756
rect 3016 11716 3792 11744
rect 3016 11704 3022 11716
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 6086 11704 6092 11756
rect 6144 11704 6150 11756
rect 6178 11704 6184 11756
rect 6236 11704 6242 11756
rect 8496 11753 8524 11784
rect 9214 11772 9220 11784
rect 9272 11812 9278 11824
rect 9950 11812 9956 11824
rect 9272 11784 9956 11812
rect 9272 11772 9278 11784
rect 9950 11772 9956 11784
rect 10008 11812 10014 11824
rect 12342 11812 12348 11824
rect 10008 11784 12348 11812
rect 10008 11772 10014 11784
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 13188 11821 13216 11852
rect 13556 11852 15016 11880
rect 13173 11815 13231 11821
rect 13173 11781 13185 11815
rect 13219 11781 13231 11815
rect 13173 11775 13231 11781
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 13556 11812 13584 11852
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 15194 11840 15200 11892
rect 15252 11840 15258 11892
rect 15473 11883 15531 11889
rect 15473 11849 15485 11883
rect 15519 11880 15531 11883
rect 16206 11880 16212 11892
rect 15519 11852 16212 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 21174 11880 21180 11892
rect 19536 11852 21180 11880
rect 13320 11784 13662 11812
rect 13320 11772 13326 11784
rect 14918 11772 14924 11824
rect 14976 11772 14982 11824
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 8904 11716 9137 11744
rect 8904 11704 8910 11716
rect 9125 11713 9137 11716
rect 9171 11744 9183 11747
rect 9582 11744 9588 11756
rect 9171 11716 9588 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 11146 11704 11152 11756
rect 11204 11744 11210 11756
rect 12066 11744 12072 11756
rect 11204 11716 12072 11744
rect 11204 11704 11210 11716
rect 12066 11704 12072 11716
rect 12124 11744 12130 11756
rect 15212 11744 15240 11840
rect 17678 11772 17684 11824
rect 17736 11812 17742 11824
rect 17736 11784 17908 11812
rect 17736 11772 17742 11784
rect 17880 11753 17908 11784
rect 19536 11753 19564 11852
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 21450 11840 21456 11892
rect 21508 11840 21514 11892
rect 24213 11883 24271 11889
rect 24213 11849 24225 11883
rect 24259 11880 24271 11883
rect 24762 11880 24768 11892
rect 24259 11852 24768 11880
rect 24259 11849 24271 11852
rect 24213 11843 24271 11849
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 25041 11883 25099 11889
rect 25041 11849 25053 11883
rect 25087 11880 25099 11883
rect 25314 11880 25320 11892
rect 25087 11852 25320 11880
rect 25087 11849 25099 11852
rect 25041 11843 25099 11849
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 25501 11883 25559 11889
rect 25501 11849 25513 11883
rect 25547 11880 25559 11883
rect 25774 11880 25780 11892
rect 25547 11852 25780 11880
rect 25547 11849 25559 11852
rect 25501 11843 25559 11849
rect 25774 11840 25780 11852
rect 25832 11840 25838 11892
rect 28626 11880 28632 11892
rect 26988 11852 28632 11880
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 12124 11716 12572 11744
rect 15212 11716 15669 11744
rect 12124 11704 12130 11716
rect 6104 11676 6132 11704
rect 6365 11679 6423 11685
rect 6365 11676 6377 11679
rect 6104 11648 6377 11676
rect 6365 11645 6377 11648
rect 6411 11645 6423 11679
rect 6365 11639 6423 11645
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 8110 11676 8116 11688
rect 7156 11648 8116 11676
rect 7156 11636 7162 11648
rect 8110 11636 8116 11648
rect 8168 11676 8174 11688
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8168 11648 8401 11676
rect 8168 11636 8174 11648
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8389 11639 8447 11645
rect 8680 11648 8769 11676
rect 8680 11552 8708 11648
rect 8757 11645 8769 11648
rect 8803 11676 8815 11679
rect 9766 11676 9772 11688
rect 8803 11648 9772 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 12434 11636 12440 11688
rect 12492 11636 12498 11688
rect 12544 11685 12572 11716
rect 15657 11713 15669 11716
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 19610 11704 19616 11756
rect 19668 11704 19674 11756
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11744 19947 11747
rect 19978 11744 19984 11756
rect 19935 11716 19984 11744
rect 19935 11713 19947 11716
rect 19889 11707 19947 11713
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 9490 11608 9496 11620
rect 8772 11580 9496 11608
rect 8772 11552 8800 11580
rect 9490 11568 9496 11580
rect 9548 11608 9554 11620
rect 9585 11611 9643 11617
rect 9585 11608 9597 11611
rect 9548 11580 9597 11608
rect 9548 11568 9554 11580
rect 9585 11577 9597 11580
rect 9631 11577 9643 11611
rect 9585 11571 9643 11577
rect 8662 11500 8668 11552
rect 8720 11500 8726 11552
rect 8754 11500 8760 11552
rect 8812 11500 8818 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8996 11512 9045 11540
rect 8996 11500 9002 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 9033 11503 9091 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10410 11540 10416 11552
rect 9456 11512 10416 11540
rect 9456 11500 9462 11512
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 12802 11540 12808 11552
rect 12308 11512 12808 11540
rect 12308 11500 12314 11512
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 12912 11540 12940 11639
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 19720 11676 19748 11707
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 21468 11744 21496 11840
rect 26988 11824 27016 11852
rect 28626 11840 28632 11852
rect 28684 11840 28690 11892
rect 28902 11840 28908 11892
rect 28960 11840 28966 11892
rect 29270 11840 29276 11892
rect 29328 11880 29334 11892
rect 29365 11883 29423 11889
rect 29365 11880 29377 11883
rect 29328 11852 29377 11880
rect 29328 11840 29334 11852
rect 29365 11849 29377 11852
rect 29411 11849 29423 11883
rect 29365 11843 29423 11849
rect 29822 11840 29828 11892
rect 29880 11880 29886 11892
rect 30009 11883 30067 11889
rect 30009 11880 30021 11883
rect 29880 11852 30021 11880
rect 29880 11840 29886 11852
rect 30009 11849 30021 11852
rect 30055 11880 30067 11883
rect 31202 11880 31208 11892
rect 30055 11852 31208 11880
rect 30055 11849 30067 11852
rect 30009 11843 30067 11849
rect 31202 11840 31208 11852
rect 31260 11840 31266 11892
rect 32950 11840 32956 11892
rect 33008 11880 33014 11892
rect 33008 11852 33640 11880
rect 33008 11840 33014 11852
rect 24486 11812 24492 11824
rect 24412 11784 24492 11812
rect 21223 11716 21496 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 22646 11704 22652 11756
rect 22704 11704 22710 11756
rect 22925 11747 22983 11753
rect 22925 11713 22937 11747
rect 22971 11744 22983 11747
rect 22971 11716 23337 11744
rect 22971 11713 22983 11716
rect 22925 11707 22983 11713
rect 13964 11648 19748 11676
rect 13964 11636 13970 11648
rect 21818 11636 21824 11688
rect 21876 11676 21882 11688
rect 22278 11676 22284 11688
rect 21876 11648 22284 11676
rect 21876 11636 21882 11648
rect 22278 11636 22284 11648
rect 22336 11676 22342 11688
rect 22940 11676 22968 11707
rect 22336 11648 22968 11676
rect 22336 11636 22342 11648
rect 19242 11568 19248 11620
rect 19300 11568 19306 11620
rect 21361 11611 21419 11617
rect 21361 11577 21373 11611
rect 21407 11608 21419 11611
rect 22462 11608 22468 11620
rect 21407 11580 22468 11608
rect 21407 11577 21419 11580
rect 21361 11571 21419 11577
rect 22462 11568 22468 11580
rect 22520 11568 22526 11620
rect 23309 11608 23337 11716
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 24029 11747 24087 11753
rect 24029 11744 24041 11747
rect 23440 11716 24041 11744
rect 23440 11704 23446 11716
rect 24029 11713 24041 11716
rect 24075 11713 24087 11747
rect 24029 11707 24087 11713
rect 24044 11676 24072 11707
rect 24302 11704 24308 11756
rect 24360 11704 24366 11756
rect 24412 11753 24440 11784
rect 24486 11772 24492 11784
rect 24544 11772 24550 11824
rect 24670 11812 24676 11824
rect 24596 11784 24676 11812
rect 24596 11753 24624 11784
rect 24670 11772 24676 11784
rect 24728 11812 24734 11824
rect 24728 11784 25636 11812
rect 24728 11772 24734 11784
rect 24397 11747 24455 11753
rect 24397 11713 24409 11747
rect 24443 11713 24455 11747
rect 24397 11707 24455 11713
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11713 24639 11747
rect 25409 11747 25467 11753
rect 25409 11744 25421 11747
rect 24581 11707 24639 11713
rect 25332 11716 25421 11744
rect 24489 11679 24547 11685
rect 24489 11676 24501 11679
rect 24044 11648 24501 11676
rect 24489 11645 24501 11648
rect 24535 11645 24547 11679
rect 24489 11639 24547 11645
rect 25332 11620 25360 11716
rect 25409 11713 25421 11716
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 25608 11685 25636 11784
rect 26786 11772 26792 11824
rect 26844 11812 26850 11824
rect 26970 11812 26976 11824
rect 26844 11784 26976 11812
rect 26844 11772 26850 11784
rect 26970 11772 26976 11784
rect 27028 11772 27034 11824
rect 27246 11821 27252 11824
rect 27189 11815 27252 11821
rect 27189 11781 27201 11815
rect 27235 11781 27252 11815
rect 27189 11775 27252 11781
rect 27246 11772 27252 11775
rect 27304 11772 27310 11824
rect 26878 11704 26884 11756
rect 26936 11744 26942 11756
rect 27338 11744 27344 11756
rect 26936 11716 27344 11744
rect 26936 11704 26942 11716
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 25593 11679 25651 11685
rect 25593 11645 25605 11679
rect 25639 11645 25651 11679
rect 28920 11676 28948 11840
rect 30653 11815 30711 11821
rect 30653 11812 30665 11815
rect 25593 11639 25651 11645
rect 26436 11648 28948 11676
rect 29012 11784 30665 11812
rect 24854 11608 24860 11620
rect 23309 11580 24860 11608
rect 24854 11568 24860 11580
rect 24912 11568 24918 11620
rect 25314 11568 25320 11620
rect 25372 11568 25378 11620
rect 14642 11540 14648 11552
rect 12912 11512 14648 11540
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15562 11540 15568 11552
rect 15068 11512 15568 11540
rect 15068 11500 15074 11512
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 17954 11500 17960 11552
rect 18012 11500 18018 11552
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 22002 11540 22008 11552
rect 20036 11512 22008 11540
rect 20036 11500 20042 11512
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 22741 11543 22799 11549
rect 22741 11509 22753 11543
rect 22787 11540 22799 11543
rect 22922 11540 22928 11552
rect 22787 11512 22928 11540
rect 22787 11509 22799 11512
rect 22741 11503 22799 11509
rect 22922 11500 22928 11512
rect 22980 11500 22986 11552
rect 24029 11543 24087 11549
rect 24029 11509 24041 11543
rect 24075 11540 24087 11543
rect 26436 11540 26464 11648
rect 27341 11611 27399 11617
rect 27341 11608 27353 11611
rect 26988 11580 27353 11608
rect 26988 11552 27016 11580
rect 27341 11577 27353 11580
rect 27387 11608 27399 11611
rect 27522 11608 27528 11620
rect 27387 11580 27528 11608
rect 27387 11577 27399 11580
rect 27341 11571 27399 11577
rect 27522 11568 27528 11580
rect 27580 11568 27586 11620
rect 27798 11568 27804 11620
rect 27856 11608 27862 11620
rect 29012 11608 29040 11784
rect 30653 11781 30665 11784
rect 30699 11781 30711 11815
rect 30653 11775 30711 11781
rect 32876 11784 33364 11812
rect 29086 11704 29092 11756
rect 29144 11704 29150 11756
rect 29181 11747 29239 11753
rect 29181 11713 29193 11747
rect 29227 11744 29239 11747
rect 29546 11744 29552 11756
rect 29227 11716 29552 11744
rect 29227 11713 29239 11716
rect 29181 11707 29239 11713
rect 29546 11704 29552 11716
rect 29604 11704 29610 11756
rect 30469 11747 30527 11753
rect 30116 11716 30328 11744
rect 29365 11679 29423 11685
rect 29365 11645 29377 11679
rect 29411 11676 29423 11679
rect 30006 11676 30012 11688
rect 29411 11648 30012 11676
rect 29411 11645 29423 11648
rect 29365 11639 29423 11645
rect 27856 11580 29040 11608
rect 27856 11568 27862 11580
rect 24075 11512 26464 11540
rect 24075 11509 24087 11512
rect 24029 11503 24087 11509
rect 26970 11500 26976 11552
rect 27028 11500 27034 11552
rect 27154 11500 27160 11552
rect 27212 11500 27218 11552
rect 28718 11500 28724 11552
rect 28776 11540 28782 11552
rect 29380 11540 29408 11639
rect 30006 11636 30012 11648
rect 30064 11636 30070 11688
rect 28776 11512 29408 11540
rect 30116 11540 30144 11716
rect 30300 11685 30328 11716
rect 30469 11713 30481 11747
rect 30515 11744 30527 11747
rect 31297 11747 31355 11753
rect 31297 11744 31309 11747
rect 30515 11716 31309 11744
rect 30515 11713 30527 11716
rect 30469 11707 30527 11713
rect 31297 11713 31309 11716
rect 31343 11713 31355 11747
rect 31297 11707 31355 11713
rect 31386 11704 31392 11756
rect 31444 11744 31450 11756
rect 32876 11753 32904 11784
rect 33336 11753 33364 11784
rect 33612 11753 33640 11852
rect 32861 11747 32919 11753
rect 32861 11744 32873 11747
rect 31444 11716 32873 11744
rect 31444 11704 31450 11716
rect 32861 11713 32873 11716
rect 32907 11713 32919 11747
rect 32861 11707 32919 11713
rect 33045 11747 33103 11753
rect 33045 11713 33057 11747
rect 33091 11713 33103 11747
rect 33045 11707 33103 11713
rect 33321 11747 33379 11753
rect 33321 11713 33333 11747
rect 33367 11713 33379 11747
rect 33321 11707 33379 11713
rect 33597 11747 33655 11753
rect 33597 11713 33609 11747
rect 33643 11713 33655 11747
rect 33597 11707 33655 11713
rect 30193 11679 30251 11685
rect 30193 11645 30205 11679
rect 30239 11645 30251 11679
rect 30193 11639 30251 11645
rect 30285 11679 30343 11685
rect 30285 11645 30297 11679
rect 30331 11645 30343 11679
rect 30285 11639 30343 11645
rect 30377 11679 30435 11685
rect 30377 11645 30389 11679
rect 30423 11676 30435 11679
rect 30558 11676 30564 11688
rect 30423 11648 30564 11676
rect 30423 11645 30435 11648
rect 30377 11639 30435 11645
rect 30208 11608 30236 11639
rect 30558 11636 30564 11648
rect 30616 11636 30622 11688
rect 30650 11636 30656 11688
rect 30708 11676 30714 11688
rect 31021 11679 31079 11685
rect 31021 11676 31033 11679
rect 30708 11648 31033 11676
rect 30708 11636 30714 11648
rect 31021 11645 31033 11648
rect 31067 11645 31079 11679
rect 31021 11639 31079 11645
rect 31110 11636 31116 11688
rect 31168 11636 31174 11688
rect 33060 11676 33088 11707
rect 33778 11704 33784 11756
rect 33836 11704 33842 11756
rect 33137 11679 33195 11685
rect 33137 11676 33149 11679
rect 33060 11648 33149 11676
rect 33137 11645 33149 11648
rect 33183 11676 33195 11679
rect 33226 11676 33232 11688
rect 33183 11648 33232 11676
rect 33183 11645 33195 11648
rect 33137 11639 33195 11645
rect 33226 11636 33232 11648
rect 33284 11636 33290 11688
rect 33796 11676 33824 11704
rect 33520 11648 33824 11676
rect 30668 11608 30696 11636
rect 30208 11580 30696 11608
rect 30466 11540 30472 11552
rect 30116 11512 30472 11540
rect 28776 11500 28782 11512
rect 30466 11500 30472 11512
rect 30524 11500 30530 11552
rect 32030 11500 32036 11552
rect 32088 11540 32094 11552
rect 33520 11549 33548 11648
rect 33870 11568 33876 11620
rect 33928 11568 33934 11620
rect 33505 11543 33563 11549
rect 33505 11540 33517 11543
rect 32088 11512 33517 11540
rect 32088 11500 32094 11512
rect 33505 11509 33517 11512
rect 33551 11509 33563 11543
rect 33505 11503 33563 11509
rect 1104 11450 38272 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38272 11450
rect 1104 11376 38272 11398
rect 1688 11308 4016 11336
rect 1688 11277 1716 11308
rect 1673 11271 1731 11277
rect 1673 11237 1685 11271
rect 1719 11237 1731 11271
rect 1673 11231 1731 11237
rect 3789 11271 3847 11277
rect 3789 11237 3801 11271
rect 3835 11237 3847 11271
rect 3988 11268 4016 11308
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 5258 11336 5264 11348
rect 4120 11308 5264 11336
rect 4120 11296 4126 11308
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 6641 11339 6699 11345
rect 6641 11336 6653 11339
rect 6236 11308 6653 11336
rect 6236 11296 6242 11308
rect 6641 11305 6653 11308
rect 6687 11305 6699 11339
rect 6641 11299 6699 11305
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 10045 11339 10103 11345
rect 10045 11336 10057 11339
rect 8260 11308 10057 11336
rect 8260 11296 8266 11308
rect 3988 11240 8064 11268
rect 3789 11231 3847 11237
rect 2774 11200 2780 11212
rect 2516 11172 2780 11200
rect 934 11092 940 11144
rect 992 11132 998 11144
rect 2516 11141 2544 11172
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 1489 11135 1547 11141
rect 1489 11132 1501 11135
rect 992 11104 1501 11132
rect 992 11092 998 11104
rect 1489 11101 1501 11104
rect 1535 11101 1547 11135
rect 1489 11095 1547 11101
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 3421 11135 3479 11141
rect 2501 11095 2559 11101
rect 2608 11104 3372 11132
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 2608 11064 2636 11104
rect 2363 11036 2636 11064
rect 2685 11067 2743 11073
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 2685 11033 2697 11067
rect 2731 11064 2743 11067
rect 2958 11064 2964 11076
rect 2731 11036 2964 11064
rect 2731 11033 2743 11036
rect 2685 11027 2743 11033
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 3344 11064 3372 11104
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3804 11132 3832 11231
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 3936 11172 4353 11200
rect 3936 11160 3942 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 4540 11172 4844 11200
rect 4540 11144 4568 11172
rect 4430 11132 4436 11144
rect 3467 11104 3832 11132
rect 3896 11104 4436 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3896 11064 3924 11104
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 4522 11092 4528 11144
rect 4580 11092 4586 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4706 11132 4712 11144
rect 4663 11104 4712 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 4816 11141 4844 11172
rect 7098 11160 7104 11212
rect 7156 11160 7162 11212
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 7374 11132 7380 11144
rect 5408 11104 7380 11132
rect 5408 11092 5414 11104
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 8036 11132 8064 11240
rect 8956 11200 8984 11308
rect 10045 11305 10057 11308
rect 10091 11336 10103 11339
rect 12250 11336 12256 11348
rect 10091 11308 12256 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 13262 11336 13268 11348
rect 12492 11308 13268 11336
rect 12492 11296 12498 11308
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 14182 11296 14188 11348
rect 14240 11296 14246 11348
rect 15286 11336 15292 11348
rect 14292 11308 15292 11336
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9585 11271 9643 11277
rect 9585 11268 9597 11271
rect 9088 11240 9597 11268
rect 9088 11228 9094 11240
rect 9585 11237 9597 11240
rect 9631 11237 9643 11271
rect 9585 11231 9643 11237
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 14292 11268 14320 11308
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 20162 11296 20168 11348
rect 20220 11296 20226 11348
rect 20622 11336 20628 11348
rect 20272 11308 20628 11336
rect 12860 11240 14320 11268
rect 14553 11271 14611 11277
rect 12860 11228 12866 11240
rect 14553 11237 14565 11271
rect 14599 11268 14611 11271
rect 14599 11240 15608 11268
rect 14599 11237 14611 11240
rect 14553 11231 14611 11237
rect 13725 11203 13783 11209
rect 13725 11200 13737 11203
rect 8956 11172 9260 11200
rect 8662 11132 8668 11144
rect 8036 11104 8668 11132
rect 8662 11092 8668 11104
rect 8720 11132 8726 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8720 11104 8953 11132
rect 8720 11092 8726 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 9232 11132 9260 11172
rect 9784 11172 10732 11200
rect 9426 11135 9484 11141
rect 9426 11132 9438 11135
rect 9232 11104 9438 11132
rect 8941 11095 8999 11101
rect 9426 11101 9438 11104
rect 9472 11101 9484 11135
rect 9426 11095 9484 11101
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9640 11104 9689 11132
rect 9640 11092 9646 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 3344 11036 3924 11064
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 7009 11067 7067 11073
rect 4203 11036 4936 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4908 11008 4936 11036
rect 7009 11033 7021 11067
rect 7055 11064 7067 11067
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 7055 11036 9321 11064
rect 7055 11033 7067 11036
rect 7009 11027 7067 11033
rect 9309 11033 9321 11036
rect 9355 11064 9367 11067
rect 9784 11064 9812 11172
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11132 9919 11135
rect 10042 11132 10048 11144
rect 9907 11104 10048 11132
rect 9907 11101 9919 11104
rect 9861 11095 9919 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10410 11092 10416 11144
rect 10468 11092 10474 11144
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 9355 11036 9812 11064
rect 10060 11064 10088 11092
rect 10520 11064 10548 11095
rect 10060 11036 10548 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 3234 10956 3240 11008
rect 3292 10956 3298 11008
rect 4249 10999 4307 11005
rect 4249 10965 4261 10999
rect 4295 10996 4307 10999
rect 4614 10996 4620 11008
rect 4295 10968 4620 10996
rect 4295 10965 4307 10968
rect 4249 10959 4307 10965
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 4706 10956 4712 11008
rect 4764 10956 4770 11008
rect 4890 10956 4896 11008
rect 4948 10956 4954 11008
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 10704 11005 10732 11172
rect 12820 11172 13737 11200
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11514 11132 11520 11144
rect 11112 11104 11520 11132
rect 11112 11092 11118 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 12820 11076 12848 11172
rect 13725 11169 13737 11172
rect 13771 11169 13783 11203
rect 13725 11163 13783 11169
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11200 15255 11203
rect 15378 11200 15384 11212
rect 15243 11172 15384 11200
rect 15243 11169 15255 11172
rect 15197 11163 15255 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 13354 11092 13360 11144
rect 13412 11092 13418 11144
rect 13446 11092 13452 11144
rect 13504 11092 13510 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13924 11104 14105 11132
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 12802 11024 12808 11076
rect 12860 11024 12866 11076
rect 13372 11064 13400 11092
rect 13722 11064 13728 11076
rect 13372 11036 13728 11064
rect 13722 11024 13728 11036
rect 13780 11064 13786 11076
rect 13924 11064 13952 11104
rect 14093 11101 14105 11104
rect 14139 11132 14151 11135
rect 14918 11132 14924 11144
rect 14139 11104 14924 11132
rect 14139 11101 14151 11104
rect 14093 11095 14151 11101
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11132 15071 11135
rect 15470 11132 15476 11144
rect 15059 11104 15476 11132
rect 15059 11101 15071 11104
rect 15013 11095 15071 11101
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15580 11141 15608 11240
rect 18064 11172 18736 11200
rect 18064 11144 18092 11172
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 17310 11092 17316 11144
rect 17368 11092 17374 11144
rect 17678 11092 17684 11144
rect 17736 11132 17742 11144
rect 18046 11132 18052 11144
rect 17736 11104 18052 11132
rect 17736 11092 17742 11104
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18230 11092 18236 11144
rect 18288 11092 18294 11144
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 18708 11141 18736 11172
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11101 18751 11135
rect 19426 11132 19432 11144
rect 18693 11095 18751 11101
rect 18800 11104 19432 11132
rect 13780 11036 13952 11064
rect 15488 11064 15516 11092
rect 17586 11064 17592 11076
rect 15488 11036 17592 11064
rect 13780 11024 13786 11036
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 18417 11067 18475 11073
rect 18417 11033 18429 11067
rect 18463 11064 18475 11067
rect 18800 11064 18828 11104
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 20180 11132 20208 11296
rect 20272 11280 20300 11308
rect 20622 11296 20628 11308
rect 20680 11336 20686 11348
rect 24489 11339 24547 11345
rect 20680 11308 24446 11336
rect 20680 11296 20686 11308
rect 20254 11228 20260 11280
rect 20312 11228 20318 11280
rect 20898 11228 20904 11280
rect 20956 11268 20962 11280
rect 21634 11268 21640 11280
rect 20956 11240 21640 11268
rect 20956 11228 20962 11240
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 24418 11200 24446 11308
rect 24489 11305 24501 11339
rect 24535 11336 24547 11339
rect 25314 11336 25320 11348
rect 24535 11308 25320 11336
rect 24535 11305 24547 11308
rect 24489 11299 24547 11305
rect 25314 11296 25320 11308
rect 25372 11296 25378 11348
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 27154 11336 27160 11348
rect 25547 11308 27160 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 27154 11296 27160 11308
rect 27212 11296 27218 11348
rect 27246 11296 27252 11348
rect 27304 11296 27310 11348
rect 27430 11296 27436 11348
rect 27488 11336 27494 11348
rect 27617 11339 27675 11345
rect 27617 11336 27629 11339
rect 27488 11308 27629 11336
rect 27488 11296 27494 11308
rect 27617 11305 27629 11308
rect 27663 11336 27675 11339
rect 29549 11339 29607 11345
rect 27663 11308 28488 11336
rect 27663 11305 27675 11308
rect 27617 11299 27675 11305
rect 25332 11268 25360 11296
rect 26694 11268 26700 11280
rect 25332 11240 26700 11268
rect 24418 11172 25452 11200
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 20180 11104 20269 11132
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 23566 11092 23572 11144
rect 23624 11132 23630 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 23624 11104 24409 11132
rect 23624 11092 23630 11104
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 24946 11132 24952 11144
rect 24627 11104 24952 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 18463 11036 18828 11064
rect 18877 11067 18935 11073
rect 18463 11033 18475 11036
rect 18417 11027 18475 11033
rect 18877 11033 18889 11067
rect 18923 11064 18935 11067
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 18923 11036 19257 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 19245 11033 19257 11036
rect 19291 11033 19303 11067
rect 19245 11027 19303 11033
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 19981 11067 20039 11073
rect 19981 11064 19993 11067
rect 19392 11036 19993 11064
rect 19392 11024 19398 11036
rect 19981 11033 19993 11036
rect 20027 11064 20039 11067
rect 20027 11036 23060 11064
rect 20027 11033 20039 11036
rect 19981 11027 20039 11033
rect 9217 10999 9275 11005
rect 9217 10996 9229 10999
rect 8720 10968 9229 10996
rect 8720 10956 8726 10968
rect 9217 10965 9229 10968
rect 9263 10965 9275 10999
rect 9217 10959 9275 10965
rect 10689 10999 10747 11005
rect 10689 10965 10701 10999
rect 10735 10996 10747 10999
rect 12434 10996 12440 11008
rect 10735 10968 12440 10996
rect 10735 10965 10747 10968
rect 10689 10959 10747 10965
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 14921 10999 14979 11005
rect 14921 10996 14933 10999
rect 14148 10968 14933 10996
rect 14148 10956 14154 10968
rect 14921 10965 14933 10968
rect 14967 10965 14979 10999
rect 14921 10959 14979 10965
rect 15381 10999 15439 11005
rect 15381 10965 15393 10999
rect 15427 10996 15439 10999
rect 15654 10996 15660 11008
rect 15427 10968 15660 10996
rect 15427 10965 15439 10968
rect 15381 10959 15439 10965
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 17604 10996 17632 11024
rect 18966 10996 18972 11008
rect 17604 10968 18972 10996
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 20162 10956 20168 11008
rect 20220 10996 20226 11008
rect 20441 10999 20499 11005
rect 20441 10996 20453 10999
rect 20220 10968 20453 10996
rect 20220 10956 20226 10968
rect 20441 10965 20453 10968
rect 20487 10965 20499 10999
rect 23032 10996 23060 11036
rect 23290 11024 23296 11076
rect 23348 11064 23354 11076
rect 24596 11064 24624 11095
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 25424 11141 25452 11172
rect 25409 11135 25467 11141
rect 25409 11101 25421 11135
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 25590 11092 25596 11144
rect 25648 11092 25654 11144
rect 25685 11135 25743 11141
rect 25685 11101 25697 11135
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 25700 11064 25728 11095
rect 25866 11092 25872 11144
rect 25924 11092 25930 11144
rect 26620 11141 26648 11240
rect 26694 11228 26700 11240
rect 26752 11228 26758 11280
rect 26786 11160 26792 11212
rect 26844 11160 26850 11212
rect 27264 11200 27292 11296
rect 27338 11228 27344 11280
rect 27396 11268 27402 11280
rect 27396 11240 28396 11268
rect 27396 11228 27402 11240
rect 27264 11172 28212 11200
rect 26605 11135 26663 11141
rect 26605 11101 26617 11135
rect 26651 11101 26663 11135
rect 26804 11132 26832 11160
rect 27154 11132 27160 11144
rect 26804 11104 27160 11132
rect 26605 11095 26663 11101
rect 27154 11092 27160 11104
rect 27212 11132 27218 11144
rect 27249 11135 27307 11141
rect 27249 11132 27261 11135
rect 27212 11104 27261 11132
rect 27212 11092 27218 11104
rect 27249 11101 27261 11104
rect 27295 11101 27307 11135
rect 27249 11095 27307 11101
rect 27338 11092 27344 11144
rect 27396 11132 27402 11144
rect 27540 11141 27568 11172
rect 27433 11135 27491 11141
rect 27433 11132 27445 11135
rect 27396 11104 27445 11132
rect 27396 11092 27402 11104
rect 27433 11101 27445 11104
rect 27479 11101 27491 11135
rect 27433 11095 27491 11101
rect 27525 11135 27583 11141
rect 27525 11101 27537 11135
rect 27571 11101 27583 11135
rect 27525 11095 27583 11101
rect 27614 11092 27620 11144
rect 27672 11132 27678 11144
rect 28184 11141 28212 11172
rect 28368 11141 28396 11240
rect 27801 11135 27859 11141
rect 27801 11132 27813 11135
rect 27672 11104 27813 11132
rect 27672 11092 27678 11104
rect 27801 11101 27813 11104
rect 27847 11101 27859 11135
rect 27801 11095 27859 11101
rect 28077 11135 28135 11141
rect 28077 11101 28089 11135
rect 28123 11101 28135 11135
rect 28077 11095 28135 11101
rect 28169 11135 28227 11141
rect 28169 11101 28181 11135
rect 28215 11101 28227 11135
rect 28169 11095 28227 11101
rect 28353 11135 28411 11141
rect 28353 11101 28365 11135
rect 28399 11101 28411 11135
rect 28460 11132 28488 11308
rect 29549 11305 29561 11339
rect 29595 11336 29607 11339
rect 29730 11336 29736 11348
rect 29595 11308 29736 11336
rect 29595 11305 29607 11308
rect 29549 11299 29607 11305
rect 29730 11296 29736 11308
rect 29788 11296 29794 11348
rect 31110 11296 31116 11348
rect 31168 11336 31174 11348
rect 31849 11339 31907 11345
rect 31849 11336 31861 11339
rect 31168 11308 31861 11336
rect 31168 11296 31174 11308
rect 31849 11305 31861 11308
rect 31895 11305 31907 11339
rect 31849 11299 31907 11305
rect 32582 11296 32588 11348
rect 32640 11296 32646 11348
rect 28626 11228 28632 11280
rect 28684 11268 28690 11280
rect 33226 11268 33232 11280
rect 28684 11240 33232 11268
rect 28684 11228 28690 11240
rect 33226 11228 33232 11240
rect 33284 11228 33290 11280
rect 32950 11160 32956 11212
rect 33008 11160 33014 11212
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 28460 11104 29745 11132
rect 28353 11095 28411 11101
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 23348 11036 24624 11064
rect 24688 11036 25728 11064
rect 23348 11024 23354 11036
rect 23474 10996 23480 11008
rect 23032 10968 23480 10996
rect 20441 10959 20499 10965
rect 23474 10956 23480 10968
rect 23532 10996 23538 11008
rect 23842 10996 23848 11008
rect 23532 10968 23848 10996
rect 23532 10956 23538 10968
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 24302 10956 24308 11008
rect 24360 10996 24366 11008
rect 24688 10996 24716 11036
rect 25774 11024 25780 11076
rect 25832 11064 25838 11076
rect 27065 11067 27123 11073
rect 25832 11036 26740 11064
rect 25832 11024 25838 11036
rect 24360 10968 24716 10996
rect 24360 10956 24366 10968
rect 25866 10956 25872 11008
rect 25924 10956 25930 11008
rect 26234 10956 26240 11008
rect 26292 10956 26298 11008
rect 26712 11005 26740 11036
rect 27065 11033 27077 11067
rect 27111 11064 27123 11067
rect 27985 11067 28043 11073
rect 27985 11064 27997 11067
rect 27111 11036 27997 11064
rect 27111 11033 27123 11036
rect 27065 11027 27123 11033
rect 27540 11008 27568 11036
rect 27985 11033 27997 11036
rect 28031 11033 28043 11067
rect 27985 11027 28043 11033
rect 26697 10999 26755 11005
rect 26697 10965 26709 10999
rect 26743 10965 26755 10999
rect 26697 10959 26755 10965
rect 27522 10956 27528 11008
rect 27580 10956 27586 11008
rect 27706 10956 27712 11008
rect 27764 10996 27770 11008
rect 28092 10996 28120 11095
rect 29914 11092 29920 11144
rect 29972 11092 29978 11144
rect 30009 11135 30067 11141
rect 30009 11101 30021 11135
rect 30055 11132 30067 11135
rect 30558 11132 30564 11144
rect 30055 11104 30564 11132
rect 30055 11101 30067 11104
rect 30009 11095 30067 11101
rect 30558 11092 30564 11104
rect 30616 11092 30622 11144
rect 31386 11092 31392 11144
rect 31444 11092 31450 11144
rect 32030 11092 32036 11144
rect 32088 11092 32094 11144
rect 32306 11092 32312 11144
rect 32364 11092 32370 11144
rect 32493 11135 32551 11141
rect 32493 11101 32505 11135
rect 32539 11132 32551 11135
rect 32769 11135 32827 11141
rect 32769 11132 32781 11135
rect 32539 11104 32781 11132
rect 32539 11101 32551 11104
rect 32493 11095 32551 11101
rect 32769 11101 32781 11104
rect 32815 11132 32827 11135
rect 32968 11132 32996 11160
rect 32815 11104 32996 11132
rect 33045 11135 33103 11141
rect 32815 11101 32827 11104
rect 32769 11095 32827 11101
rect 33045 11101 33057 11135
rect 33091 11101 33103 11135
rect 33045 11095 33103 11101
rect 28261 11067 28319 11073
rect 28261 11033 28273 11067
rect 28307 11064 28319 11067
rect 31404 11064 31432 11092
rect 33060 11064 33088 11095
rect 33134 11092 33140 11144
rect 33192 11132 33198 11144
rect 33229 11135 33287 11141
rect 33229 11132 33241 11135
rect 33192 11104 33241 11132
rect 33192 11092 33198 11104
rect 33229 11101 33241 11104
rect 33275 11101 33287 11135
rect 33229 11095 33287 11101
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 37553 11135 37611 11141
rect 37553 11132 37565 11135
rect 37332 11104 37565 11132
rect 37332 11092 37338 11104
rect 37553 11101 37565 11104
rect 37599 11101 37611 11135
rect 37553 11095 37611 11101
rect 28307 11036 31432 11064
rect 32600 11036 33088 11064
rect 28307 11033 28319 11036
rect 28261 11027 28319 11033
rect 32600 11008 32628 11036
rect 37918 11024 37924 11076
rect 37976 11024 37982 11076
rect 29822 10996 29828 11008
rect 27764 10968 29828 10996
rect 27764 10956 27770 10968
rect 29822 10956 29828 10968
rect 29880 10956 29886 11008
rect 32582 10956 32588 11008
rect 32640 10956 32646 11008
rect 1104 10906 38272 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38272 10906
rect 1104 10832 38272 10854
rect 3234 10752 3240 10804
rect 3292 10752 3298 10804
rect 4614 10752 4620 10804
rect 4672 10752 4678 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 5077 10795 5135 10801
rect 5077 10792 5089 10795
rect 4764 10764 5089 10792
rect 4764 10752 4770 10764
rect 5077 10761 5089 10764
rect 5123 10761 5135 10795
rect 5077 10755 5135 10761
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10100 10764 10456 10792
rect 10100 10752 10106 10764
rect 3053 10727 3111 10733
rect 3053 10693 3065 10727
rect 3099 10724 3111 10727
rect 3252 10724 3280 10752
rect 6089 10727 6147 10733
rect 3099 10696 3280 10724
rect 5000 10696 6040 10724
rect 3099 10693 3111 10696
rect 3053 10687 3111 10693
rect 5000 10665 5028 10696
rect 4985 10659 5043 10665
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 2777 10591 2835 10597
rect 2777 10588 2789 10591
rect 1452 10560 2789 10588
rect 1452 10548 1458 10560
rect 2777 10557 2789 10560
rect 2823 10557 2835 10591
rect 2777 10551 2835 10557
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 4172 10452 4200 10642
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5074 10616 5080 10668
rect 5132 10656 5138 10668
rect 5442 10656 5448 10668
rect 5132 10628 5448 10656
rect 5132 10616 5138 10628
rect 5442 10616 5448 10628
rect 5500 10656 5506 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5500 10628 5733 10656
rect 5500 10616 5506 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 6012 10656 6040 10696
rect 6089 10693 6101 10727
rect 6135 10724 6147 10727
rect 6135 10696 10364 10724
rect 6135 10693 6147 10696
rect 6089 10687 6147 10693
rect 6012 10628 6500 10656
rect 5905 10619 5963 10625
rect 4430 10548 4436 10600
rect 4488 10588 4494 10600
rect 5092 10588 5120 10616
rect 4488 10560 5120 10588
rect 4488 10548 4494 10560
rect 5166 10548 5172 10600
rect 5224 10548 5230 10600
rect 4525 10523 4583 10529
rect 4525 10489 4537 10523
rect 4571 10520 4583 10523
rect 4890 10520 4896 10532
rect 4571 10492 4896 10520
rect 4571 10489 4583 10492
rect 4525 10483 4583 10489
rect 4890 10480 4896 10492
rect 4948 10520 4954 10532
rect 5920 10520 5948 10619
rect 6086 10548 6092 10600
rect 6144 10548 6150 10600
rect 6472 10588 6500 10628
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 9766 10656 9772 10668
rect 7892 10628 9772 10656
rect 7892 10616 7898 10628
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 6472 10560 9260 10588
rect 4948 10492 5948 10520
rect 6104 10520 6132 10548
rect 9122 10520 9128 10532
rect 6104 10492 9128 10520
rect 4948 10480 4954 10492
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 9232 10520 9260 10560
rect 10134 10548 10140 10600
rect 10192 10588 10198 10600
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 10192 10560 10241 10588
rect 10192 10548 10198 10560
rect 10229 10557 10241 10560
rect 10275 10557 10287 10591
rect 10336 10588 10364 10696
rect 10428 10665 10456 10764
rect 11790 10752 11796 10804
rect 11848 10752 11854 10804
rect 11974 10752 11980 10804
rect 12032 10752 12038 10804
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 14148 10764 14289 10792
rect 14148 10752 14154 10764
rect 14277 10761 14289 10764
rect 14323 10761 14335 10795
rect 15654 10792 15660 10804
rect 14277 10755 14335 10761
rect 15304 10764 15660 10792
rect 11992 10665 12020 10752
rect 13538 10684 13544 10736
rect 13596 10724 13602 10736
rect 14918 10724 14924 10736
rect 13596 10696 14924 10724
rect 13596 10684 13602 10696
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 15013 10727 15071 10733
rect 15013 10693 15025 10727
rect 15059 10724 15071 10727
rect 15304 10724 15332 10764
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 20162 10792 20168 10804
rect 20088 10764 20168 10792
rect 15059 10696 15332 10724
rect 15059 10693 15071 10696
rect 15013 10687 15071 10693
rect 15562 10684 15568 10736
rect 15620 10684 15626 10736
rect 17586 10684 17592 10736
rect 17644 10684 17650 10736
rect 19426 10684 19432 10736
rect 19484 10684 19490 10736
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 12124 10628 13461 10656
rect 12124 10616 12130 10628
rect 13449 10625 13461 10628
rect 13495 10656 13507 10659
rect 13495 10628 14596 10656
rect 13495 10625 13507 10628
rect 13449 10619 13507 10625
rect 10336 10560 13492 10588
rect 10229 10551 10287 10557
rect 13081 10523 13139 10529
rect 13081 10520 13093 10523
rect 9232 10492 13093 10520
rect 13081 10489 13093 10492
rect 13127 10489 13139 10523
rect 13464 10520 13492 10560
rect 13722 10548 13728 10600
rect 13780 10548 13786 10600
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 14366 10588 14372 10600
rect 14364 10548 14372 10588
rect 14424 10548 14430 10600
rect 14458 10548 14464 10600
rect 14516 10548 14522 10600
rect 14568 10588 14596 10628
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14700 10628 14749 10656
rect 14700 10616 14706 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 14737 10619 14795 10625
rect 16500 10628 16865 10656
rect 16500 10597 16528 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 18046 10616 18052 10668
rect 18104 10616 18110 10668
rect 18506 10616 18512 10668
rect 18564 10656 18570 10668
rect 18693 10659 18751 10665
rect 18693 10656 18705 10659
rect 18564 10628 18705 10656
rect 18564 10616 18570 10628
rect 18693 10625 18705 10628
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 16485 10591 16543 10597
rect 14568 10560 16068 10588
rect 13924 10520 13952 10548
rect 13464 10492 13952 10520
rect 14364 10520 14392 10548
rect 16040 10520 16068 10560
rect 16485 10557 16497 10591
rect 16531 10557 16543 10591
rect 19444 10588 19472 10684
rect 20088 10665 20116 10764
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 21266 10792 21272 10804
rect 20680 10764 21272 10792
rect 20680 10752 20686 10764
rect 21266 10752 21272 10764
rect 21324 10792 21330 10804
rect 21361 10795 21419 10801
rect 21361 10792 21373 10795
rect 21324 10764 21373 10792
rect 21324 10752 21330 10764
rect 21361 10761 21373 10764
rect 21407 10792 21419 10795
rect 22833 10795 22891 10801
rect 22833 10792 22845 10795
rect 21407 10764 22845 10792
rect 21407 10761 21419 10764
rect 21361 10755 21419 10761
rect 22833 10761 22845 10764
rect 22879 10761 22891 10795
rect 22833 10755 22891 10761
rect 23566 10752 23572 10804
rect 23624 10752 23630 10804
rect 25866 10752 25872 10804
rect 25924 10752 25930 10804
rect 26602 10752 26608 10804
rect 26660 10752 26666 10804
rect 30558 10752 30564 10804
rect 30616 10792 30622 10804
rect 30616 10764 33088 10792
rect 30616 10752 30622 10764
rect 21910 10724 21916 10736
rect 20180 10696 20944 10724
rect 20180 10665 20208 10696
rect 20916 10668 20944 10696
rect 21116 10696 21916 10724
rect 20073 10659 20131 10665
rect 20073 10625 20085 10659
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 20165 10659 20223 10665
rect 20165 10625 20177 10659
rect 20211 10625 20223 10659
rect 20165 10619 20223 10625
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 20272 10588 20300 10619
rect 20438 10616 20444 10668
rect 20496 10656 20502 10668
rect 20496 10628 20857 10656
rect 20496 10616 20502 10628
rect 20530 10588 20536 10600
rect 19444 10560 20536 10588
rect 16485 10551 16543 10557
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 20829 10588 20857 10628
rect 20898 10616 20904 10668
rect 20956 10616 20962 10668
rect 21116 10588 21144 10696
rect 21468 10665 21496 10696
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 22005 10727 22063 10733
rect 22005 10693 22017 10727
rect 22051 10724 22063 10727
rect 23382 10724 23388 10736
rect 22051 10696 23388 10724
rect 22051 10693 22063 10696
rect 22005 10687 22063 10693
rect 23382 10684 23388 10696
rect 23440 10684 23446 10736
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10625 21235 10659
rect 21177 10619 21235 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 21453 10619 21511 10625
rect 20829 10560 21144 10588
rect 21192 10588 21220 10619
rect 21818 10616 21824 10668
rect 21876 10616 21882 10668
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 22235 10628 22477 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22465 10625 22477 10628
rect 22511 10625 22523 10659
rect 22465 10619 22523 10625
rect 21542 10588 21548 10600
rect 21192 10560 21548 10588
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 19061 10523 19119 10529
rect 14364 10492 14780 10520
rect 16040 10492 18828 10520
rect 13081 10483 13139 10489
rect 5350 10452 5356 10464
rect 3844 10424 5356 10452
rect 3844 10412 3850 10424
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 8754 10412 8760 10464
rect 8812 10452 8818 10464
rect 10134 10452 10140 10464
rect 8812 10424 10140 10452
rect 8812 10412 8818 10424
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 13909 10455 13967 10461
rect 13909 10421 13921 10455
rect 13955 10452 13967 10455
rect 14642 10452 14648 10464
rect 13955 10424 14648 10452
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 14752 10452 14780 10492
rect 18800 10464 18828 10492
rect 19061 10489 19073 10523
rect 19107 10520 19119 10523
rect 19150 10520 19156 10532
rect 19107 10492 19156 10520
rect 19107 10489 19119 10492
rect 19061 10483 19119 10489
rect 19150 10480 19156 10492
rect 19208 10520 19214 10532
rect 20254 10520 20260 10532
rect 19208 10492 20260 10520
rect 19208 10480 19214 10492
rect 20254 10480 20260 10492
rect 20312 10480 20318 10532
rect 20441 10523 20499 10529
rect 20441 10489 20453 10523
rect 20487 10520 20499 10523
rect 20806 10520 20812 10532
rect 20487 10492 20812 10520
rect 20487 10489 20499 10492
rect 20441 10483 20499 10489
rect 20806 10480 20812 10492
rect 20864 10520 20870 10532
rect 22112 10520 22140 10619
rect 22554 10616 22560 10668
rect 22612 10656 22618 10668
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 22612 10628 22661 10656
rect 22612 10616 22618 10628
rect 22649 10625 22661 10628
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 22925 10659 22983 10665
rect 22925 10625 22937 10659
rect 22971 10656 22983 10659
rect 23106 10656 23112 10668
rect 22971 10628 23112 10656
rect 22971 10625 22983 10628
rect 22925 10619 22983 10625
rect 23106 10616 23112 10628
rect 23164 10616 23170 10668
rect 23290 10616 23296 10668
rect 23348 10656 23354 10668
rect 23584 10665 23612 10752
rect 23477 10659 23535 10665
rect 23477 10656 23489 10659
rect 23348 10628 23489 10656
rect 23348 10616 23354 10628
rect 23477 10625 23489 10628
rect 23523 10625 23535 10659
rect 23477 10619 23535 10625
rect 23569 10659 23627 10665
rect 23569 10625 23581 10659
rect 23615 10625 23627 10659
rect 25884 10656 25912 10752
rect 26620 10724 26648 10752
rect 26620 10696 27384 10724
rect 27356 10668 27384 10696
rect 28460 10696 29132 10724
rect 28460 10668 28488 10696
rect 26973 10659 27031 10665
rect 26973 10656 26985 10659
rect 25884 10628 26985 10656
rect 23569 10619 23627 10625
rect 26973 10625 26985 10628
rect 27019 10625 27031 10659
rect 26973 10619 27031 10625
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 25222 10588 25228 10600
rect 23584 10560 25228 10588
rect 23584 10532 23612 10560
rect 25222 10548 25228 10560
rect 25280 10548 25286 10600
rect 26418 10548 26424 10600
rect 26476 10588 26482 10600
rect 27172 10588 27200 10619
rect 27338 10616 27344 10668
rect 27396 10616 27402 10668
rect 27522 10616 27528 10668
rect 27580 10616 27586 10668
rect 28442 10616 28448 10668
rect 28500 10616 28506 10668
rect 28534 10616 28540 10668
rect 28592 10616 28598 10668
rect 28644 10665 28672 10696
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10625 28687 10659
rect 28629 10619 28687 10625
rect 28718 10616 28724 10668
rect 28776 10656 28782 10668
rect 29104 10665 29132 10696
rect 28905 10659 28963 10665
rect 28905 10656 28917 10659
rect 28776 10628 28917 10656
rect 28776 10616 28782 10628
rect 28905 10625 28917 10628
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 29089 10659 29147 10665
rect 29089 10625 29101 10659
rect 29135 10625 29147 10659
rect 29089 10619 29147 10625
rect 26476 10560 27200 10588
rect 26476 10548 26482 10560
rect 27246 10548 27252 10600
rect 27304 10548 27310 10600
rect 28920 10588 28948 10619
rect 30466 10616 30472 10668
rect 30524 10656 30530 10668
rect 30742 10656 30748 10668
rect 30524 10628 30748 10656
rect 30524 10616 30530 10628
rect 30742 10616 30748 10628
rect 30800 10616 30806 10668
rect 30929 10659 30987 10665
rect 30929 10625 30941 10659
rect 30975 10656 30987 10659
rect 31938 10656 31944 10668
rect 30975 10628 31944 10656
rect 30975 10625 30987 10628
rect 30929 10619 30987 10625
rect 31938 10616 31944 10628
rect 31996 10656 32002 10668
rect 32306 10656 32312 10668
rect 31996 10628 32312 10656
rect 31996 10616 32002 10628
rect 32306 10616 32312 10628
rect 32364 10616 32370 10668
rect 32490 10616 32496 10668
rect 32548 10656 32554 10668
rect 32677 10659 32735 10665
rect 32677 10656 32689 10659
rect 32548 10628 32689 10656
rect 32548 10616 32554 10628
rect 32677 10625 32689 10628
rect 32723 10625 32735 10659
rect 33060 10656 33088 10764
rect 34882 10752 34888 10804
rect 34940 10752 34946 10804
rect 33870 10724 33876 10736
rect 33244 10696 33876 10724
rect 33137 10659 33195 10665
rect 33137 10656 33149 10659
rect 33060 10628 33149 10656
rect 32677 10619 32735 10625
rect 33137 10625 33149 10628
rect 33183 10656 33195 10659
rect 33244 10656 33272 10696
rect 33870 10684 33876 10696
rect 33928 10684 33934 10736
rect 33183 10628 33272 10656
rect 33183 10625 33195 10628
rect 33137 10619 33195 10625
rect 33686 10616 33692 10668
rect 33744 10656 33750 10668
rect 34517 10659 34575 10665
rect 34517 10656 34529 10659
rect 33744 10628 34529 10656
rect 33744 10616 33750 10628
rect 34517 10625 34529 10628
rect 34563 10625 34575 10659
rect 34517 10619 34575 10625
rect 36538 10616 36544 10668
rect 36596 10616 36602 10668
rect 36630 10616 36636 10668
rect 36688 10656 36694 10668
rect 36725 10659 36783 10665
rect 36725 10656 36737 10659
rect 36688 10628 36737 10656
rect 36688 10616 36694 10628
rect 36725 10625 36737 10628
rect 36771 10625 36783 10659
rect 36725 10619 36783 10625
rect 30650 10588 30656 10600
rect 27356 10560 30656 10588
rect 20864 10492 22140 10520
rect 20864 10480 20870 10492
rect 23566 10480 23572 10532
rect 23624 10480 23630 10532
rect 24854 10480 24860 10532
rect 24912 10520 24918 10532
rect 27356 10520 27384 10560
rect 30650 10548 30656 10560
rect 30708 10548 30714 10600
rect 30837 10591 30895 10597
rect 30837 10557 30849 10591
rect 30883 10588 30895 10591
rect 32582 10588 32588 10600
rect 30883 10560 32588 10588
rect 30883 10557 30895 10560
rect 30837 10551 30895 10557
rect 32582 10548 32588 10560
rect 32640 10548 32646 10600
rect 34606 10548 34612 10600
rect 34664 10548 34670 10600
rect 24912 10492 27384 10520
rect 24912 10480 24918 10492
rect 28626 10480 28632 10532
rect 28684 10520 28690 10532
rect 28721 10523 28779 10529
rect 28721 10520 28733 10523
rect 28684 10492 28733 10520
rect 28684 10480 28690 10492
rect 28721 10489 28733 10492
rect 28767 10489 28779 10523
rect 28721 10483 28779 10489
rect 29181 10523 29239 10529
rect 29181 10489 29193 10523
rect 29227 10489 29239 10523
rect 33045 10523 33103 10529
rect 33045 10520 33057 10523
rect 29181 10483 29239 10489
rect 30484 10492 33057 10520
rect 17310 10452 17316 10464
rect 14752 10424 17316 10452
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18414 10452 18420 10464
rect 17920 10424 18420 10452
rect 17920 10412 17926 10424
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18782 10412 18788 10464
rect 18840 10412 18846 10464
rect 21177 10455 21235 10461
rect 21177 10421 21189 10455
rect 21223 10452 21235 10455
rect 21634 10452 21640 10464
rect 21223 10424 21640 10452
rect 21223 10421 21235 10424
rect 21177 10415 21235 10421
rect 21634 10412 21640 10424
rect 21692 10412 21698 10464
rect 22370 10412 22376 10464
rect 22428 10412 22434 10464
rect 23750 10412 23756 10464
rect 23808 10412 23814 10464
rect 24210 10412 24216 10464
rect 24268 10452 24274 10464
rect 26878 10452 26884 10464
rect 24268 10424 26884 10452
rect 24268 10412 24274 10424
rect 26878 10412 26884 10424
rect 26936 10412 26942 10464
rect 27706 10412 27712 10464
rect 27764 10412 27770 10464
rect 29196 10452 29224 10483
rect 30484 10464 30512 10492
rect 33045 10489 33057 10492
rect 33091 10520 33103 10523
rect 33870 10520 33876 10532
rect 33091 10492 33876 10520
rect 33091 10489 33103 10492
rect 33045 10483 33103 10489
rect 33870 10480 33876 10492
rect 33928 10480 33934 10532
rect 29362 10452 29368 10464
rect 29196 10424 29368 10452
rect 29362 10412 29368 10424
rect 29420 10452 29426 10464
rect 29638 10452 29644 10464
rect 29420 10424 29644 10452
rect 29420 10412 29426 10424
rect 29638 10412 29644 10424
rect 29696 10412 29702 10464
rect 30466 10412 30472 10464
rect 30524 10412 30530 10464
rect 32490 10412 32496 10464
rect 32548 10452 32554 10464
rect 33134 10452 33140 10464
rect 32548 10424 33140 10452
rect 32548 10412 32554 10424
rect 33134 10412 33140 10424
rect 33192 10452 33198 10464
rect 33229 10455 33287 10461
rect 33229 10452 33241 10455
rect 33192 10424 33241 10452
rect 33192 10412 33198 10424
rect 33229 10421 33241 10424
rect 33275 10421 33287 10455
rect 33229 10415 33287 10421
rect 36906 10412 36912 10464
rect 36964 10412 36970 10464
rect 1104 10362 38272 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38272 10362
rect 1104 10288 38272 10310
rect 4614 10208 4620 10260
rect 4672 10208 4678 10260
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 4798 10248 4804 10260
rect 4755 10220 4804 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5984 10251 6042 10257
rect 5984 10217 5996 10251
rect 6030 10248 6042 10251
rect 6362 10248 6368 10260
rect 6030 10220 6368 10248
rect 6030 10217 6042 10220
rect 5984 10211 6042 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8662 10248 8668 10260
rect 8067 10220 8668 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 9398 10208 9404 10260
rect 9456 10208 9462 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9548 10220 12434 10248
rect 9548 10208 9554 10220
rect 2866 10140 2872 10192
rect 2924 10180 2930 10192
rect 3234 10180 3240 10192
rect 2924 10152 3240 10180
rect 2924 10140 2930 10152
rect 3234 10140 3240 10152
rect 3292 10140 3298 10192
rect 8570 10180 8576 10192
rect 7944 10152 8576 10180
rect 4249 10115 4307 10121
rect 2884 10084 3372 10112
rect 2884 10056 2912 10084
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 2792 9976 2820 10007
rect 2866 10004 2872 10056
rect 2924 10004 2930 10056
rect 2958 10004 2964 10056
rect 3016 10004 3022 10056
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3234 10044 3240 10056
rect 3191 10016 3240 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3344 10044 3372 10084
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 5721 10115 5779 10121
rect 4295 10084 4936 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 4908 10056 4936 10084
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 6086 10112 6092 10124
rect 5767 10084 6092 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 7650 10112 7656 10124
rect 6420 10084 7656 10112
rect 6420 10072 6426 10084
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7944 10112 7972 10152
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 7852 10084 7972 10112
rect 8113 10115 8171 10121
rect 4338 10044 4344 10056
rect 3344 10016 4344 10044
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4706 10044 4712 10056
rect 4479 10016 4712 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4890 10004 4896 10056
rect 4948 10004 4954 10056
rect 7852 10053 7880 10084
rect 8113 10081 8125 10115
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 7926 10004 7932 10056
rect 7984 10004 7990 10056
rect 6270 9976 6276 9988
rect 2792 9948 6276 9976
rect 6270 9936 6276 9948
rect 6328 9936 6334 9988
rect 7374 9976 7380 9988
rect 7222 9948 7380 9976
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 7745 9979 7803 9985
rect 7745 9945 7757 9979
rect 7791 9945 7803 9979
rect 8128 9976 8156 10075
rect 8386 10072 8392 10124
rect 8444 10072 8450 10124
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8588 10112 8616 10140
rect 8527 10084 8616 10112
rect 8665 10115 8723 10121
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 8665 10081 8677 10115
rect 8711 10112 8723 10115
rect 9030 10112 9036 10124
rect 8711 10084 9036 10112
rect 8711 10081 8723 10084
rect 8665 10075 8723 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 9140 10112 9168 10208
rect 12406 10180 12434 10220
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14240 10220 14504 10248
rect 14240 10208 14246 10220
rect 14093 10183 14151 10189
rect 14093 10180 14105 10183
rect 12406 10152 14105 10180
rect 14093 10149 14105 10152
rect 14139 10149 14151 10183
rect 14093 10143 14151 10149
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 9140 10084 10333 10112
rect 10321 10081 10333 10084
rect 10367 10112 10379 10115
rect 11054 10112 11060 10124
rect 10367 10084 11060 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8754 10044 8760 10056
rect 8619 10016 8760 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10044 8999 10047
rect 9122 10044 9128 10056
rect 8987 10016 9128 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 7745 9939 7803 9945
rect 7944 9948 8156 9976
rect 1486 9868 1492 9920
rect 1544 9908 1550 9920
rect 2501 9911 2559 9917
rect 2501 9908 2513 9911
rect 1544 9880 2513 9908
rect 1544 9868 1550 9880
rect 2501 9877 2513 9880
rect 2547 9877 2559 9911
rect 2501 9871 2559 9877
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7760 9908 7788 9939
rect 7944 9920 7972 9948
rect 8846 9936 8852 9988
rect 8904 9976 8910 9988
rect 9030 9976 9036 9988
rect 8904 9948 9036 9976
rect 8904 9936 8910 9948
rect 9030 9936 9036 9948
rect 9088 9976 9094 9988
rect 9232 9976 9260 10007
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 9401 10047 9459 10053
rect 9401 10044 9413 10047
rect 9364 10016 9413 10044
rect 9364 10004 9370 10016
rect 9401 10013 9413 10016
rect 9447 10044 9459 10047
rect 9582 10044 9588 10056
rect 9447 10016 9588 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 10597 9979 10655 9985
rect 10597 9976 10609 9979
rect 9088 9948 9260 9976
rect 10060 9948 10609 9976
rect 9088 9936 9094 9948
rect 6972 9880 7788 9908
rect 6972 9868 6978 9880
rect 7926 9868 7932 9920
rect 7984 9868 7990 9920
rect 8110 9868 8116 9920
rect 8168 9908 8174 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 8168 9880 8217 9908
rect 8168 9868 8174 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 10060 9917 10088 9948
rect 10597 9945 10609 9948
rect 10643 9945 10655 9979
rect 11822 9948 12434 9976
rect 10597 9939 10655 9945
rect 9585 9911 9643 9917
rect 9585 9908 9597 9911
rect 8628 9880 9597 9908
rect 8628 9868 8634 9880
rect 9585 9877 9597 9880
rect 9631 9877 9643 9911
rect 9585 9871 9643 9877
rect 10045 9911 10103 9917
rect 10045 9877 10057 9911
rect 10091 9877 10103 9911
rect 10045 9871 10103 9877
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 11900 9908 11928 9948
rect 11020 9880 11928 9908
rect 11020 9868 11026 9880
rect 12066 9868 12072 9920
rect 12124 9868 12130 9920
rect 12406 9908 12434 9948
rect 12802 9908 12808 9920
rect 12406 9880 12808 9908
rect 12802 9868 12808 9880
rect 12860 9908 12866 9920
rect 13538 9908 13544 9920
rect 12860 9880 13544 9908
rect 12860 9868 12866 9880
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 14292 9908 14320 10007
rect 14366 10004 14372 10056
rect 14424 10004 14430 10056
rect 14476 10044 14504 10220
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 16945 10251 17003 10257
rect 14976 10220 16804 10248
rect 14976 10208 14982 10220
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 15197 10115 15255 10121
rect 15197 10112 15209 10115
rect 14792 10084 15209 10112
rect 14792 10072 14798 10084
rect 15197 10081 15209 10084
rect 15243 10081 15255 10115
rect 15197 10075 15255 10081
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 16666 10112 16672 10124
rect 15620 10084 16672 10112
rect 15620 10072 15626 10084
rect 16666 10072 16672 10084
rect 16724 10072 16730 10124
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14476 10016 14565 10044
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 14642 10004 14648 10056
rect 14700 10044 14706 10056
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 14700 10016 15025 10044
rect 14700 10004 14706 10016
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 16776 10044 16804 10220
rect 16945 10217 16957 10251
rect 16991 10248 17003 10251
rect 17310 10248 17316 10260
rect 16991 10220 17316 10248
rect 16991 10217 17003 10220
rect 16945 10211 17003 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 24486 10248 24492 10260
rect 17420 10220 19012 10248
rect 17420 10121 17448 10220
rect 17512 10152 18920 10180
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 17512 10044 17540 10152
rect 17862 10072 17868 10124
rect 17920 10072 17926 10124
rect 18506 10112 18512 10124
rect 18156 10084 18512 10112
rect 16776 10016 17540 10044
rect 17773 10047 17831 10053
rect 15013 10007 15071 10013
rect 17773 10013 17785 10047
rect 17819 10044 17831 10047
rect 17954 10044 17960 10056
rect 17819 10016 17960 10044
rect 17819 10013 17831 10016
rect 17773 10007 17831 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18156 10053 18184 10084
rect 18506 10072 18512 10084
rect 18564 10112 18570 10124
rect 18564 10084 18736 10112
rect 18564 10072 18570 10084
rect 18141 10047 18199 10053
rect 18141 10013 18153 10047
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18230 10004 18236 10056
rect 18288 10044 18294 10056
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 18288 10016 18337 10044
rect 18288 10004 18294 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 14384 9976 14412 10004
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 14384 9948 14473 9976
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 14461 9939 14519 9945
rect 15473 9979 15531 9985
rect 15473 9945 15485 9979
rect 15519 9945 15531 9979
rect 15473 9939 15531 9945
rect 14734 9908 14740 9920
rect 14292 9880 14740 9908
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 14829 9911 14887 9917
rect 14829 9877 14841 9911
rect 14875 9908 14887 9911
rect 15488 9908 15516 9939
rect 15562 9936 15568 9988
rect 15620 9976 15626 9988
rect 17972 9976 18000 10004
rect 18432 9976 18460 10007
rect 18598 10004 18604 10056
rect 18656 10004 18662 10056
rect 18708 10053 18736 10084
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10013 18751 10047
rect 18693 10007 18751 10013
rect 18782 10004 18788 10056
rect 18840 10004 18846 10056
rect 18892 10044 18920 10152
rect 18984 10112 19012 10220
rect 19076 10220 24492 10248
rect 19076 10189 19104 10220
rect 24486 10208 24492 10220
rect 24544 10208 24550 10260
rect 24596 10220 31432 10248
rect 19061 10183 19119 10189
rect 19061 10149 19073 10183
rect 19107 10149 19119 10183
rect 20254 10180 20260 10192
rect 19061 10143 19119 10149
rect 19168 10152 20260 10180
rect 19168 10112 19196 10152
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 20806 10140 20812 10192
rect 20864 10140 20870 10192
rect 21082 10140 21088 10192
rect 21140 10140 21146 10192
rect 21300 10152 21496 10180
rect 18984 10084 19196 10112
rect 19242 10072 19248 10124
rect 19300 10072 19306 10124
rect 20622 10072 20628 10124
rect 20680 10072 20686 10124
rect 19429 10047 19487 10053
rect 19429 10044 19441 10047
rect 18892 10016 19441 10044
rect 19429 10013 19441 10016
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 20073 10047 20131 10053
rect 20073 10044 20085 10047
rect 19944 10016 20085 10044
rect 19944 10004 19950 10016
rect 20073 10013 20085 10016
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 20349 10047 20407 10053
rect 20349 10013 20361 10047
rect 20395 10044 20407 10047
rect 20438 10044 20444 10056
rect 20395 10016 20444 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 20824 10053 20852 10140
rect 21300 10112 21328 10152
rect 20916 10084 21328 10112
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 20809 10047 20867 10053
rect 20809 10013 20821 10047
rect 20855 10013 20867 10047
rect 20809 10007 20867 10013
rect 20548 9976 20576 10007
rect 15620 9948 15962 9976
rect 17972 9948 18460 9976
rect 20272 9948 20576 9976
rect 15620 9936 15626 9948
rect 20272 9920 20300 9948
rect 14875 9880 15516 9908
rect 14875 9877 14887 9880
rect 14829 9871 14887 9877
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 18230 9908 18236 9920
rect 16172 9880 18236 9908
rect 16172 9868 16178 9880
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19484 9880 19625 9908
rect 19484 9868 19490 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 20165 9911 20223 9917
rect 20165 9877 20177 9911
rect 20211 9908 20223 9911
rect 20254 9908 20260 9920
rect 20211 9880 20260 9908
rect 20211 9877 20223 9880
rect 20165 9871 20223 9877
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 20441 9911 20499 9917
rect 20441 9877 20453 9911
rect 20487 9908 20499 9911
rect 20916 9908 20944 10084
rect 21358 10072 21364 10124
rect 21416 10072 21422 10124
rect 21468 10121 21496 10152
rect 22186 10140 22192 10192
rect 22244 10140 22250 10192
rect 22646 10180 22652 10192
rect 22296 10152 22652 10180
rect 21453 10115 21511 10121
rect 21453 10081 21465 10115
rect 21499 10081 21511 10115
rect 21453 10075 21511 10081
rect 21545 10115 21603 10121
rect 21545 10081 21557 10115
rect 21591 10112 21603 10115
rect 21634 10112 21640 10124
rect 21591 10084 21640 10112
rect 21591 10081 21603 10084
rect 21545 10075 21603 10081
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 22296 10112 22324 10152
rect 22646 10140 22652 10152
rect 22704 10140 22710 10192
rect 24397 10183 24455 10189
rect 24397 10149 24409 10183
rect 24443 10180 24455 10183
rect 24596 10180 24624 10220
rect 24443 10152 24624 10180
rect 24443 10149 24455 10152
rect 24397 10143 24455 10149
rect 27706 10140 27712 10192
rect 27764 10140 27770 10192
rect 29914 10180 29920 10192
rect 29656 10152 29920 10180
rect 24857 10115 24915 10121
rect 24857 10112 24869 10115
rect 21744 10084 22324 10112
rect 22388 10084 24869 10112
rect 21744 10053 21772 10084
rect 22388 10053 22416 10084
rect 24857 10081 24869 10084
rect 24903 10081 24915 10115
rect 24857 10075 24915 10081
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10081 25007 10115
rect 27724 10112 27752 10140
rect 24949 10075 25007 10081
rect 27172 10084 27752 10112
rect 29012 10084 29408 10112
rect 21269 10047 21327 10053
rect 21269 10013 21281 10047
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10013 21787 10047
rect 22373 10047 22431 10053
rect 22373 10044 22385 10047
rect 21729 10007 21787 10013
rect 21836 10016 22385 10044
rect 20993 9979 21051 9985
rect 20993 9945 21005 9979
rect 21039 9976 21051 9979
rect 21284 9976 21312 10007
rect 21836 9976 21864 10016
rect 22373 10013 22385 10016
rect 22419 10013 22431 10047
rect 22373 10007 22431 10013
rect 22462 10004 22468 10056
rect 22520 10004 22526 10056
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 21039 9948 21864 9976
rect 21039 9945 21051 9948
rect 20993 9939 21051 9945
rect 21910 9936 21916 9988
rect 21968 9976 21974 9988
rect 22664 9976 22692 10007
rect 22738 10004 22744 10056
rect 22796 10004 22802 10056
rect 23014 10004 23020 10056
rect 23072 10004 23078 10056
rect 23106 10004 23112 10056
rect 23164 10004 23170 10056
rect 23198 10004 23204 10056
rect 23256 10004 23262 10056
rect 23474 10004 23480 10056
rect 23532 10004 23538 10056
rect 23750 10004 23756 10056
rect 23808 10004 23814 10056
rect 24118 10004 24124 10056
rect 24176 10044 24182 10056
rect 24578 10044 24584 10056
rect 24176 10016 24584 10044
rect 24176 10004 24182 10016
rect 24578 10004 24584 10016
rect 24636 10044 24642 10056
rect 24964 10044 24992 10075
rect 24636 10016 24992 10044
rect 24636 10004 24642 10016
rect 26234 10004 26240 10056
rect 26292 10004 26298 10056
rect 26970 10004 26976 10056
rect 27028 10004 27034 10056
rect 27062 10004 27068 10056
rect 27120 10004 27126 10056
rect 27172 10053 27200 10084
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10013 27215 10047
rect 27157 10007 27215 10013
rect 27341 10047 27399 10053
rect 27341 10013 27353 10047
rect 27387 10013 27399 10047
rect 27341 10007 27399 10013
rect 23216 9976 23244 10004
rect 21968 9948 22692 9976
rect 22756 9948 23244 9976
rect 23339 9979 23397 9985
rect 21968 9936 21974 9948
rect 20487 9880 20944 9908
rect 20487 9877 20499 9880
rect 20441 9871 20499 9877
rect 22278 9868 22284 9920
rect 22336 9908 22342 9920
rect 22756 9908 22784 9948
rect 23339 9945 23351 9979
rect 23385 9976 23397 9979
rect 23768 9976 23796 10004
rect 23385 9948 23796 9976
rect 23385 9945 23397 9948
rect 23339 9939 23397 9945
rect 24486 9936 24492 9988
rect 24544 9976 24550 9988
rect 26252 9976 26280 10004
rect 27356 9976 27384 10007
rect 28442 10004 28448 10056
rect 28500 10044 28506 10056
rect 28537 10047 28595 10053
rect 28537 10044 28549 10047
rect 28500 10016 28549 10044
rect 28500 10004 28506 10016
rect 28537 10013 28549 10016
rect 28583 10013 28595 10047
rect 28537 10007 28595 10013
rect 28718 10004 28724 10056
rect 28776 10004 28782 10056
rect 29012 10053 29040 10084
rect 29380 10056 29408 10084
rect 29656 10063 29684 10152
rect 29914 10140 29920 10152
rect 29972 10140 29978 10192
rect 30466 10180 30472 10192
rect 30392 10152 30472 10180
rect 29641 10057 29699 10063
rect 28997 10047 29055 10053
rect 28997 10013 29009 10047
rect 29043 10013 29055 10047
rect 28997 10007 29055 10013
rect 29086 10004 29092 10056
rect 29144 10044 29150 10056
rect 29181 10047 29239 10053
rect 29181 10044 29193 10047
rect 29144 10016 29193 10044
rect 29144 10004 29150 10016
rect 29181 10013 29193 10016
rect 29227 10013 29239 10047
rect 29181 10007 29239 10013
rect 29362 10004 29368 10056
rect 29420 10004 29426 10056
rect 29641 10023 29653 10057
rect 29687 10023 29699 10057
rect 29641 10017 29699 10023
rect 29822 10004 29828 10056
rect 29880 10004 29886 10056
rect 30392 10053 30420 10152
rect 30466 10140 30472 10152
rect 30524 10140 30530 10192
rect 30650 10140 30656 10192
rect 30708 10180 30714 10192
rect 30708 10152 31340 10180
rect 30708 10140 30714 10152
rect 30834 10112 30840 10124
rect 30576 10084 30840 10112
rect 30193 10047 30251 10053
rect 30193 10013 30205 10047
rect 30239 10013 30251 10047
rect 30193 10007 30251 10013
rect 30377 10047 30435 10053
rect 30377 10013 30389 10047
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 30208 9976 30236 10007
rect 30466 10004 30472 10056
rect 30524 10004 30530 10056
rect 30576 10053 30604 10084
rect 30834 10072 30840 10084
rect 30892 10072 30898 10124
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10013 30619 10047
rect 30561 10007 30619 10013
rect 30650 10004 30656 10056
rect 30708 10044 30714 10056
rect 30745 10047 30803 10053
rect 30745 10044 30757 10047
rect 30708 10016 30757 10044
rect 30708 10004 30714 10016
rect 30745 10013 30757 10016
rect 30791 10013 30803 10047
rect 30745 10007 30803 10013
rect 31205 10047 31263 10053
rect 31205 10013 31217 10047
rect 31251 10013 31263 10047
rect 31205 10007 31263 10013
rect 31220 9976 31248 10007
rect 24544 9948 24900 9976
rect 26252 9948 27384 9976
rect 28828 9948 30236 9976
rect 30300 9948 31248 9976
rect 31312 9976 31340 10152
rect 31404 10112 31432 10220
rect 34606 10208 34612 10260
rect 34664 10248 34670 10260
rect 35161 10251 35219 10257
rect 35161 10248 35173 10251
rect 34664 10220 35173 10248
rect 34664 10208 34670 10220
rect 35161 10217 35173 10220
rect 35207 10217 35219 10251
rect 35161 10211 35219 10217
rect 34241 10183 34299 10189
rect 34241 10149 34253 10183
rect 34287 10180 34299 10183
rect 34287 10152 34928 10180
rect 34287 10149 34299 10152
rect 34241 10143 34299 10149
rect 34793 10115 34851 10121
rect 34793 10112 34805 10115
rect 31404 10084 34805 10112
rect 34793 10081 34805 10084
rect 34839 10081 34851 10115
rect 34793 10075 34851 10081
rect 31573 10047 31631 10053
rect 31573 10013 31585 10047
rect 31619 10044 31631 10047
rect 32490 10044 32496 10056
rect 31619 10016 32496 10044
rect 31619 10013 31631 10016
rect 31573 10007 31631 10013
rect 32490 10004 32496 10016
rect 32548 10004 32554 10056
rect 33781 10047 33839 10053
rect 33781 10044 33793 10047
rect 33244 10016 33793 10044
rect 33244 9976 33272 10016
rect 33781 10013 33793 10016
rect 33827 10013 33839 10047
rect 33781 10007 33839 10013
rect 33870 10004 33876 10056
rect 33928 10004 33934 10056
rect 33962 10004 33968 10056
rect 34020 10004 34026 10056
rect 34054 10004 34060 10056
rect 34112 10044 34118 10056
rect 34900 10053 34928 10152
rect 34149 10047 34207 10053
rect 34149 10044 34161 10047
rect 34112 10016 34161 10044
rect 34112 10004 34118 10016
rect 34149 10013 34161 10016
rect 34195 10013 34207 10047
rect 34517 10047 34575 10053
rect 34517 10044 34529 10047
rect 34149 10007 34207 10013
rect 34348 10016 34529 10044
rect 34348 9988 34376 10016
rect 34517 10013 34529 10016
rect 34563 10013 34575 10047
rect 34517 10007 34575 10013
rect 34885 10047 34943 10053
rect 34885 10013 34897 10047
rect 34931 10013 34943 10047
rect 34885 10007 34943 10013
rect 31312 9948 33272 9976
rect 33505 9979 33563 9985
rect 24544 9936 24550 9948
rect 22336 9880 22784 9908
rect 22336 9868 22342 9880
rect 22830 9868 22836 9920
rect 22888 9868 22894 9920
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 24762 9908 24768 9920
rect 23532 9880 24768 9908
rect 23532 9868 23538 9880
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 24872 9908 24900 9948
rect 26510 9908 26516 9920
rect 24872 9880 26516 9908
rect 26510 9868 26516 9880
rect 26568 9868 26574 9920
rect 26697 9911 26755 9917
rect 26697 9877 26709 9911
rect 26743 9908 26755 9911
rect 28828 9908 28856 9948
rect 26743 9880 28856 9908
rect 26743 9877 26755 9880
rect 26697 9871 26755 9877
rect 28902 9868 28908 9920
rect 28960 9868 28966 9920
rect 29086 9868 29092 9920
rect 29144 9868 29150 9920
rect 29825 9911 29883 9917
rect 29825 9877 29837 9911
rect 29871 9908 29883 9911
rect 30300 9908 30328 9948
rect 33505 9945 33517 9979
rect 33551 9976 33563 9979
rect 34241 9979 34299 9985
rect 34241 9976 34253 9979
rect 33551 9948 34253 9976
rect 33551 9945 33563 9948
rect 33505 9939 33563 9945
rect 34241 9945 34253 9948
rect 34287 9945 34299 9979
rect 34241 9939 34299 9945
rect 34330 9936 34336 9988
rect 34388 9936 34394 9988
rect 29871 9880 30328 9908
rect 29871 9877 29883 9880
rect 29825 9871 29883 9877
rect 30374 9868 30380 9920
rect 30432 9908 30438 9920
rect 30834 9908 30840 9920
rect 30432 9880 30840 9908
rect 30432 9868 30438 9880
rect 30834 9868 30840 9880
rect 30892 9868 30898 9920
rect 30926 9868 30932 9920
rect 30984 9868 30990 9920
rect 32122 9868 32128 9920
rect 32180 9908 32186 9920
rect 32217 9911 32275 9917
rect 32217 9908 32229 9911
rect 32180 9880 32229 9908
rect 32180 9868 32186 9880
rect 32217 9877 32229 9880
rect 32263 9877 32275 9911
rect 32217 9871 32275 9877
rect 33226 9868 33232 9920
rect 33284 9908 33290 9920
rect 34425 9911 34483 9917
rect 34425 9908 34437 9911
rect 33284 9880 34437 9908
rect 33284 9868 33290 9880
rect 34425 9877 34437 9880
rect 34471 9877 34483 9911
rect 34425 9871 34483 9877
rect 1104 9818 38272 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38272 9818
rect 1104 9744 38272 9766
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 6457 9707 6515 9713
rect 4396 9676 5580 9704
rect 4396 9664 4402 9676
rect 3050 9596 3056 9648
rect 3108 9636 3114 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 3108 9608 4537 9636
rect 3108 9596 3114 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 4525 9599 4583 9605
rect 1394 9528 1400 9580
rect 1452 9528 1458 9580
rect 3786 9568 3792 9580
rect 2806 9540 3792 9568
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 4080 9540 4169 9568
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 4080 9376 4108 9540
rect 4157 9537 4169 9540
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4356 9500 4384 9531
rect 4430 9528 4436 9580
rect 4488 9528 4494 9580
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 4908 9577 4936 9676
rect 4781 9571 4839 9577
rect 4781 9568 4793 9571
rect 4724 9540 4793 9568
rect 4632 9500 4660 9528
rect 4356 9472 4660 9500
rect 4724 9500 4752 9540
rect 4781 9537 4793 9540
rect 4827 9537 4839 9571
rect 4781 9531 4839 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5442 9568 5448 9580
rect 5215 9540 5448 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5552 9568 5580 9676
rect 6457 9673 6469 9707
rect 6503 9704 6515 9707
rect 6546 9704 6552 9716
rect 6503 9676 6552 9704
rect 6503 9673 6515 9676
rect 6457 9667 6515 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 7892 9676 9076 9704
rect 7892 9664 7898 9676
rect 6825 9639 6883 9645
rect 6825 9605 6837 9639
rect 6871 9636 6883 9639
rect 7852 9636 7880 9664
rect 6871 9608 7880 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 8570 9636 8576 9648
rect 8260 9608 8432 9636
rect 8260 9596 8266 9608
rect 8294 9568 8300 9580
rect 5552 9540 8300 9568
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 8404 9577 8432 9608
rect 8496 9608 8576 9636
rect 8496 9577 8524 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 8772 9577 8800 9676
rect 9048 9636 9076 9676
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10284 9676 10609 9704
rect 10284 9664 10290 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 10597 9667 10655 9673
rect 11057 9707 11115 9713
rect 11057 9673 11069 9707
rect 11103 9704 11115 9707
rect 12066 9704 12072 9716
rect 11103 9676 12072 9704
rect 11103 9673 11115 9676
rect 11057 9667 11115 9673
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 14274 9704 14280 9716
rect 12492 9676 14280 9704
rect 12492 9664 12498 9676
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 20070 9704 20076 9716
rect 14792 9676 20076 9704
rect 14792 9664 14798 9676
rect 20070 9664 20076 9676
rect 20128 9664 20134 9716
rect 20806 9704 20812 9716
rect 20732 9676 20812 9704
rect 9048 9608 10640 9636
rect 10612 9580 10640 9608
rect 10870 9596 10876 9648
rect 10928 9636 10934 9648
rect 10965 9639 11023 9645
rect 10965 9636 10977 9639
rect 10928 9608 10977 9636
rect 10928 9596 10934 9608
rect 10965 9605 10977 9608
rect 11011 9605 11023 9639
rect 10965 9599 11023 9605
rect 11072 9608 12756 9636
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 8846 9528 8852 9580
rect 8904 9577 8910 9580
rect 8904 9568 8913 9577
rect 9033 9571 9091 9577
rect 8904 9540 8949 9568
rect 8904 9531 8913 9540
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 10226 9568 10232 9580
rect 9079 9540 10232 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 8904 9528 8910 9531
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 11072 9568 11100 9608
rect 10652 9540 11100 9568
rect 12253 9571 12311 9577
rect 10652 9528 10658 9540
rect 12253 9537 12265 9571
rect 12299 9568 12311 9571
rect 12299 9540 12388 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 7101 9503 7159 9509
rect 4724 9472 7052 9500
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 5350 9432 5356 9444
rect 4203 9404 5356 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 7024 9432 7052 9472
rect 7101 9469 7113 9503
rect 7147 9500 7159 9503
rect 7282 9500 7288 9512
rect 7147 9472 7288 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 7282 9460 7288 9472
rect 7340 9500 7346 9512
rect 7834 9500 7840 9512
rect 7340 9472 7840 9500
rect 7340 9460 7346 9472
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 7984 9472 8953 9500
rect 7984 9460 7990 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 10134 9460 10140 9512
rect 10192 9500 10198 9512
rect 11146 9500 11152 9512
rect 10192 9472 11152 9500
rect 10192 9460 10198 9472
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 12360 9441 12388 9540
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 12728 9577 12756 9608
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 19521 9639 19579 9645
rect 19521 9636 19533 9639
rect 19484 9608 19533 9636
rect 19484 9596 19490 9608
rect 19521 9605 19533 9608
rect 19567 9605 19579 9639
rect 20732 9636 20760 9676
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 22278 9704 22284 9716
rect 21100 9676 22284 9704
rect 21100 9648 21128 9676
rect 22278 9664 22284 9676
rect 22336 9664 22342 9716
rect 22370 9664 22376 9716
rect 22428 9664 22434 9716
rect 22738 9664 22744 9716
rect 22796 9704 22802 9716
rect 22925 9707 22983 9713
rect 22925 9704 22937 9707
rect 22796 9676 22937 9704
rect 22796 9664 22802 9676
rect 22925 9673 22937 9676
rect 22971 9673 22983 9707
rect 22925 9667 22983 9673
rect 24486 9664 24492 9716
rect 24544 9674 24550 9716
rect 25041 9707 25099 9713
rect 24544 9664 24588 9674
rect 25041 9673 25053 9707
rect 25087 9673 25099 9707
rect 25041 9667 25099 9673
rect 20732 9608 21036 9636
rect 19521 9599 19579 9605
rect 12713 9571 12771 9577
rect 12713 9537 12725 9571
rect 12759 9568 12771 9571
rect 13078 9568 13084 9580
rect 12759 9540 13084 9568
rect 12759 9537 12771 9540
rect 12713 9531 12771 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9568 14243 9571
rect 14734 9568 14740 9580
rect 14231 9540 14740 9568
rect 14231 9537 14243 9540
rect 14185 9531 14243 9537
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 15252 9540 17877 9568
rect 15252 9528 15258 9540
rect 17865 9537 17877 9540
rect 17911 9568 17923 9571
rect 18506 9568 18512 9580
rect 17911 9540 18512 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9568 20683 9571
rect 20714 9568 20720 9580
rect 20671 9540 20720 9568
rect 20671 9537 20683 9540
rect 20625 9531 20683 9537
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 12636 9500 12664 9528
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12636 9472 12817 9500
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 12894 9460 12900 9512
rect 12952 9460 12958 9512
rect 13814 9500 13820 9512
rect 13004 9472 13820 9500
rect 12345 9435 12403 9441
rect 7024 9404 12204 9432
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 4062 9364 4068 9376
rect 3191 9336 4068 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 4798 9364 4804 9376
rect 4488 9336 4804 9364
rect 4488 9324 4494 9336
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 5166 9364 5172 9376
rect 4948 9336 5172 9364
rect 4948 9324 4954 9336
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 8202 9324 8208 9376
rect 8260 9324 8266 9376
rect 12066 9324 12072 9376
rect 12124 9324 12130 9376
rect 12176 9364 12204 9404
rect 12345 9401 12357 9435
rect 12391 9401 12403 9435
rect 12345 9395 12403 9401
rect 12526 9392 12532 9444
rect 12584 9432 12590 9444
rect 13004 9432 13032 9472
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 15010 9500 15016 9512
rect 14507 9472 15016 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14292 9432 14320 9463
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 18012 9472 18153 9500
rect 18012 9460 18018 9472
rect 18141 9469 18153 9472
rect 18187 9500 18199 9503
rect 19978 9500 19984 9512
rect 18187 9472 19984 9500
rect 18187 9469 18199 9472
rect 18141 9463 18199 9469
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 20530 9460 20536 9512
rect 20588 9500 20594 9512
rect 20824 9500 20852 9531
rect 20898 9528 20904 9580
rect 20956 9528 20962 9580
rect 21008 9568 21036 9608
rect 21082 9596 21088 9648
rect 21140 9596 21146 9648
rect 21285 9639 21343 9645
rect 21285 9636 21297 9639
rect 21192 9608 21297 9636
rect 21192 9568 21220 9608
rect 21285 9605 21297 9608
rect 21331 9605 21343 9639
rect 21285 9599 21343 9605
rect 21008 9540 21220 9568
rect 22388 9568 22416 9664
rect 24504 9646 24588 9664
rect 22557 9571 22615 9577
rect 22557 9568 22569 9571
rect 22388 9540 22569 9568
rect 22557 9537 22569 9540
rect 22603 9537 22615 9571
rect 22557 9531 22615 9537
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 22830 9568 22836 9580
rect 22787 9540 22836 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 24560 9577 24588 9646
rect 24765 9639 24823 9645
rect 24765 9605 24777 9639
rect 24811 9636 24823 9639
rect 25056 9636 25084 9667
rect 28534 9664 28540 9716
rect 28592 9704 28598 9716
rect 29825 9707 29883 9713
rect 28592 9676 29040 9704
rect 28592 9664 28598 9676
rect 24811 9608 24992 9636
rect 25056 9608 27200 9636
rect 24811 9605 24823 9608
rect 24765 9599 24823 9605
rect 24964 9580 24992 9608
rect 24535 9571 24593 9577
rect 24535 9537 24547 9571
rect 24581 9537 24593 9571
rect 24535 9531 24593 9537
rect 24670 9528 24676 9580
rect 24728 9528 24734 9580
rect 24857 9571 24915 9577
rect 24857 9537 24869 9571
rect 24903 9537 24915 9571
rect 24857 9531 24915 9537
rect 20588 9472 20852 9500
rect 20588 9460 20594 9472
rect 21266 9460 21272 9512
rect 21324 9500 21330 9512
rect 21450 9500 21456 9512
rect 21324 9472 21456 9500
rect 21324 9460 21330 9472
rect 21450 9460 21456 9472
rect 21508 9460 21514 9512
rect 14826 9432 14832 9444
rect 12584 9404 13032 9432
rect 13740 9404 13952 9432
rect 14292 9404 14832 9432
rect 12584 9392 12590 9404
rect 13740 9364 13768 9404
rect 12176 9336 13768 9364
rect 13814 9324 13820 9376
rect 13872 9324 13878 9376
rect 13924 9364 13952 9404
rect 14826 9392 14832 9404
rect 14884 9432 14890 9444
rect 14884 9404 18092 9432
rect 14884 9392 14890 9404
rect 18064 9376 18092 9404
rect 19794 9392 19800 9444
rect 19852 9392 19858 9444
rect 21468 9432 21496 9460
rect 21376 9404 21496 9432
rect 17218 9364 17224 9376
rect 13924 9336 17224 9364
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 18046 9324 18052 9376
rect 18104 9324 18110 9376
rect 20625 9367 20683 9373
rect 20625 9333 20637 9367
rect 20671 9364 20683 9367
rect 21174 9364 21180 9376
rect 20671 9336 21180 9364
rect 20671 9333 20683 9336
rect 20625 9327 20683 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 21269 9367 21327 9373
rect 21269 9333 21281 9367
rect 21315 9364 21327 9367
rect 21376 9364 21404 9404
rect 23842 9392 23848 9444
rect 23900 9432 23906 9444
rect 24872 9432 24900 9531
rect 24946 9528 24952 9580
rect 25004 9528 25010 9580
rect 25038 9528 25044 9580
rect 25096 9568 25102 9580
rect 25590 9568 25596 9580
rect 25096 9540 25596 9568
rect 25096 9528 25102 9540
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 25866 9528 25872 9580
rect 25924 9528 25930 9580
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 27172 9577 27200 9608
rect 27246 9596 27252 9648
rect 27304 9636 27310 9648
rect 29012 9636 29040 9676
rect 29825 9673 29837 9707
rect 29871 9704 29883 9707
rect 30558 9704 30564 9716
rect 29871 9676 29960 9704
rect 29871 9673 29883 9676
rect 29825 9667 29883 9673
rect 29932 9636 29960 9676
rect 30300 9676 30564 9704
rect 30190 9636 30196 9648
rect 27304 9608 28948 9636
rect 29012 9608 29868 9636
rect 29932 9608 30196 9636
rect 27304 9596 27310 9608
rect 26237 9571 26295 9577
rect 26237 9568 26249 9571
rect 26016 9540 26249 9568
rect 26016 9528 26022 9540
rect 26237 9537 26249 9540
rect 26283 9537 26295 9571
rect 26237 9531 26295 9537
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27338 9528 27344 9580
rect 27396 9568 27402 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 27396 9540 27445 9568
rect 27396 9528 27402 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27614 9528 27620 9580
rect 27672 9528 27678 9580
rect 28920 9577 28948 9608
rect 28905 9571 28963 9577
rect 28905 9537 28917 9571
rect 28951 9568 28963 9571
rect 28994 9568 29000 9580
rect 28951 9540 29000 9568
rect 28951 9537 28963 9540
rect 28905 9531 28963 9537
rect 28994 9528 29000 9540
rect 29052 9528 29058 9580
rect 29089 9571 29147 9577
rect 29089 9537 29101 9571
rect 29135 9568 29147 9571
rect 29362 9568 29368 9580
rect 29135 9540 29368 9568
rect 29135 9537 29147 9540
rect 29089 9531 29147 9537
rect 29362 9528 29368 9540
rect 29420 9528 29426 9580
rect 29733 9571 29791 9577
rect 29733 9537 29745 9571
rect 29779 9537 29791 9571
rect 29733 9531 29791 9537
rect 25884 9500 25912 9528
rect 26053 9503 26111 9509
rect 26053 9500 26065 9503
rect 25884 9472 26065 9500
rect 26053 9469 26065 9472
rect 26099 9469 26111 9503
rect 26053 9463 26111 9469
rect 26421 9503 26479 9509
rect 26421 9469 26433 9503
rect 26467 9500 26479 9503
rect 27706 9500 27712 9512
rect 26467 9472 27712 9500
rect 26467 9469 26479 9472
rect 26421 9463 26479 9469
rect 27706 9460 27712 9472
rect 27764 9460 27770 9512
rect 28534 9460 28540 9512
rect 28592 9500 28598 9512
rect 29748 9500 29776 9531
rect 28592 9472 29776 9500
rect 29840 9500 29868 9608
rect 30190 9596 30196 9608
rect 30248 9596 30254 9648
rect 29917 9571 29975 9577
rect 29917 9537 29929 9571
rect 29963 9568 29975 9571
rect 30300 9568 30328 9676
rect 30558 9664 30564 9676
rect 30616 9664 30622 9716
rect 32048 9676 32812 9704
rect 32048 9636 32076 9676
rect 29963 9540 30328 9568
rect 30392 9608 32076 9636
rect 29963 9537 29975 9540
rect 29917 9531 29975 9537
rect 30392 9500 30420 9608
rect 32214 9596 32220 9648
rect 32272 9636 32278 9648
rect 32677 9639 32735 9645
rect 32677 9636 32689 9639
rect 32272 9608 32689 9636
rect 32272 9596 32278 9608
rect 32677 9605 32689 9608
rect 32723 9605 32735 9639
rect 32784 9636 32812 9676
rect 33962 9664 33968 9716
rect 34020 9664 34026 9716
rect 32858 9636 32864 9648
rect 32784 9608 32864 9636
rect 32677 9599 32735 9605
rect 32858 9596 32864 9608
rect 32916 9596 32922 9648
rect 33045 9639 33103 9645
rect 33045 9605 33057 9639
rect 33091 9636 33103 9639
rect 33134 9636 33140 9648
rect 33091 9608 33140 9636
rect 33091 9605 33103 9608
rect 33045 9599 33103 9605
rect 33134 9596 33140 9608
rect 33192 9636 33198 9648
rect 33980 9636 34008 9664
rect 33192 9608 34008 9636
rect 33192 9596 33198 9608
rect 30834 9528 30840 9580
rect 30892 9528 30898 9580
rect 30926 9528 30932 9580
rect 30984 9568 30990 9580
rect 31205 9571 31263 9577
rect 31205 9568 31217 9571
rect 30984 9540 31217 9568
rect 30984 9528 30990 9540
rect 31205 9537 31217 9540
rect 31251 9537 31263 9571
rect 31205 9531 31263 9537
rect 31665 9571 31723 9577
rect 31665 9537 31677 9571
rect 31711 9568 31723 9571
rect 32582 9568 32588 9580
rect 31711 9540 32588 9568
rect 31711 9537 31723 9540
rect 31665 9531 31723 9537
rect 32582 9528 32588 9540
rect 32640 9528 32646 9580
rect 29840 9472 30420 9500
rect 28592 9460 28598 9472
rect 23900 9404 24900 9432
rect 23900 9392 23906 9404
rect 25038 9392 25044 9444
rect 25096 9432 25102 9444
rect 29546 9432 29552 9444
rect 25096 9404 29552 9432
rect 25096 9392 25102 9404
rect 29546 9392 29552 9404
rect 29604 9392 29610 9444
rect 21315 9336 21404 9364
rect 21453 9367 21511 9373
rect 21315 9333 21327 9336
rect 21269 9327 21327 9333
rect 21453 9333 21465 9367
rect 21499 9364 21511 9367
rect 21542 9364 21548 9376
rect 21499 9336 21548 9364
rect 21499 9333 21511 9336
rect 21453 9327 21511 9333
rect 21542 9324 21548 9336
rect 21600 9364 21606 9376
rect 21910 9364 21916 9376
rect 21600 9336 21916 9364
rect 21600 9324 21606 9336
rect 21910 9324 21916 9336
rect 21968 9324 21974 9376
rect 22738 9324 22744 9376
rect 22796 9324 22802 9376
rect 22830 9324 22836 9376
rect 22888 9364 22894 9376
rect 23566 9364 23572 9376
rect 22888 9336 23572 9364
rect 22888 9324 22894 9336
rect 23566 9324 23572 9336
rect 23624 9324 23630 9376
rect 23934 9324 23940 9376
rect 23992 9364 23998 9376
rect 24946 9364 24952 9376
rect 23992 9336 24952 9364
rect 23992 9324 23998 9336
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 25685 9367 25743 9373
rect 25685 9333 25697 9367
rect 25731 9364 25743 9367
rect 26234 9364 26240 9376
rect 25731 9336 26240 9364
rect 25731 9333 25743 9336
rect 25685 9327 25743 9333
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 26326 9324 26332 9376
rect 26384 9364 26390 9376
rect 26786 9364 26792 9376
rect 26384 9336 26792 9364
rect 26384 9324 26390 9336
rect 26786 9324 26792 9336
rect 26844 9324 26850 9376
rect 26973 9367 27031 9373
rect 26973 9333 26985 9367
rect 27019 9364 27031 9367
rect 28810 9364 28816 9376
rect 27019 9336 28816 9364
rect 27019 9333 27031 9336
rect 26973 9327 27031 9333
rect 28810 9324 28816 9336
rect 28868 9324 28874 9376
rect 29270 9324 29276 9376
rect 29328 9324 29334 9376
rect 29656 9364 29684 9472
rect 30650 9460 30656 9512
rect 30708 9460 30714 9512
rect 31202 9392 31208 9444
rect 31260 9392 31266 9444
rect 31386 9392 31392 9444
rect 31444 9432 31450 9444
rect 31938 9432 31944 9444
rect 31444 9404 31944 9432
rect 31444 9392 31450 9404
rect 31938 9392 31944 9404
rect 31996 9392 32002 9444
rect 33226 9392 33232 9444
rect 33284 9432 33290 9444
rect 34330 9432 34336 9444
rect 33284 9404 34336 9432
rect 33284 9392 33290 9404
rect 34330 9392 34336 9404
rect 34388 9392 34394 9444
rect 32030 9364 32036 9376
rect 29656 9336 32036 9364
rect 32030 9324 32036 9336
rect 32088 9324 32094 9376
rect 1104 9274 38272 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38272 9274
rect 1104 9200 38272 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1728 9132 1961 9160
rect 1728 9120 1734 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 4890 9160 4896 9172
rect 1949 9123 2007 9129
rect 4356 9132 4896 9160
rect 2317 9095 2375 9101
rect 2317 9061 2329 9095
rect 2363 9061 2375 9095
rect 3973 9095 4031 9101
rect 3973 9092 3985 9095
rect 2317 9055 2375 9061
rect 2792 9064 3985 9092
rect 1486 8916 1492 8968
rect 1544 8916 1550 8968
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2332 8956 2360 9055
rect 2792 9033 2820 9064
rect 3973 9061 3985 9064
rect 4019 9061 4031 9095
rect 3973 9055 4031 9061
rect 2777 9027 2835 9033
rect 2777 8993 2789 9027
rect 2823 8993 2835 9027
rect 2777 8987 2835 8993
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 3878 9024 3884 9036
rect 3007 8996 3884 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 3878 8984 3884 8996
rect 3936 9024 3942 9036
rect 4246 9024 4252 9036
rect 3936 8996 4252 9024
rect 3936 8984 3942 8996
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 2179 8928 2360 8956
rect 2685 8959 2743 8965
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 2731 8928 3341 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 3329 8925 3341 8928
rect 3375 8956 3387 8959
rect 4062 8956 4068 8968
rect 3375 8928 4068 8956
rect 3375 8925 3387 8928
rect 3329 8919 3387 8925
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4356 8956 4384 9132
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 5040 9132 5181 9160
rect 5040 9120 5046 9132
rect 5169 9129 5181 9132
rect 5215 9129 5227 9163
rect 5169 9123 5227 9129
rect 5350 9120 5356 9172
rect 5408 9120 5414 9172
rect 8018 9120 8024 9172
rect 8076 9120 8082 9172
rect 12066 9120 12072 9172
rect 12124 9160 12130 9172
rect 12234 9163 12292 9169
rect 12234 9160 12246 9163
rect 12124 9132 12246 9160
rect 12124 9120 12130 9132
rect 12234 9129 12246 9132
rect 12280 9129 12292 9163
rect 12234 9123 12292 9129
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 15010 9160 15016 9172
rect 12492 9132 15016 9160
rect 12492 9120 12498 9132
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 17678 9120 17684 9172
rect 17736 9120 17742 9172
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 22462 9160 22468 9172
rect 18564 9132 22468 9160
rect 18564 9120 18570 9132
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 22738 9120 22744 9172
rect 22796 9120 22802 9172
rect 22830 9120 22836 9172
rect 22888 9120 22894 9172
rect 23382 9160 23388 9172
rect 22940 9132 23388 9160
rect 5261 9095 5319 9101
rect 5261 9092 5273 9095
rect 4448 9064 5273 9092
rect 4448 9033 4476 9064
rect 5261 9061 5273 9064
rect 5307 9061 5319 9095
rect 5261 9055 5319 9061
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4433 8987 4491 8993
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 8993 4583 9027
rect 5074 9024 5080 9036
rect 4525 8987 4583 8993
rect 4632 8996 5080 9024
rect 4540 8956 4568 8987
rect 4356 8928 4568 8956
rect 3145 8891 3203 8897
rect 3145 8857 3157 8891
rect 3191 8888 3203 8891
rect 4632 8888 4660 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 4764 8928 5273 8956
rect 4764 8916 4770 8928
rect 5261 8925 5273 8928
rect 5307 8925 5319 8959
rect 5368 8956 5396 9120
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 13630 9092 13636 9104
rect 5500 9064 10456 9092
rect 5500 9052 5506 9064
rect 8202 8984 8208 9036
rect 8260 8984 8266 9036
rect 10318 9024 10324 9036
rect 9876 8996 10324 9024
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5368 8928 5457 8956
rect 5261 8919 5319 8925
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 8570 8956 8576 8968
rect 8343 8928 8576 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9876 8965 9904 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 9953 8959 10011 8965
rect 9953 8925 9965 8959
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 4801 8891 4859 8897
rect 4801 8888 4813 8891
rect 3191 8860 4813 8888
rect 3191 8857 3203 8860
rect 3145 8851 3203 8857
rect 4801 8857 4813 8860
rect 4847 8857 4859 8891
rect 4801 8851 4859 8857
rect 4890 8848 4896 8900
rect 4948 8888 4954 8900
rect 4985 8891 5043 8897
rect 4985 8888 4997 8891
rect 4948 8860 4997 8888
rect 4948 8848 4954 8860
rect 4985 8857 4997 8860
rect 5031 8857 5043 8891
rect 4985 8851 5043 8857
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 8389 8891 8447 8897
rect 8389 8888 8401 8891
rect 8260 8860 8401 8888
rect 8260 8848 8266 8860
rect 8389 8857 8401 8860
rect 8435 8857 8447 8891
rect 8389 8851 8447 8857
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9968 8888 9996 8919
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8956 10287 8959
rect 10428 8956 10456 9064
rect 11164 9064 12112 9092
rect 11164 9036 11192 9064
rect 11146 8984 11152 9036
rect 11204 8984 11210 9036
rect 12084 9024 12112 9064
rect 13280 9064 13636 9092
rect 13280 9036 13308 9064
rect 13630 9052 13636 9064
rect 13688 9092 13694 9104
rect 13688 9064 15516 9092
rect 13688 9052 13694 9064
rect 12802 9024 12808 9036
rect 12084 8996 12808 9024
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 13262 8984 13268 9036
rect 13320 8984 13326 9036
rect 15488 9033 15516 9064
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 22848 9092 22876 9120
rect 17276 9064 22876 9092
rect 17276 9052 17282 9064
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 8993 15531 9027
rect 17773 9027 17831 9033
rect 15473 8987 15531 8993
rect 17328 8996 17724 9024
rect 10275 8928 10456 8956
rect 10275 8925 10287 8928
rect 10229 8919 10287 8925
rect 8536 8860 9996 8888
rect 10244 8888 10272 8919
rect 11974 8916 11980 8968
rect 12032 8916 12038 8968
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 14458 8956 14464 8968
rect 14332 8928 14464 8956
rect 14332 8916 14338 8928
rect 14458 8916 14464 8928
rect 14516 8956 14522 8968
rect 17328 8965 17356 8996
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14516 8928 15301 8956
rect 14516 8916 14522 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 15289 8919 15347 8925
rect 16408 8928 17325 8956
rect 13538 8888 13544 8900
rect 10244 8860 12434 8888
rect 13478 8860 13544 8888
rect 8536 8848 8542 8860
rect 12406 8832 12434 8860
rect 13538 8848 13544 8860
rect 13596 8888 13602 8900
rect 13596 8860 14688 8888
rect 13596 8848 13602 8860
rect 14660 8832 14688 8860
rect 15010 8848 15016 8900
rect 15068 8888 15074 8900
rect 16408 8888 16436 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 17494 8916 17500 8968
rect 17552 8916 17558 8968
rect 17696 8956 17724 8996
rect 17773 8993 17785 9027
rect 17819 9024 17831 9027
rect 17862 9024 17868 9036
rect 17819 8996 17868 9024
rect 17819 8993 17831 8996
rect 17773 8987 17831 8993
rect 17862 8984 17868 8996
rect 17920 8984 17926 9036
rect 20622 8984 20628 9036
rect 20680 8984 20686 9036
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 22940 9033 22968 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 23658 9120 23664 9172
rect 23716 9160 23722 9172
rect 23753 9163 23811 9169
rect 23753 9160 23765 9163
rect 23716 9132 23765 9160
rect 23716 9120 23722 9132
rect 23753 9129 23765 9132
rect 23799 9160 23811 9163
rect 26326 9160 26332 9172
rect 23799 9132 26332 9160
rect 23799 9129 23811 9132
rect 23753 9123 23811 9129
rect 26326 9120 26332 9132
rect 26384 9160 26390 9172
rect 26384 9132 26648 9160
rect 26384 9120 26390 9132
rect 24302 9092 24308 9104
rect 23216 9064 24308 9092
rect 21177 9027 21235 9033
rect 21177 9024 21189 9027
rect 20956 8996 21189 9024
rect 20956 8984 20962 8996
rect 21177 8993 21189 8996
rect 21223 8993 21235 9027
rect 22925 9027 22983 9033
rect 22925 9024 22937 9027
rect 21177 8987 21235 8993
rect 22066 8996 22937 9024
rect 17954 8956 17960 8968
rect 17696 8928 17960 8956
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 18104 8928 19349 8956
rect 18104 8916 18110 8928
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 19576 8928 20177 8956
rect 19576 8916 19582 8928
rect 20165 8925 20177 8928
rect 20211 8925 20223 8959
rect 20165 8919 20223 8925
rect 20530 8916 20536 8968
rect 20588 8916 20594 8968
rect 20640 8956 20668 8984
rect 20806 8956 20812 8968
rect 20640 8928 20812 8956
rect 20806 8916 20812 8928
rect 20864 8956 20870 8968
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 20864 8928 21097 8956
rect 20864 8916 20870 8928
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21085 8919 21143 8925
rect 15068 8860 16436 8888
rect 15068 8848 15074 8860
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 18141 8891 18199 8897
rect 18141 8888 18153 8891
rect 16540 8860 18153 8888
rect 16540 8848 16546 8860
rect 18141 8857 18153 8860
rect 18187 8857 18199 8891
rect 18141 8851 18199 8857
rect 18322 8848 18328 8900
rect 18380 8848 18386 8900
rect 22066 8888 22094 8996
rect 22925 8993 22937 8996
rect 22971 9024 22983 9027
rect 23106 9024 23112 9036
rect 22971 8996 23112 9024
rect 22971 8993 22983 8996
rect 22925 8987 22983 8993
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 22554 8916 22560 8968
rect 22612 8916 22618 8968
rect 22830 8916 22836 8968
rect 22888 8956 22894 8968
rect 23017 8959 23075 8965
rect 23017 8956 23029 8959
rect 22888 8928 23029 8956
rect 22888 8916 22894 8928
rect 23017 8925 23029 8928
rect 23063 8925 23075 8959
rect 23216 8956 23244 9064
rect 24302 9052 24308 9064
rect 24360 9092 24366 9104
rect 26418 9092 26424 9104
rect 24360 9064 24900 9092
rect 24360 9052 24366 9064
rect 23290 8984 23296 9036
rect 23348 9024 23354 9036
rect 24762 9024 24768 9036
rect 23348 8996 24768 9024
rect 23348 8984 23354 8996
rect 23385 8959 23443 8965
rect 23385 8956 23397 8959
rect 23216 8928 23397 8956
rect 23017 8919 23075 8925
rect 23385 8925 23397 8928
rect 23431 8956 23443 8959
rect 23661 8959 23719 8965
rect 23661 8956 23673 8959
rect 23431 8928 23673 8956
rect 23431 8925 23443 8928
rect 23385 8919 23443 8925
rect 23661 8925 23673 8928
rect 23707 8925 23719 8959
rect 23934 8956 23940 8968
rect 23661 8919 23719 8925
rect 23768 8928 23940 8956
rect 20732 8860 22094 8888
rect 22572 8888 22600 8916
rect 23768 8888 23796 8928
rect 23934 8916 23940 8928
rect 23992 8956 23998 8968
rect 24029 8959 24087 8965
rect 24029 8956 24041 8959
rect 23992 8928 24041 8956
rect 23992 8916 23998 8928
rect 24029 8925 24041 8928
rect 24075 8925 24087 8959
rect 24029 8919 24087 8925
rect 24118 8916 24124 8968
rect 24176 8916 24182 8968
rect 24213 8959 24271 8965
rect 24213 8925 24225 8959
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 22572 8860 23796 8888
rect 934 8780 940 8832
rect 992 8820 998 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 992 8792 1593 8820
rect 992 8780 998 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 3510 8780 3516 8832
rect 3568 8780 3574 8832
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 8294 8820 8300 8832
rect 4387 8792 8300 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9490 8820 9496 8832
rect 8812 8792 9496 8820
rect 8812 8780 8818 8792
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9582 8780 9588 8832
rect 9640 8780 9646 8832
rect 12406 8792 12440 8832
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 13725 8823 13783 8829
rect 13725 8820 13737 8823
rect 12676 8792 13737 8820
rect 12676 8780 12682 8792
rect 13725 8789 13737 8792
rect 13771 8789 13783 8823
rect 13725 8783 13783 8789
rect 14642 8780 14648 8832
rect 14700 8780 14706 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15194 8820 15200 8832
rect 14967 8792 15200 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 15381 8823 15439 8829
rect 15381 8789 15393 8823
rect 15427 8820 15439 8823
rect 18340 8820 18368 8848
rect 15427 8792 18368 8820
rect 15427 8789 15439 8792
rect 15381 8783 15439 8789
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 20622 8820 20628 8832
rect 20220 8792 20628 8820
rect 20220 8780 20226 8792
rect 20622 8780 20628 8792
rect 20680 8820 20686 8832
rect 20732 8829 20760 8860
rect 23842 8848 23848 8900
rect 23900 8888 23906 8900
rect 24228 8888 24256 8919
rect 24394 8916 24400 8968
rect 24452 8916 24458 8968
rect 24504 8965 24532 8996
rect 24762 8984 24768 8996
rect 24820 8984 24826 9036
rect 24872 8965 24900 9064
rect 25424 9064 26424 9092
rect 24490 8959 24548 8965
rect 24490 8925 24502 8959
rect 24536 8925 24548 8959
rect 24490 8919 24548 8925
rect 24862 8959 24920 8965
rect 24862 8925 24874 8959
rect 24908 8925 24920 8959
rect 25424 8956 25452 9064
rect 26418 9052 26424 9064
rect 26476 9052 26482 9104
rect 25774 8984 25780 9036
rect 25832 8984 25838 9036
rect 26620 9024 26648 9132
rect 27154 9120 27160 9172
rect 27212 9120 27218 9172
rect 27617 9163 27675 9169
rect 27617 9129 27629 9163
rect 27663 9160 27675 9163
rect 28718 9160 28724 9172
rect 27663 9132 28724 9160
rect 27663 9129 27675 9132
rect 27617 9123 27675 9129
rect 28718 9120 28724 9132
rect 28776 9120 28782 9172
rect 29270 9120 29276 9172
rect 29328 9160 29334 9172
rect 29733 9163 29791 9169
rect 29733 9160 29745 9163
rect 29328 9132 29745 9160
rect 29328 9120 29334 9132
rect 29733 9129 29745 9132
rect 29779 9129 29791 9163
rect 29733 9123 29791 9129
rect 27172 9092 27200 9120
rect 29748 9092 29776 9123
rect 30834 9120 30840 9172
rect 30892 9160 30898 9172
rect 31849 9163 31907 9169
rect 31849 9160 31861 9163
rect 30892 9132 31861 9160
rect 30892 9120 30898 9132
rect 31849 9129 31861 9132
rect 31895 9129 31907 9163
rect 31849 9123 31907 9129
rect 32582 9120 32588 9172
rect 32640 9120 32646 9172
rect 33045 9163 33103 9169
rect 33045 9129 33057 9163
rect 33091 9160 33103 9163
rect 33134 9160 33140 9172
rect 33091 9132 33140 9160
rect 33091 9129 33103 9132
rect 33045 9123 33103 9129
rect 33134 9120 33140 9132
rect 33192 9120 33198 9172
rect 33505 9163 33563 9169
rect 33505 9129 33517 9163
rect 33551 9160 33563 9163
rect 33594 9160 33600 9172
rect 33551 9132 33600 9160
rect 33551 9129 33563 9132
rect 33505 9123 33563 9129
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 27172 9064 27476 9092
rect 26252 8996 26556 9024
rect 26620 8996 27292 9024
rect 26252 8968 26280 8996
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25424 8928 25513 8956
rect 24862 8919 24920 8925
rect 25501 8925 25513 8928
rect 25547 8925 25559 8959
rect 25501 8919 25559 8925
rect 25590 8916 25596 8968
rect 25648 8916 25654 8968
rect 25682 8916 25688 8968
rect 25740 8956 25746 8968
rect 25869 8959 25927 8965
rect 25869 8956 25881 8959
rect 25740 8928 25881 8956
rect 25740 8916 25746 8928
rect 25869 8925 25881 8928
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 26234 8916 26240 8968
rect 26292 8916 26298 8968
rect 26326 8916 26332 8968
rect 26384 8916 26390 8968
rect 26421 8959 26479 8965
rect 26421 8925 26433 8959
rect 26467 8925 26479 8959
rect 26421 8919 26479 8925
rect 24670 8888 24676 8900
rect 23900 8860 24256 8888
rect 24320 8860 24676 8888
rect 23900 8848 23906 8860
rect 20717 8823 20775 8829
rect 20717 8820 20729 8823
rect 20680 8792 20729 8820
rect 20680 8780 20686 8792
rect 20717 8789 20729 8792
rect 20763 8789 20775 8823
rect 20717 8783 20775 8789
rect 21358 8780 21364 8832
rect 21416 8780 21422 8832
rect 23014 8780 23020 8832
rect 23072 8820 23078 8832
rect 24320 8820 24348 8860
rect 24670 8848 24676 8860
rect 24728 8848 24734 8900
rect 24765 8891 24823 8897
rect 24765 8857 24777 8891
rect 24811 8888 24823 8891
rect 25317 8891 25375 8897
rect 24811 8860 25268 8888
rect 24811 8857 24823 8860
rect 24765 8851 24823 8857
rect 23072 8792 24348 8820
rect 23072 8780 23078 8792
rect 24486 8780 24492 8832
rect 24544 8820 24550 8832
rect 24780 8820 24808 8851
rect 24544 8792 24808 8820
rect 25041 8823 25099 8829
rect 24544 8780 24550 8792
rect 25041 8789 25053 8823
rect 25087 8820 25099 8823
rect 25130 8820 25136 8832
rect 25087 8792 25136 8820
rect 25087 8789 25099 8792
rect 25041 8783 25099 8789
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 25240 8820 25268 8860
rect 25317 8857 25329 8891
rect 25363 8888 25375 8891
rect 26436 8888 26464 8919
rect 25363 8860 26464 8888
rect 26528 8888 26556 8996
rect 26605 8959 26663 8965
rect 26605 8925 26617 8959
rect 26651 8956 26663 8959
rect 26786 8956 26792 8968
rect 26651 8928 26792 8956
rect 26651 8925 26663 8928
rect 26605 8919 26663 8925
rect 26786 8916 26792 8928
rect 26844 8916 26850 8968
rect 26878 8916 26884 8968
rect 26936 8916 26942 8968
rect 26970 8916 26976 8968
rect 27028 8956 27034 8968
rect 27264 8965 27292 8996
rect 27448 8965 27476 9064
rect 27816 9064 28994 9092
rect 29748 9064 31754 9092
rect 27816 9036 27844 9064
rect 27798 8984 27804 9036
rect 27856 8984 27862 9036
rect 28442 8965 28448 8968
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 27028 8928 27077 8956
rect 27028 8916 27034 8928
rect 27065 8925 27077 8928
rect 27111 8925 27123 8959
rect 27065 8919 27123 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 27249 8959 27307 8965
rect 27249 8925 27261 8959
rect 27295 8925 27307 8959
rect 27249 8919 27307 8925
rect 27433 8959 27491 8965
rect 27433 8925 27445 8959
rect 27479 8925 27491 8959
rect 27433 8919 27491 8925
rect 28425 8959 28448 8965
rect 28425 8925 28437 8959
rect 28425 8919 28448 8925
rect 27172 8888 27200 8919
rect 28442 8916 28448 8919
rect 28500 8916 28506 8968
rect 28552 8965 28580 9064
rect 28537 8959 28595 8965
rect 28537 8925 28549 8959
rect 28583 8925 28595 8959
rect 28537 8919 28595 8925
rect 28629 8959 28687 8965
rect 28629 8925 28641 8959
rect 28675 8925 28687 8959
rect 28629 8919 28687 8925
rect 28644 8888 28672 8919
rect 28810 8916 28816 8968
rect 28868 8916 28874 8968
rect 28718 8888 28724 8900
rect 26528 8860 27292 8888
rect 28644 8860 28724 8888
rect 25363 8857 25375 8860
rect 25317 8851 25375 8857
rect 27264 8832 27292 8860
rect 28718 8848 28724 8860
rect 28776 8848 28782 8900
rect 28966 8888 28994 9064
rect 29086 8984 29092 9036
rect 29144 9024 29150 9036
rect 29641 9027 29699 9033
rect 29641 9024 29653 9027
rect 29144 8996 29653 9024
rect 29144 8984 29150 8996
rect 29641 8993 29653 8996
rect 29687 9024 29699 9027
rect 31386 9024 31392 9036
rect 29687 8996 31392 9024
rect 29687 8993 29699 8996
rect 29641 8987 29699 8993
rect 31386 8984 31392 8996
rect 31444 8984 31450 9036
rect 31726 9024 31754 9064
rect 32030 9052 32036 9104
rect 32088 9092 32094 9104
rect 32217 9095 32275 9101
rect 32217 9092 32229 9095
rect 32088 9064 32229 9092
rect 32088 9052 32094 9064
rect 32217 9061 32229 9064
rect 32263 9061 32275 9095
rect 32217 9055 32275 9061
rect 33060 9064 33548 9092
rect 32950 9024 32956 9036
rect 31726 8996 32956 9024
rect 29546 8916 29552 8968
rect 29604 8956 29610 8968
rect 30098 8956 30104 8968
rect 29604 8928 30104 8956
rect 29604 8916 29610 8928
rect 30098 8916 30104 8928
rect 30156 8916 30162 8968
rect 30374 8916 30380 8968
rect 30432 8916 30438 8968
rect 31573 8959 31631 8965
rect 31573 8956 31585 8959
rect 31404 8928 31585 8956
rect 30392 8888 30420 8916
rect 31404 8900 31432 8928
rect 31573 8925 31585 8928
rect 31619 8925 31631 8959
rect 31573 8919 31631 8925
rect 31665 8959 31723 8965
rect 31665 8925 31677 8959
rect 31711 8956 31723 8959
rect 31846 8956 31852 8968
rect 31711 8928 31852 8956
rect 31711 8925 31723 8928
rect 31665 8919 31723 8925
rect 28966 8860 30420 8888
rect 31386 8848 31392 8900
rect 31444 8848 31450 8900
rect 31588 8888 31616 8919
rect 31846 8916 31852 8928
rect 31904 8916 31910 8968
rect 31938 8916 31944 8968
rect 31996 8916 32002 8968
rect 32140 8965 32168 8996
rect 32950 8984 32956 8996
rect 33008 9024 33014 9036
rect 33060 9024 33088 9064
rect 33008 8996 33088 9024
rect 33008 8984 33014 8996
rect 32125 8959 32183 8965
rect 32125 8925 32137 8959
rect 32171 8925 32183 8959
rect 32125 8919 32183 8925
rect 32490 8916 32496 8968
rect 32548 8956 32554 8968
rect 32769 8959 32827 8965
rect 32769 8956 32781 8959
rect 32548 8928 32781 8956
rect 32548 8916 32554 8928
rect 32769 8925 32781 8928
rect 32815 8925 32827 8959
rect 32769 8919 32827 8925
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8925 32919 8959
rect 32861 8919 32919 8925
rect 32214 8888 32220 8900
rect 31588 8860 32220 8888
rect 32214 8848 32220 8860
rect 32272 8848 32278 8900
rect 32876 8888 32904 8919
rect 33134 8916 33140 8968
rect 33192 8916 33198 8968
rect 33520 8965 33548 9064
rect 36630 8984 36636 9036
rect 36688 9024 36694 9036
rect 37645 9027 37703 9033
rect 37645 9024 37657 9027
rect 36688 8996 37657 9024
rect 36688 8984 36694 8996
rect 37645 8993 37657 8996
rect 37691 8993 37703 9027
rect 37645 8987 37703 8993
rect 33229 8959 33287 8965
rect 33229 8925 33241 8959
rect 33275 8925 33287 8959
rect 33229 8919 33287 8925
rect 33505 8959 33563 8965
rect 33505 8925 33517 8959
rect 33551 8925 33563 8959
rect 33505 8919 33563 8925
rect 33689 8959 33747 8965
rect 33689 8925 33701 8959
rect 33735 8956 33747 8959
rect 33778 8956 33784 8968
rect 33735 8928 33784 8956
rect 33735 8925 33747 8928
rect 33689 8919 33747 8925
rect 33244 8888 33272 8919
rect 33778 8916 33784 8928
rect 33836 8916 33842 8968
rect 37461 8959 37519 8965
rect 37461 8925 37473 8959
rect 37507 8956 37519 8959
rect 38102 8956 38108 8968
rect 37507 8928 38108 8956
rect 37507 8925 37519 8928
rect 37461 8919 37519 8925
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 32876 8860 33272 8888
rect 33152 8832 33180 8860
rect 25682 8820 25688 8832
rect 25240 8792 25688 8820
rect 25682 8780 25688 8792
rect 25740 8780 25746 8832
rect 25958 8780 25964 8832
rect 26016 8780 26022 8832
rect 26234 8780 26240 8832
rect 26292 8820 26298 8832
rect 26970 8820 26976 8832
rect 26292 8792 26976 8820
rect 26292 8780 26298 8792
rect 26970 8780 26976 8792
rect 27028 8780 27034 8832
rect 27246 8780 27252 8832
rect 27304 8780 27310 8832
rect 28169 8823 28227 8829
rect 28169 8789 28181 8823
rect 28215 8820 28227 8823
rect 29178 8820 29184 8832
rect 28215 8792 29184 8820
rect 28215 8789 28227 8792
rect 28169 8783 28227 8789
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 29914 8780 29920 8832
rect 29972 8780 29978 8832
rect 30834 8780 30840 8832
rect 30892 8820 30898 8832
rect 31205 8823 31263 8829
rect 31205 8820 31217 8823
rect 30892 8792 31217 8820
rect 30892 8780 30898 8792
rect 31205 8789 31217 8792
rect 31251 8789 31263 8823
rect 31205 8783 31263 8789
rect 33134 8780 33140 8832
rect 33192 8780 33198 8832
rect 1104 8730 38272 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38272 8730
rect 1104 8656 38272 8678
rect 2866 8576 2872 8628
rect 2924 8576 2930 8628
rect 3510 8576 3516 8628
rect 3568 8576 3574 8628
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4541 8619 4599 8625
rect 4541 8616 4553 8619
rect 4120 8588 4553 8616
rect 4120 8576 4126 8588
rect 4541 8585 4553 8588
rect 4587 8585 4599 8619
rect 4541 8579 4599 8585
rect 4706 8576 4712 8628
rect 4764 8576 4770 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7653 8619 7711 8625
rect 7653 8616 7665 8619
rect 7147 8588 7665 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7653 8585 7665 8588
rect 7699 8585 7711 8619
rect 7653 8579 7711 8585
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 8754 8616 8760 8628
rect 8067 8588 8760 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 10042 8616 10048 8628
rect 8895 8588 10048 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 13814 8616 13820 8628
rect 12406 8588 13820 8616
rect 2884 8548 2912 8576
rect 3528 8548 3556 8576
rect 2884 8520 3004 8548
rect 2976 8489 3004 8520
rect 3068 8520 3556 8548
rect 4341 8551 4399 8557
rect 3068 8489 3096 8520
rect 4341 8517 4353 8551
rect 4387 8517 4399 8551
rect 4341 8511 4399 8517
rect 5184 8520 8248 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2869 8483 2927 8489
rect 2869 8480 2881 8483
rect 2363 8452 2881 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2746 8412 2774 8452
rect 2869 8449 2881 8452
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 4356 8480 4384 8511
rect 5184 8492 5212 8520
rect 4706 8480 4712 8492
rect 4356 8452 4712 8480
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6932 8452 7021 8480
rect 4080 8412 4108 8440
rect 2746 8384 4108 8412
rect 2590 8304 2596 8356
rect 2648 8304 2654 8356
rect 6932 8344 6960 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7190 8372 7196 8424
rect 7248 8372 7254 8424
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 8220 8421 8248 8520
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 12406 8548 12434 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 14608 8588 16528 8616
rect 14608 8576 14614 8588
rect 14568 8548 14596 8576
rect 8352 8520 12434 8548
rect 14384 8520 14596 8548
rect 8352 8508 8358 8520
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8536 8452 8677 8480
rect 8536 8440 8542 8452
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8665 8443 8723 8449
rect 8772 8452 8861 8480
rect 8113 8415 8171 8421
rect 8113 8412 8125 8415
rect 7984 8384 8125 8412
rect 7984 8372 7990 8384
rect 8113 8381 8125 8384
rect 8159 8381 8171 8415
rect 8113 8375 8171 8381
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 7466 8344 7472 8356
rect 6564 8316 7472 8344
rect 4525 8279 4583 8285
rect 4525 8245 4537 8279
rect 4571 8276 4583 8279
rect 4982 8276 4988 8288
rect 4571 8248 4988 8276
rect 4571 8245 4583 8248
rect 4525 8239 4583 8245
rect 4982 8236 4988 8248
rect 5040 8276 5046 8288
rect 6564 8276 6592 8316
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 8128 8344 8156 8375
rect 8772 8344 8800 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 12345 8483 12403 8489
rect 12345 8480 12357 8483
rect 11940 8452 12357 8480
rect 11940 8440 11946 8452
rect 12345 8449 12357 8452
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 14274 8440 14280 8492
rect 14332 8440 14338 8492
rect 14384 8489 14412 8520
rect 14642 8508 14648 8560
rect 14700 8548 14706 8560
rect 14700 8520 15134 8548
rect 14700 8508 14706 8520
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8449 14427 8483
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 14369 8443 14427 8449
rect 15856 8452 16405 8480
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 14384 8412 14412 8443
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 12032 8384 14412 8412
rect 14476 8384 14657 8412
rect 12032 8372 12038 8384
rect 8128 8316 8800 8344
rect 12406 8288 12434 8384
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8344 14151 8347
rect 14476 8344 14504 8384
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 15194 8372 15200 8424
rect 15252 8412 15258 8424
rect 15856 8412 15884 8452
rect 16393 8449 16405 8452
rect 16439 8449 16451 8483
rect 16500 8480 16528 8588
rect 16666 8576 16672 8628
rect 16724 8576 16730 8628
rect 19978 8616 19984 8628
rect 19536 8588 19984 8616
rect 16684 8548 16712 8576
rect 16684 8520 17434 8548
rect 18322 8508 18328 8560
rect 18380 8548 18386 8560
rect 19245 8551 19303 8557
rect 19245 8548 19257 8551
rect 18380 8520 19257 8548
rect 18380 8508 18386 8520
rect 19245 8517 19257 8520
rect 19291 8517 19303 8551
rect 19245 8511 19303 8517
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16500 8452 16681 8480
rect 16393 8443 16451 8449
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 16669 8443 16727 8449
rect 18432 8452 18521 8480
rect 15252 8384 15884 8412
rect 15252 8372 15258 8384
rect 16114 8372 16120 8424
rect 16172 8372 16178 8424
rect 18432 8421 18460 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 19334 8440 19340 8492
rect 19392 8480 19398 8492
rect 19536 8489 19564 8588
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20806 8616 20812 8628
rect 20128 8588 20812 8616
rect 20128 8576 20134 8588
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 22830 8616 22836 8628
rect 22480 8588 22836 8616
rect 19613 8551 19671 8557
rect 19613 8517 19625 8551
rect 19659 8548 19671 8551
rect 19659 8520 22416 8548
rect 19659 8517 19671 8520
rect 19613 8511 19671 8517
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19392 8452 19533 8480
rect 19392 8440 19398 8452
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 16945 8415 17003 8421
rect 16945 8412 16957 8415
rect 16224 8384 16957 8412
rect 16132 8344 16160 8372
rect 16224 8353 16252 8384
rect 16945 8381 16957 8384
rect 16991 8381 17003 8415
rect 16945 8375 17003 8381
rect 18417 8415 18475 8421
rect 18417 8381 18429 8415
rect 18463 8381 18475 8415
rect 18417 8375 18475 8381
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 19720 8412 19748 8443
rect 20070 8440 20076 8492
rect 20128 8440 20134 8492
rect 20162 8440 20168 8492
rect 20220 8440 20226 8492
rect 20254 8440 20260 8492
rect 20312 8440 20318 8492
rect 20622 8440 20628 8492
rect 20680 8440 20686 8492
rect 20898 8440 20904 8492
rect 20956 8440 20962 8492
rect 22388 8489 22416 8520
rect 22480 8489 22508 8588
rect 22830 8576 22836 8588
rect 22888 8616 22894 8628
rect 23198 8616 23204 8628
rect 22888 8588 23204 8616
rect 22888 8576 22894 8588
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 23842 8616 23848 8628
rect 23624 8588 23848 8616
rect 23624 8576 23630 8588
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 24118 8576 24124 8628
rect 24176 8616 24182 8628
rect 25133 8619 25191 8625
rect 25133 8616 25145 8619
rect 24176 8588 25145 8616
rect 24176 8576 24182 8588
rect 25133 8585 25145 8588
rect 25179 8616 25191 8619
rect 26234 8616 26240 8628
rect 25179 8588 26240 8616
rect 25179 8585 25191 8588
rect 25133 8579 25191 8585
rect 26234 8576 26240 8588
rect 26292 8576 26298 8628
rect 26878 8576 26884 8628
rect 26936 8616 26942 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26936 8588 27353 8616
rect 26936 8576 26942 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27341 8579 27399 8585
rect 28166 8576 28172 8628
rect 28224 8576 28230 8628
rect 28905 8619 28963 8625
rect 28905 8585 28917 8619
rect 28951 8616 28963 8619
rect 29546 8616 29552 8628
rect 28951 8588 29552 8616
rect 28951 8585 28963 8588
rect 28905 8579 28963 8585
rect 29546 8576 29552 8588
rect 29604 8576 29610 8628
rect 29914 8576 29920 8628
rect 29972 8576 29978 8628
rect 30650 8576 30656 8628
rect 30708 8616 30714 8628
rect 31389 8619 31447 8625
rect 31389 8616 31401 8619
rect 30708 8588 31401 8616
rect 30708 8576 30714 8588
rect 31389 8585 31401 8588
rect 31435 8616 31447 8619
rect 31754 8616 31760 8628
rect 31435 8588 31760 8616
rect 31435 8585 31447 8588
rect 31389 8579 31447 8585
rect 31754 8576 31760 8588
rect 31812 8576 31818 8628
rect 32950 8576 32956 8628
rect 33008 8576 33014 8628
rect 23290 8548 23296 8560
rect 22572 8520 23296 8548
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8449 22431 8483
rect 22373 8443 22431 8449
rect 22465 8483 22523 8489
rect 22465 8449 22477 8483
rect 22511 8449 22523 8483
rect 22465 8443 22523 8449
rect 19208 8384 19748 8412
rect 19208 8372 19214 8384
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20916 8412 20944 8440
rect 20036 8384 20944 8412
rect 22388 8412 22416 8443
rect 22572 8412 22600 8520
rect 23290 8508 23296 8520
rect 23348 8508 23354 8560
rect 24946 8508 24952 8560
rect 25004 8548 25010 8560
rect 27157 8551 27215 8557
rect 25004 8520 27108 8548
rect 25004 8508 25010 8520
rect 22646 8440 22652 8492
rect 22704 8480 22710 8492
rect 23106 8489 23112 8492
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 22704 8452 22845 8480
rect 22704 8440 22710 8452
rect 22833 8449 22845 8452
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8449 22983 8483
rect 22925 8443 22983 8449
rect 23073 8483 23112 8489
rect 23073 8449 23085 8483
rect 23073 8443 23112 8449
rect 22388 8384 22600 8412
rect 20036 8372 20042 8384
rect 22738 8372 22744 8424
rect 22796 8372 22802 8424
rect 14139 8316 14504 8344
rect 15672 8316 16160 8344
rect 16209 8347 16267 8353
rect 14139 8313 14151 8316
rect 14093 8307 14151 8313
rect 5040 8248 6592 8276
rect 5040 8236 5046 8248
rect 6638 8236 6644 8288
rect 6696 8236 6702 8288
rect 12342 8236 12348 8288
rect 12400 8248 12434 8288
rect 12621 8279 12679 8285
rect 12400 8236 12406 8248
rect 12621 8245 12633 8279
rect 12667 8276 12679 8279
rect 13262 8276 13268 8288
rect 12667 8248 13268 8276
rect 12667 8245 12679 8248
rect 12621 8239 12679 8245
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 15672 8276 15700 8316
rect 16209 8313 16221 8347
rect 16255 8313 16267 8347
rect 16209 8307 16267 8313
rect 19797 8347 19855 8353
rect 19797 8313 19809 8347
rect 19843 8344 19855 8347
rect 19886 8344 19892 8356
rect 19843 8316 19892 8344
rect 19843 8313 19855 8316
rect 19797 8307 19855 8313
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 22189 8347 22247 8353
rect 22189 8313 22201 8347
rect 22235 8344 22247 8347
rect 22940 8344 22968 8443
rect 23106 8440 23112 8443
rect 23164 8440 23170 8492
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 23431 8483 23489 8489
rect 23431 8449 23443 8483
rect 23477 8480 23489 8483
rect 23750 8480 23756 8492
rect 23477 8452 23756 8480
rect 23477 8449 23489 8452
rect 23431 8443 23489 8449
rect 23216 8412 23244 8443
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 25774 8480 25780 8492
rect 25240 8452 25780 8480
rect 25240 8421 25268 8452
rect 25774 8440 25780 8452
rect 25832 8480 25838 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 25832 8452 26985 8480
rect 25832 8440 25838 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 27080 8480 27108 8520
rect 27157 8517 27169 8551
rect 27203 8548 27215 8551
rect 27706 8548 27712 8560
rect 27203 8520 27712 8548
rect 27203 8517 27215 8520
rect 27157 8511 27215 8517
rect 27706 8508 27712 8520
rect 27764 8548 27770 8560
rect 28184 8548 28212 8576
rect 29362 8548 29368 8560
rect 27764 8520 28212 8548
rect 28276 8520 29368 8548
rect 27764 8508 27770 8520
rect 28276 8480 28304 8520
rect 29362 8508 29368 8520
rect 29420 8508 29426 8560
rect 27080 8452 28304 8480
rect 26973 8443 27031 8449
rect 28350 8440 28356 8492
rect 28408 8440 28414 8492
rect 28537 8483 28595 8489
rect 28537 8449 28549 8483
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 25225 8415 25283 8421
rect 25225 8412 25237 8415
rect 23032 8384 23244 8412
rect 23400 8384 25237 8412
rect 23032 8356 23060 8384
rect 22235 8316 22968 8344
rect 22235 8313 22247 8316
rect 22189 8307 22247 8313
rect 23014 8304 23020 8356
rect 23072 8304 23078 8356
rect 23198 8304 23204 8356
rect 23256 8344 23262 8356
rect 23400 8344 23428 8384
rect 25225 8381 25237 8384
rect 25271 8381 25283 8415
rect 25225 8375 25283 8381
rect 25317 8415 25375 8421
rect 25317 8381 25329 8415
rect 25363 8412 25375 8415
rect 25590 8412 25596 8424
rect 25363 8384 25596 8412
rect 25363 8381 25375 8384
rect 25317 8375 25375 8381
rect 23256 8316 23428 8344
rect 24765 8347 24823 8353
rect 23256 8304 23262 8316
rect 24765 8313 24777 8347
rect 24811 8344 24823 8347
rect 24946 8344 24952 8356
rect 24811 8316 24952 8344
rect 24811 8313 24823 8316
rect 24765 8307 24823 8313
rect 24946 8304 24952 8316
rect 25004 8304 25010 8356
rect 14792 8248 15700 8276
rect 20441 8279 20499 8285
rect 14792 8236 14798 8248
rect 20441 8245 20453 8279
rect 20487 8276 20499 8279
rect 20806 8276 20812 8288
rect 20487 8248 20812 8276
rect 20487 8245 20499 8248
rect 20441 8239 20499 8245
rect 20806 8236 20812 8248
rect 20864 8236 20870 8288
rect 23566 8236 23572 8288
rect 23624 8236 23630 8288
rect 23934 8236 23940 8288
rect 23992 8276 23998 8288
rect 25332 8276 25360 8375
rect 25590 8372 25596 8384
rect 25648 8372 25654 8424
rect 26878 8372 26884 8424
rect 26936 8412 26942 8424
rect 28552 8412 28580 8443
rect 28718 8440 28724 8492
rect 28776 8440 28782 8492
rect 28810 8440 28816 8492
rect 28868 8440 28874 8492
rect 29932 8489 29960 8576
rect 28997 8483 29055 8489
rect 28997 8449 29009 8483
rect 29043 8449 29055 8483
rect 28997 8443 29055 8449
rect 29917 8483 29975 8489
rect 29917 8449 29929 8483
rect 29963 8449 29975 8483
rect 29917 8443 29975 8449
rect 26936 8384 28580 8412
rect 28736 8412 28764 8440
rect 29012 8412 29040 8443
rect 30006 8440 30012 8492
rect 30064 8480 30070 8492
rect 30101 8483 30159 8489
rect 30101 8480 30113 8483
rect 30064 8452 30113 8480
rect 30064 8440 30070 8452
rect 30101 8449 30113 8452
rect 30147 8449 30159 8483
rect 30101 8443 30159 8449
rect 31386 8440 31392 8492
rect 31444 8440 31450 8492
rect 31573 8483 31631 8489
rect 31573 8449 31585 8483
rect 31619 8449 31631 8483
rect 31573 8443 31631 8449
rect 28736 8384 29040 8412
rect 30285 8415 30343 8421
rect 26936 8372 26942 8384
rect 27614 8304 27620 8356
rect 27672 8344 27678 8356
rect 28552 8344 28580 8384
rect 30285 8381 30297 8415
rect 30331 8412 30343 8415
rect 30558 8412 30564 8424
rect 30331 8384 30564 8412
rect 30331 8381 30343 8384
rect 30285 8375 30343 8381
rect 30558 8372 30564 8384
rect 30616 8412 30622 8424
rect 31588 8412 31616 8443
rect 30616 8384 31616 8412
rect 30616 8372 30622 8384
rect 31754 8372 31760 8424
rect 31812 8372 31818 8424
rect 32968 8421 32996 8576
rect 33045 8483 33103 8489
rect 33045 8449 33057 8483
rect 33091 8480 33103 8483
rect 33778 8480 33784 8492
rect 33091 8452 33784 8480
rect 33091 8449 33103 8452
rect 33045 8443 33103 8449
rect 33778 8440 33784 8452
rect 33836 8440 33842 8492
rect 32953 8415 33011 8421
rect 32953 8381 32965 8415
rect 32999 8381 33011 8415
rect 33318 8412 33324 8424
rect 32953 8375 33011 8381
rect 33152 8384 33324 8412
rect 29362 8344 29368 8356
rect 27672 8316 28488 8344
rect 28552 8316 29368 8344
rect 27672 8304 27678 8316
rect 23992 8248 25360 8276
rect 23992 8236 23998 8248
rect 26510 8236 26516 8288
rect 26568 8276 26574 8288
rect 28258 8276 28264 8288
rect 26568 8248 28264 8276
rect 26568 8236 26574 8248
rect 28258 8236 28264 8248
rect 28316 8236 28322 8288
rect 28350 8236 28356 8288
rect 28408 8236 28414 8288
rect 28460 8276 28488 8316
rect 29362 8304 29368 8316
rect 29420 8304 29426 8356
rect 30834 8344 30840 8356
rect 29472 8316 30840 8344
rect 28626 8276 28632 8288
rect 28460 8248 28632 8276
rect 28626 8236 28632 8248
rect 28684 8276 28690 8288
rect 29472 8276 29500 8316
rect 30834 8304 30840 8316
rect 30892 8304 30898 8356
rect 33152 8344 33180 8384
rect 33318 8372 33324 8384
rect 33376 8372 33382 8424
rect 31726 8316 33180 8344
rect 28684 8248 29500 8276
rect 28684 8236 28690 8248
rect 29546 8236 29552 8288
rect 29604 8276 29610 8288
rect 31726 8276 31754 8316
rect 33226 8304 33232 8356
rect 33284 8344 33290 8356
rect 33413 8347 33471 8353
rect 33413 8344 33425 8347
rect 33284 8316 33425 8344
rect 33284 8304 33290 8316
rect 33413 8313 33425 8316
rect 33459 8313 33471 8347
rect 33413 8307 33471 8313
rect 29604 8248 31754 8276
rect 29604 8236 29610 8248
rect 1104 8186 38272 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38272 8186
rect 1104 8112 38272 8134
rect 4982 8032 4988 8084
rect 5040 8032 5046 8084
rect 7466 8032 7472 8084
rect 7524 8032 7530 8084
rect 7926 8032 7932 8084
rect 7984 8032 7990 8084
rect 9398 8072 9404 8084
rect 8128 8044 9404 8072
rect 5000 8004 5028 8032
rect 4724 7976 5028 8004
rect 4724 7945 4752 7976
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 4982 7896 4988 7948
rect 5040 7896 5046 7948
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7936 5779 7939
rect 6086 7936 6092 7948
rect 5767 7908 6092 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 7484 7868 7512 8032
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8128 8004 8156 8044
rect 9398 8032 9404 8044
rect 9456 8072 9462 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 9456 8044 10885 8072
rect 9456 8032 9462 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 11977 8075 12035 8081
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12158 8072 12164 8084
rect 12023 8044 12164 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 12860 8044 14228 8072
rect 12860 8032 12866 8044
rect 7892 7976 8156 8004
rect 12713 8007 12771 8013
rect 7892 7964 7898 7976
rect 12713 7973 12725 8007
rect 12759 8004 12771 8007
rect 14200 8004 14228 8044
rect 14274 8032 14280 8084
rect 14332 8032 14338 8084
rect 25682 8032 25688 8084
rect 25740 8072 25746 8084
rect 26878 8072 26884 8084
rect 25740 8044 26884 8072
rect 25740 8032 25746 8044
rect 26878 8032 26884 8044
rect 26936 8032 26942 8084
rect 27154 8032 27160 8084
rect 27212 8072 27218 8084
rect 27338 8072 27344 8084
rect 27212 8044 27344 8072
rect 27212 8032 27218 8044
rect 27338 8032 27344 8044
rect 27396 8032 27402 8084
rect 28718 8072 28724 8084
rect 28368 8044 28724 8072
rect 14366 8004 14372 8016
rect 12759 7976 13768 8004
rect 14200 7976 14372 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 10689 7939 10747 7945
rect 7944 7908 10456 7936
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 4663 7840 4752 7868
rect 7484 7840 7849 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4724 7812 4752 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 4706 7760 4712 7812
rect 4764 7760 4770 7812
rect 5994 7760 6000 7812
rect 6052 7760 6058 7812
rect 7466 7800 7472 7812
rect 7222 7772 7472 7800
rect 7466 7760 7472 7772
rect 7524 7800 7530 7812
rect 7944 7800 7972 7908
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 7524 7772 7972 7800
rect 7524 7760 7530 7772
rect 8956 7732 8984 7831
rect 9214 7760 9220 7812
rect 9272 7760 9278 7812
rect 10428 7800 10456 7908
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 11514 7936 11520 7948
rect 10735 7908 11520 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7868 11023 7871
rect 11054 7868 11060 7880
rect 11011 7840 11060 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11348 7877 11376 7908
rect 11514 7896 11520 7908
rect 11572 7936 11578 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11572 7908 11897 7936
rect 11572 7896 11578 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 13044 7908 13185 7936
rect 13044 7896 13050 7908
rect 13173 7905 13185 7908
rect 13219 7905 13231 7939
rect 13173 7899 13231 7905
rect 13262 7896 13268 7948
rect 13320 7896 13326 7948
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11606 7828 11612 7880
rect 11664 7828 11670 7880
rect 13078 7828 13084 7880
rect 13136 7828 13142 7880
rect 13740 7877 13768 7976
rect 14366 7964 14372 7976
rect 14424 8004 14430 8016
rect 14424 7976 14872 8004
rect 14424 7964 14430 7976
rect 14844 7948 14872 7976
rect 19426 7964 19432 8016
rect 19484 8004 19490 8016
rect 19705 8007 19763 8013
rect 19705 8004 19717 8007
rect 19484 7976 19717 8004
rect 19484 7964 19490 7976
rect 19705 7973 19717 7976
rect 19751 7973 19763 8007
rect 19705 7967 19763 7973
rect 28368 7948 28396 8044
rect 28718 8032 28724 8044
rect 28776 8072 28782 8084
rect 28813 8075 28871 8081
rect 28813 8072 28825 8075
rect 28776 8044 28825 8072
rect 28776 8032 28782 8044
rect 28813 8041 28825 8044
rect 28859 8041 28871 8075
rect 28813 8035 28871 8041
rect 29181 8075 29239 8081
rect 29181 8041 29193 8075
rect 29227 8072 29239 8075
rect 30006 8072 30012 8084
rect 29227 8044 30012 8072
rect 29227 8041 29239 8044
rect 29181 8035 29239 8041
rect 30006 8032 30012 8044
rect 30064 8032 30070 8084
rect 31846 8032 31852 8084
rect 31904 8072 31910 8084
rect 31941 8075 31999 8081
rect 31941 8072 31953 8075
rect 31904 8044 31953 8072
rect 31904 8032 31910 8044
rect 31941 8041 31953 8044
rect 31987 8041 31999 8075
rect 31941 8035 31999 8041
rect 30558 7964 30564 8016
rect 30616 8004 30622 8016
rect 31662 8004 31668 8016
rect 30616 7976 31668 8004
rect 30616 7964 30622 7976
rect 14734 7896 14740 7948
rect 14792 7896 14798 7948
rect 14826 7896 14832 7948
rect 14884 7896 14890 7948
rect 19720 7908 20208 7936
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 14516 7840 14657 7868
rect 14516 7828 14522 7840
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 18138 7868 18144 7880
rect 17644 7840 18144 7868
rect 17644 7828 17650 7840
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 19720 7877 19748 7908
rect 20180 7880 20208 7908
rect 20530 7896 20536 7948
rect 20588 7936 20594 7948
rect 22462 7936 22468 7948
rect 20588 7908 22468 7936
rect 20588 7896 20594 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 27065 7939 27123 7945
rect 23124 7908 23520 7936
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19978 7828 19984 7880
rect 20036 7828 20042 7880
rect 20070 7828 20076 7880
rect 20128 7828 20134 7880
rect 20162 7828 20168 7880
rect 20220 7828 20226 7880
rect 23124 7868 23152 7908
rect 23492 7880 23520 7908
rect 27065 7905 27077 7939
rect 27111 7936 27123 7939
rect 28350 7936 28356 7948
rect 27111 7908 28356 7936
rect 27111 7905 27123 7908
rect 27065 7899 27123 7905
rect 28350 7896 28356 7908
rect 28408 7896 28414 7948
rect 28442 7896 28448 7948
rect 28500 7936 28506 7948
rect 30469 7939 30527 7945
rect 28500 7908 29776 7936
rect 28500 7896 28506 7908
rect 22066 7840 23152 7868
rect 23201 7871 23259 7877
rect 19889 7803 19947 7809
rect 10428 7786 12296 7800
rect 10442 7772 12296 7786
rect 12268 7744 12296 7772
rect 19889 7769 19901 7803
rect 19935 7800 19947 7803
rect 20088 7800 20116 7828
rect 19935 7772 20116 7800
rect 19935 7769 19947 7772
rect 19889 7763 19947 7769
rect 20530 7760 20536 7812
rect 20588 7800 20594 7812
rect 22066 7800 22094 7840
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 20588 7772 22094 7800
rect 23216 7800 23244 7831
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 23566 7828 23572 7880
rect 23624 7828 23630 7880
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7868 23719 7871
rect 24026 7868 24032 7880
rect 23707 7840 24032 7868
rect 23707 7837 23719 7840
rect 23661 7831 23719 7837
rect 24026 7828 24032 7840
rect 24084 7828 24090 7880
rect 25958 7828 25964 7880
rect 26016 7868 26022 7880
rect 26789 7871 26847 7877
rect 26789 7868 26801 7871
rect 26016 7840 26801 7868
rect 26016 7828 26022 7840
rect 26789 7837 26801 7840
rect 26835 7837 26847 7871
rect 26789 7831 26847 7837
rect 26970 7828 26976 7880
rect 27028 7828 27034 7880
rect 27154 7828 27160 7880
rect 27212 7828 27218 7880
rect 27341 7871 27399 7877
rect 27341 7837 27353 7871
rect 27387 7837 27399 7871
rect 27341 7831 27399 7837
rect 23584 7800 23612 7828
rect 23216 7772 23612 7800
rect 20588 7760 20594 7772
rect 27356 7744 27384 7831
rect 28166 7828 28172 7880
rect 28224 7868 28230 7880
rect 28810 7868 28816 7880
rect 28224 7840 28816 7868
rect 28224 7828 28230 7840
rect 28810 7828 28816 7840
rect 28868 7828 28874 7880
rect 28905 7871 28963 7877
rect 28905 7837 28917 7871
rect 28951 7837 28963 7871
rect 28905 7831 28963 7837
rect 27448 7772 28488 7800
rect 27448 7744 27476 7772
rect 9490 7732 9496 7744
rect 8956 7704 9496 7732
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 12158 7692 12164 7744
rect 12216 7692 12222 7744
rect 12250 7692 12256 7744
rect 12308 7692 12314 7744
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 13320 7704 13553 7732
rect 13320 7692 13326 7704
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13541 7695 13599 7701
rect 20346 7692 20352 7744
rect 20404 7732 20410 7744
rect 20622 7732 20628 7744
rect 20404 7704 20628 7732
rect 20404 7692 20410 7704
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 23014 7692 23020 7744
rect 23072 7692 23078 7744
rect 27338 7692 27344 7744
rect 27396 7692 27402 7744
rect 27430 7692 27436 7744
rect 27488 7692 27494 7744
rect 27522 7692 27528 7744
rect 27580 7692 27586 7744
rect 28460 7732 28488 7772
rect 28534 7760 28540 7812
rect 28592 7800 28598 7812
rect 28920 7800 28948 7831
rect 29546 7828 29552 7880
rect 29604 7828 29610 7880
rect 29748 7877 29776 7908
rect 30469 7905 30481 7939
rect 30515 7936 30527 7939
rect 30515 7908 30696 7936
rect 30515 7905 30527 7908
rect 30469 7899 30527 7905
rect 30668 7880 30696 7908
rect 30760 7908 31340 7936
rect 29733 7871 29791 7877
rect 29733 7837 29745 7871
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 30193 7871 30251 7877
rect 30193 7837 30205 7871
rect 30239 7837 30251 7871
rect 30193 7831 30251 7837
rect 28592 7772 28948 7800
rect 28592 7760 28598 7772
rect 29564 7732 29592 7828
rect 29641 7803 29699 7809
rect 29641 7769 29653 7803
rect 29687 7800 29699 7803
rect 30208 7800 30236 7831
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 30377 7871 30435 7877
rect 30377 7868 30389 7871
rect 30340 7840 30389 7868
rect 30340 7828 30346 7840
rect 30377 7837 30389 7840
rect 30423 7837 30435 7871
rect 30377 7831 30435 7837
rect 30558 7828 30564 7880
rect 30616 7828 30622 7880
rect 30650 7828 30656 7880
rect 30708 7828 30714 7880
rect 30760 7877 30788 7908
rect 31312 7880 31340 7908
rect 30745 7871 30803 7877
rect 30745 7837 30757 7871
rect 30791 7837 30803 7871
rect 30745 7831 30803 7837
rect 30834 7828 30840 7880
rect 30892 7868 30898 7880
rect 31021 7871 31079 7877
rect 31021 7868 31033 7871
rect 30892 7840 31033 7868
rect 30892 7828 30898 7840
rect 31021 7837 31033 7840
rect 31067 7837 31079 7871
rect 31021 7831 31079 7837
rect 31294 7828 31300 7880
rect 31352 7828 31358 7880
rect 31404 7877 31432 7976
rect 31662 7964 31668 7976
rect 31720 7964 31726 8016
rect 31754 7936 31760 7948
rect 31588 7908 31760 7936
rect 31588 7877 31616 7908
rect 31754 7896 31760 7908
rect 31812 7896 31818 7948
rect 31389 7871 31447 7877
rect 31389 7837 31401 7871
rect 31435 7837 31447 7871
rect 31389 7831 31447 7837
rect 31481 7871 31539 7877
rect 31481 7837 31493 7871
rect 31527 7868 31539 7871
rect 31573 7871 31631 7877
rect 31573 7868 31585 7871
rect 31527 7840 31585 7868
rect 31527 7837 31539 7840
rect 31481 7831 31539 7837
rect 31573 7837 31585 7840
rect 31619 7837 31631 7871
rect 31573 7831 31631 7837
rect 29687 7772 30236 7800
rect 30944 7772 31524 7800
rect 29687 7769 29699 7772
rect 29641 7763 29699 7769
rect 30944 7741 30972 7772
rect 31496 7744 31524 7772
rect 31662 7760 31668 7812
rect 31720 7800 31726 7812
rect 31757 7803 31815 7809
rect 31757 7800 31769 7803
rect 31720 7772 31769 7800
rect 31720 7760 31726 7772
rect 31757 7769 31769 7772
rect 31803 7769 31815 7803
rect 31757 7763 31815 7769
rect 28460 7704 29592 7732
rect 30929 7735 30987 7741
rect 30929 7701 30941 7735
rect 30975 7701 30987 7735
rect 30929 7695 30987 7701
rect 31294 7692 31300 7744
rect 31352 7692 31358 7744
rect 31478 7692 31484 7744
rect 31536 7692 31542 7744
rect 1104 7642 38272 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38272 7642
rect 1104 7568 38272 7590
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4479 7500 4905 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4893 7497 4905 7500
rect 4939 7497 4951 7531
rect 4893 7491 4951 7497
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5040 7500 5365 7528
rect 5040 7488 5046 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6052 7500 6377 7528
rect 6052 7488 6058 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6638 7488 6644 7540
rect 6696 7488 6702 7540
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 9272 7500 9321 7528
rect 9272 7488 9278 7500
rect 9309 7497 9321 7500
rect 9355 7497 9367 7531
rect 9309 7491 9367 7497
rect 13262 7488 13268 7540
rect 13320 7488 13326 7540
rect 15286 7488 15292 7540
rect 15344 7488 15350 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 17236 7500 17693 7528
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4706 7392 4712 7404
rect 4387 7364 4712 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 5258 7352 5264 7404
rect 5316 7352 5322 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 6656 7392 6684 7488
rect 10134 7460 10140 7472
rect 9232 7432 10140 7460
rect 9232 7401 9260 7432
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7460 13047 7463
rect 13280 7460 13308 7488
rect 14274 7460 14280 7472
rect 13035 7432 13308 7460
rect 14214 7432 14280 7460
rect 13035 7429 13047 7432
rect 12989 7423 13047 7429
rect 14274 7420 14280 7432
rect 14332 7460 14338 7472
rect 15102 7460 15108 7472
rect 14332 7432 15108 7460
rect 14332 7420 14338 7432
rect 15102 7420 15108 7432
rect 15160 7420 15166 7472
rect 17236 7469 17264 7500
rect 17681 7497 17693 7500
rect 17727 7497 17739 7531
rect 17681 7491 17739 7497
rect 19426 7488 19432 7540
rect 19484 7488 19490 7540
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 19944 7500 20484 7528
rect 19944 7488 19950 7500
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7429 17279 7463
rect 17221 7423 17279 7429
rect 6595 7364 6684 7392
rect 9217 7395 9275 7401
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9398 7352 9404 7404
rect 9456 7352 9462 7404
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 11606 7352 11612 7404
rect 11664 7352 11670 7404
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7392 15439 7395
rect 17034 7392 17040 7404
rect 15427 7364 17040 7392
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17586 7392 17592 7404
rect 17543 7364 17592 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7361 17831 7395
rect 19444 7392 19472 7488
rect 19613 7463 19671 7469
rect 19613 7429 19625 7463
rect 19659 7460 19671 7463
rect 20456 7460 20484 7500
rect 20530 7488 20536 7540
rect 20588 7488 20594 7540
rect 22370 7528 22376 7540
rect 20824 7500 22376 7528
rect 20824 7460 20852 7500
rect 22370 7488 22376 7500
rect 22428 7528 22434 7540
rect 22738 7528 22744 7540
rect 22428 7500 22744 7528
rect 22428 7488 22434 7500
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 23014 7488 23020 7540
rect 23072 7488 23078 7540
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 26789 7531 26847 7537
rect 24412 7500 26740 7528
rect 19659 7432 20392 7460
rect 20456 7432 20852 7460
rect 19659 7429 19671 7432
rect 19613 7423 19671 7429
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19444 7364 19533 7392
rect 17773 7355 17831 7361
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7392 19763 7395
rect 19886 7392 19892 7404
rect 19751 7364 19892 7392
rect 19751 7361 19763 7364
rect 19705 7355 19763 7361
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 5074 7324 5080 7336
rect 4672 7296 5080 7324
rect 4672 7284 4678 7296
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5224 7296 5457 7324
rect 5224 7284 5230 7296
rect 5445 7293 5457 7296
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 9548 7296 9597 7324
rect 9548 7284 9554 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7324 9919 7327
rect 11333 7327 11391 7333
rect 9907 7296 11100 7324
rect 9907 7293 9919 7296
rect 9861 7287 9919 7293
rect 11072 7268 11100 7296
rect 11333 7293 11345 7327
rect 11379 7324 11391 7327
rect 11624 7324 11652 7352
rect 11379 7296 11652 7324
rect 11379 7293 11391 7296
rect 11333 7287 11391 7293
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 12342 7324 12348 7336
rect 11756 7296 12348 7324
rect 11756 7284 11762 7296
rect 12342 7284 12348 7296
rect 12400 7324 12406 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12400 7296 12725 7324
rect 12400 7284 12406 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 14737 7327 14795 7333
rect 14737 7324 14749 7327
rect 13044 7296 14749 7324
rect 13044 7284 13050 7296
rect 14737 7293 14749 7296
rect 14783 7293 14795 7327
rect 14737 7287 14795 7293
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 14884 7296 15485 7324
rect 14884 7284 14890 7296
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 17052 7324 17080 7352
rect 17788 7324 17816 7355
rect 17052 7296 17816 7324
rect 19536 7324 19564 7355
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 19981 7395 20039 7401
rect 19981 7361 19993 7395
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 19996 7324 20024 7355
rect 20162 7352 20168 7404
rect 20220 7352 20226 7404
rect 20254 7352 20260 7404
rect 20312 7352 20318 7404
rect 20364 7401 20392 7432
rect 20824 7401 20852 7432
rect 21634 7420 21640 7472
rect 21692 7460 21698 7472
rect 21692 7432 22232 7460
rect 21692 7420 21698 7432
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 20533 7395 20591 7401
rect 20533 7361 20545 7395
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 19536 7296 20024 7324
rect 15473 7287 15531 7293
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 9306 7256 9312 7268
rect 1719 7228 9312 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 11054 7216 11060 7268
rect 11112 7216 11118 7268
rect 14274 7216 14280 7268
rect 14332 7216 14338 7268
rect 19797 7259 19855 7265
rect 19797 7225 19809 7259
rect 19843 7256 19855 7259
rect 20346 7256 20352 7268
rect 19843 7228 20352 7256
rect 19843 7225 19855 7228
rect 19797 7219 19855 7225
rect 20346 7216 20352 7228
rect 20404 7256 20410 7268
rect 20548 7256 20576 7355
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22204 7392 22232 7432
rect 22922 7420 22928 7472
rect 22980 7420 22986 7472
rect 22327 7395 22385 7401
rect 22327 7392 22339 7395
rect 22204 7364 22339 7392
rect 22327 7361 22339 7364
rect 22373 7361 22385 7395
rect 22327 7355 22385 7361
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7392 22891 7395
rect 23032 7392 23060 7488
rect 22879 7364 23060 7392
rect 23492 7392 23520 7488
rect 24029 7463 24087 7469
rect 24029 7429 24041 7463
rect 24075 7460 24087 7463
rect 24075 7432 24256 7460
rect 24075 7429 24087 7432
rect 24029 7423 24087 7429
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23492 7364 23949 7392
rect 22879 7361 22891 7364
rect 22833 7355 22891 7361
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24228 7401 24256 7432
rect 24412 7401 24440 7500
rect 26712 7472 26740 7500
rect 26789 7497 26801 7531
rect 26835 7528 26847 7531
rect 27338 7528 27344 7540
rect 26835 7500 27344 7528
rect 26835 7497 26847 7500
rect 26789 7491 26847 7497
rect 27338 7488 27344 7500
rect 27396 7528 27402 7540
rect 27396 7500 27476 7528
rect 27396 7488 27402 7500
rect 24946 7420 24952 7472
rect 25004 7460 25010 7472
rect 25041 7463 25099 7469
rect 25041 7460 25053 7463
rect 25004 7432 25053 7460
rect 25004 7420 25010 7432
rect 25041 7429 25053 7432
rect 25087 7429 25099 7463
rect 25869 7463 25927 7469
rect 25869 7460 25881 7463
rect 25041 7423 25099 7429
rect 25516 7432 25881 7460
rect 24213 7395 24271 7401
rect 24213 7361 24225 7395
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 24578 7352 24584 7404
rect 24636 7352 24642 7404
rect 24762 7352 24768 7404
rect 24820 7352 24826 7404
rect 25516 7401 25544 7432
rect 25869 7429 25881 7432
rect 25915 7429 25927 7463
rect 25869 7423 25927 7429
rect 26510 7420 26516 7472
rect 26568 7420 26574 7472
rect 26694 7420 26700 7472
rect 26752 7420 26758 7472
rect 26878 7460 26884 7472
rect 26804 7432 26884 7460
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 25777 7395 25835 7401
rect 25777 7361 25789 7395
rect 25823 7361 25835 7395
rect 25777 7355 25835 7361
rect 25961 7395 26019 7401
rect 25961 7361 25973 7395
rect 26007 7361 26019 7395
rect 26528 7390 26556 7420
rect 26804 7401 26832 7432
rect 26878 7420 26884 7432
rect 26936 7420 26942 7472
rect 26789 7395 26847 7401
rect 26605 7390 26663 7391
rect 26528 7385 26663 7390
rect 26528 7362 26617 7385
rect 25961 7355 26019 7361
rect 20901 7327 20959 7333
rect 20901 7293 20913 7327
rect 20947 7324 20959 7327
rect 21358 7324 21364 7336
rect 20947 7296 21364 7324
rect 20947 7293 20959 7296
rect 20901 7287 20959 7293
rect 21358 7284 21364 7296
rect 21416 7324 21422 7336
rect 21726 7324 21732 7336
rect 21416 7296 21732 7324
rect 21416 7284 21422 7296
rect 21726 7284 21732 7296
rect 21784 7284 21790 7336
rect 21821 7327 21879 7333
rect 21821 7293 21833 7327
rect 21867 7324 21879 7327
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 21867 7296 22753 7324
rect 21867 7293 21879 7296
rect 21821 7287 21879 7293
rect 22741 7293 22753 7296
rect 22787 7293 22799 7327
rect 22741 7287 22799 7293
rect 23106 7284 23112 7336
rect 23164 7324 23170 7336
rect 24489 7327 24547 7333
rect 24489 7324 24501 7327
rect 23164 7296 24501 7324
rect 23164 7284 23170 7296
rect 24489 7293 24501 7296
rect 24535 7293 24547 7327
rect 24489 7287 24547 7293
rect 25409 7327 25467 7333
rect 25409 7293 25421 7327
rect 25455 7324 25467 7327
rect 25590 7324 25596 7336
rect 25455 7296 25596 7324
rect 25455 7293 25467 7296
rect 25409 7287 25467 7293
rect 25590 7284 25596 7296
rect 25648 7284 25654 7336
rect 20404 7228 20576 7256
rect 20404 7216 20410 7228
rect 21174 7216 21180 7268
rect 21232 7216 21238 7268
rect 22557 7259 22615 7265
rect 22557 7225 22569 7259
rect 22603 7256 22615 7259
rect 23658 7256 23664 7268
rect 22603 7228 23664 7256
rect 22603 7225 22615 7228
rect 22557 7219 22615 7225
rect 23658 7216 23664 7228
rect 23716 7216 23722 7268
rect 25792 7256 25820 7355
rect 24872 7228 25820 7256
rect 25976 7256 26004 7355
rect 26605 7351 26617 7362
rect 26651 7351 26663 7385
rect 26789 7361 26801 7395
rect 26835 7361 26847 7395
rect 26789 7355 26847 7361
rect 27246 7352 27252 7404
rect 27304 7352 27310 7404
rect 27338 7352 27344 7404
rect 27396 7352 27402 7404
rect 27448 7401 27476 7500
rect 31294 7488 31300 7540
rect 31352 7488 31358 7540
rect 31478 7488 31484 7540
rect 31536 7528 31542 7540
rect 31536 7500 33364 7528
rect 31536 7488 31542 7500
rect 28166 7460 28172 7472
rect 27540 7432 28172 7460
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 26605 7345 26663 7351
rect 26973 7327 27031 7333
rect 26973 7293 26985 7327
rect 27019 7324 27031 7327
rect 27540 7324 27568 7432
rect 28166 7420 28172 7432
rect 28224 7420 28230 7472
rect 30745 7463 30803 7469
rect 29196 7432 30328 7460
rect 27617 7395 27675 7401
rect 27617 7361 27629 7395
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 27019 7296 27568 7324
rect 27019 7293 27031 7296
rect 26973 7287 27031 7293
rect 26418 7256 26424 7268
rect 25976 7228 26424 7256
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 3973 7191 4031 7197
rect 3973 7188 3985 7191
rect 3752 7160 3985 7188
rect 3752 7148 3758 7160
rect 3973 7157 3985 7160
rect 4019 7157 4031 7191
rect 3973 7151 4031 7157
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 11480 7160 12173 7188
rect 11480 7148 11486 7160
rect 12161 7157 12173 7160
rect 12207 7157 12219 7191
rect 12161 7151 12219 7157
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 14292 7188 14320 7216
rect 12308 7160 14320 7188
rect 14921 7191 14979 7197
rect 12308 7148 12314 7160
rect 14921 7157 14933 7191
rect 14967 7188 14979 7191
rect 15194 7188 15200 7200
rect 14967 7160 15200 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 17218 7148 17224 7200
rect 17276 7148 17282 7200
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 20162 7188 20168 7200
rect 19392 7160 20168 7188
rect 19392 7148 19398 7160
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 22281 7191 22339 7197
rect 22281 7188 22293 7191
rect 20772 7160 22293 7188
rect 20772 7148 20778 7160
rect 22281 7157 22293 7160
rect 22327 7188 22339 7191
rect 24872 7188 24900 7228
rect 22327 7160 24900 7188
rect 22327 7157 22339 7160
rect 22281 7151 22339 7157
rect 24946 7148 24952 7200
rect 25004 7148 25010 7200
rect 25130 7148 25136 7200
rect 25188 7148 25194 7200
rect 25682 7148 25688 7200
rect 25740 7148 25746 7200
rect 25792 7188 25820 7228
rect 26418 7216 26424 7228
rect 26476 7256 26482 7268
rect 27632 7256 27660 7355
rect 28442 7352 28448 7404
rect 28500 7352 28506 7404
rect 29196 7401 29224 7432
rect 30300 7404 30328 7432
rect 30745 7429 30757 7463
rect 30791 7460 30803 7463
rect 31018 7460 31024 7472
rect 30791 7432 31024 7460
rect 30791 7429 30803 7432
rect 30745 7423 30803 7429
rect 31018 7420 31024 7432
rect 31076 7420 31082 7472
rect 31312 7460 31340 7488
rect 31312 7432 31984 7460
rect 29181 7395 29239 7401
rect 29181 7361 29193 7395
rect 29227 7361 29239 7395
rect 29181 7355 29239 7361
rect 29270 7352 29276 7404
rect 29328 7352 29334 7404
rect 29362 7352 29368 7404
rect 29420 7392 29426 7404
rect 29549 7395 29607 7401
rect 29549 7392 29561 7395
rect 29420 7364 29561 7392
rect 29420 7352 29426 7364
rect 29549 7361 29561 7364
rect 29595 7361 29607 7395
rect 29549 7355 29607 7361
rect 29825 7395 29883 7401
rect 29825 7361 29837 7395
rect 29871 7361 29883 7395
rect 29825 7355 29883 7361
rect 29086 7284 29092 7336
rect 29144 7284 29150 7336
rect 26476 7228 27660 7256
rect 29840 7256 29868 7355
rect 30282 7352 30288 7404
rect 30340 7352 30346 7404
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7392 31447 7395
rect 31757 7395 31815 7401
rect 31846 7395 31852 7404
rect 31435 7364 31616 7392
rect 31435 7361 31447 7364
rect 31389 7355 31447 7361
rect 31294 7284 31300 7336
rect 31352 7284 31358 7336
rect 31588 7324 31616 7364
rect 31757 7361 31769 7395
rect 31803 7367 31852 7395
rect 31803 7361 31815 7367
rect 31757 7355 31815 7361
rect 31846 7352 31852 7367
rect 31904 7352 31910 7404
rect 31956 7401 31984 7432
rect 33336 7401 33364 7500
rect 33686 7488 33692 7540
rect 33744 7488 33750 7540
rect 31941 7395 31999 7401
rect 31941 7361 31953 7395
rect 31987 7361 31999 7395
rect 31941 7355 31999 7361
rect 33321 7395 33379 7401
rect 33321 7361 33333 7395
rect 33367 7361 33379 7395
rect 33321 7355 33379 7361
rect 32122 7324 32128 7336
rect 31588 7296 32128 7324
rect 32122 7284 32128 7296
rect 32180 7284 32186 7336
rect 33229 7327 33287 7333
rect 33229 7293 33241 7327
rect 33275 7293 33287 7327
rect 33229 7287 33287 7293
rect 33244 7256 33272 7287
rect 33318 7256 33324 7268
rect 29840 7228 33180 7256
rect 33244 7228 33324 7256
rect 26476 7216 26482 7228
rect 27154 7188 27160 7200
rect 25792 7160 27160 7188
rect 27154 7148 27160 7160
rect 27212 7148 27218 7200
rect 29362 7148 29368 7200
rect 29420 7188 29426 7200
rect 31754 7188 31760 7200
rect 29420 7160 31760 7188
rect 29420 7148 29426 7160
rect 31754 7148 31760 7160
rect 31812 7148 31818 7200
rect 33152 7188 33180 7228
rect 33318 7216 33324 7228
rect 33376 7216 33382 7268
rect 34054 7188 34060 7200
rect 33152 7160 34060 7188
rect 34054 7148 34060 7160
rect 34112 7148 34118 7200
rect 1104 7098 38272 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38272 7098
rect 1104 7024 38272 7046
rect 5258 6944 5264 6996
rect 5316 6984 5322 6996
rect 5316 6956 11008 6984
rect 5316 6944 5322 6956
rect 5074 6876 5080 6928
rect 5132 6916 5138 6928
rect 10980 6916 11008 6956
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11241 6987 11299 6993
rect 11241 6984 11253 6987
rect 11112 6956 11253 6984
rect 11112 6944 11118 6956
rect 11241 6953 11253 6956
rect 11287 6953 11299 6987
rect 11241 6947 11299 6953
rect 11514 6944 11520 6996
rect 11572 6944 11578 6996
rect 17218 6984 17224 6996
rect 12406 6956 17224 6984
rect 12406 6916 12434 6956
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 17773 6987 17831 6993
rect 17773 6984 17785 6987
rect 17460 6956 17785 6984
rect 17460 6944 17466 6956
rect 17773 6953 17785 6956
rect 17819 6984 17831 6987
rect 18598 6984 18604 6996
rect 17819 6956 18604 6984
rect 17819 6953 17831 6956
rect 17773 6947 17831 6953
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 19886 6944 19892 6996
rect 19944 6984 19950 6996
rect 20070 6984 20076 6996
rect 19944 6956 20076 6984
rect 19944 6944 19950 6956
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 20162 6944 20168 6996
rect 20220 6984 20226 6996
rect 21634 6984 21640 6996
rect 20220 6956 21640 6984
rect 20220 6944 20226 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22462 6944 22468 6996
rect 22520 6984 22526 6996
rect 23934 6984 23940 6996
rect 22520 6956 23940 6984
rect 22520 6944 22526 6956
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 25590 6944 25596 6996
rect 25648 6944 25654 6996
rect 27522 6944 27528 6996
rect 27580 6944 27586 6996
rect 28258 6944 28264 6996
rect 28316 6984 28322 6996
rect 29914 6984 29920 6996
rect 28316 6956 29920 6984
rect 28316 6944 28322 6956
rect 29914 6944 29920 6956
rect 29972 6944 29978 6996
rect 31294 6944 31300 6996
rect 31352 6944 31358 6996
rect 33134 6944 33140 6996
rect 33192 6944 33198 6996
rect 5132 6888 6316 6916
rect 5132 6876 5138 6888
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 6178 6848 6184 6860
rect 3835 6820 6184 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6288 6848 6316 6888
rect 8036 6888 8708 6916
rect 10980 6888 12434 6916
rect 7190 6848 7196 6860
rect 6288 6820 7196 6848
rect 7190 6808 7196 6820
rect 7248 6848 7254 6860
rect 8036 6848 8064 6888
rect 7248 6820 8064 6848
rect 7248 6808 7254 6820
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 8168 6820 8493 6848
rect 8168 6808 8174 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 8570 6808 8576 6860
rect 8628 6808 8634 6860
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3694 6780 3700 6792
rect 3651 6752 3700 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7524 6766 7590 6780
rect 7524 6752 7604 6766
rect 7524 6740 7530 6752
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 3436 6684 4077 6712
rect 3436 6653 3464 6684
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 5290 6684 5764 6712
rect 4065 6675 4123 6681
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 4764 6616 5549 6644
rect 4764 6604 4770 6616
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5736 6644 5764 6684
rect 6454 6672 6460 6724
rect 6512 6672 6518 6724
rect 7576 6644 7604 6752
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8202 6780 8208 6792
rect 7984 6752 8208 6780
rect 7984 6740 7990 6752
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8294 6712 8300 6724
rect 7944 6684 8300 6712
rect 7944 6653 7972 6684
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 8680 6712 8708 6888
rect 17034 6876 17040 6928
rect 17092 6916 17098 6928
rect 17586 6916 17592 6928
rect 17092 6888 17592 6916
rect 17092 6876 17098 6888
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 18141 6919 18199 6925
rect 18141 6885 18153 6919
rect 18187 6916 18199 6919
rect 20254 6916 20260 6928
rect 18187 6888 20260 6916
rect 18187 6885 18199 6888
rect 18141 6879 18199 6885
rect 11256 6820 11560 6848
rect 11256 6789 11284 6820
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 11532 6789 11560 6820
rect 11606 6808 11612 6860
rect 11664 6808 11670 6860
rect 17497 6851 17555 6857
rect 17497 6817 17509 6851
rect 17543 6848 17555 6851
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17543 6820 17969 6848
rect 17543 6817 17555 6820
rect 17497 6811 17555 6817
rect 17957 6817 17969 6820
rect 18003 6848 18015 6851
rect 18414 6848 18420 6860
rect 18003 6820 18420 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 18414 6808 18420 6820
rect 18472 6848 18478 6860
rect 19245 6851 19303 6857
rect 18472 6820 18736 6848
rect 18472 6808 18478 6820
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 12066 6780 12072 6792
rect 11563 6752 12072 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 13170 6740 13176 6792
rect 13228 6740 13234 6792
rect 15194 6740 15200 6792
rect 15252 6740 15258 6792
rect 15286 6740 15292 6792
rect 15344 6740 15350 6792
rect 17405 6773 17463 6779
rect 17405 6739 17417 6773
rect 17451 6770 17463 6773
rect 17451 6742 17540 6770
rect 17451 6739 17463 6742
rect 17405 6733 17463 6739
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 8680 6684 12112 6712
rect 5736 6616 7604 6644
rect 7929 6647 7987 6653
rect 5537 6607 5595 6613
rect 7929 6613 7941 6647
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8018 6604 8024 6656
rect 8076 6604 8082 6656
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 11238 6644 11244 6656
rect 10468 6616 11244 6644
rect 10468 6604 10474 6616
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11882 6604 11888 6656
rect 11940 6604 11946 6656
rect 12084 6653 12112 6684
rect 15028 6684 15577 6712
rect 15028 6653 15056 6684
rect 15565 6681 15577 6684
rect 15611 6681 15623 6715
rect 15565 6675 15623 6681
rect 16574 6672 16580 6724
rect 16632 6672 16638 6724
rect 17512 6712 17540 6742
rect 17586 6740 17592 6792
rect 17644 6740 17650 6792
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 17727 6752 17828 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 17800 6712 17828 6752
rect 18046 6740 18052 6792
rect 18104 6740 18110 6792
rect 18506 6780 18512 6792
rect 18156 6752 18512 6780
rect 18156 6712 18184 6752
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18598 6740 18604 6792
rect 18656 6740 18662 6792
rect 18708 6789 18736 6820
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 19334 6848 19340 6860
rect 19291 6820 19340 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 19444 6789 19472 6888
rect 20254 6876 20260 6888
rect 20312 6876 20318 6928
rect 21726 6876 21732 6928
rect 21784 6876 21790 6928
rect 22278 6876 22284 6928
rect 22336 6916 22342 6928
rect 23661 6919 23719 6925
rect 22336 6888 23336 6916
rect 22336 6876 22342 6888
rect 22094 6848 22100 6860
rect 19536 6820 22100 6848
rect 18877 6783 18935 6789
rect 18877 6780 18889 6783
rect 18840 6752 18889 6780
rect 18840 6740 18846 6752
rect 18877 6749 18889 6752
rect 18923 6749 18935 6783
rect 18877 6743 18935 6749
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 17512 6684 17828 6712
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6613 15071 6647
rect 17800 6644 17828 6684
rect 17972 6684 18184 6712
rect 18233 6715 18291 6721
rect 17972 6644 18000 6684
rect 18233 6681 18245 6715
rect 18279 6712 18291 6715
rect 19536 6712 19564 6820
rect 21174 6740 21180 6792
rect 21232 6740 21238 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 21634 6780 21640 6792
rect 21591 6752 21640 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 21836 6789 21864 6820
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 23106 6848 23112 6860
rect 22296 6820 23112 6848
rect 21821 6783 21879 6789
rect 21821 6749 21833 6783
rect 21867 6749 21879 6783
rect 21821 6743 21879 6749
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 21968 6752 22201 6780
rect 21968 6740 21974 6752
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 18279 6684 19564 6712
rect 19613 6715 19671 6721
rect 18279 6681 18291 6684
rect 18233 6675 18291 6681
rect 19613 6681 19625 6715
rect 19659 6712 19671 6715
rect 19981 6715 20039 6721
rect 19981 6712 19993 6715
rect 19659 6684 19993 6712
rect 19659 6681 19671 6684
rect 19613 6675 19671 6681
rect 19981 6681 19993 6684
rect 20027 6681 20039 6715
rect 21192 6712 21220 6740
rect 22005 6715 22063 6721
rect 22005 6712 22017 6715
rect 21192 6684 22017 6712
rect 19981 6675 20039 6681
rect 22005 6681 22017 6684
rect 22051 6712 22063 6715
rect 22296 6712 22324 6820
rect 23106 6808 23112 6820
rect 23164 6808 23170 6860
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6780 22431 6783
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 22419 6752 22477 6780
rect 22419 6749 22431 6752
rect 22373 6743 22431 6749
rect 22465 6749 22477 6752
rect 22511 6749 22523 6783
rect 22741 6783 22799 6789
rect 22741 6780 22753 6783
rect 22465 6743 22523 6749
rect 22572 6752 22753 6780
rect 22051 6684 22324 6712
rect 22051 6681 22063 6684
rect 22005 6675 22063 6681
rect 22572 6656 22600 6752
rect 22741 6749 22753 6752
rect 22787 6749 22799 6783
rect 22741 6743 22799 6749
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6749 22891 6783
rect 22833 6743 22891 6749
rect 22848 6656 22876 6743
rect 23198 6672 23204 6724
rect 23256 6672 23262 6724
rect 23308 6712 23336 6888
rect 23661 6885 23673 6919
rect 23707 6916 23719 6919
rect 23842 6916 23848 6928
rect 23707 6888 23848 6916
rect 23707 6885 23719 6888
rect 23661 6879 23719 6885
rect 23842 6876 23848 6888
rect 23900 6876 23906 6928
rect 27246 6876 27252 6928
rect 27304 6876 27310 6928
rect 24946 6808 24952 6860
rect 25004 6848 25010 6860
rect 25041 6851 25099 6857
rect 25041 6848 25053 6851
rect 25004 6820 25053 6848
rect 25004 6808 25010 6820
rect 25041 6817 25053 6820
rect 25087 6817 25099 6851
rect 27264 6848 27292 6876
rect 25041 6811 25099 6817
rect 25608 6820 27292 6848
rect 27433 6851 27491 6857
rect 25130 6740 25136 6792
rect 25188 6740 25194 6792
rect 25498 6740 25504 6792
rect 25556 6780 25562 6792
rect 25608 6789 25636 6820
rect 27433 6817 27445 6851
rect 27479 6848 27491 6851
rect 27540 6848 27568 6944
rect 27798 6916 27804 6928
rect 27479 6820 27568 6848
rect 27632 6888 27804 6916
rect 27479 6817 27491 6820
rect 27433 6811 27491 6817
rect 25593 6783 25651 6789
rect 25593 6780 25605 6783
rect 25556 6752 25605 6780
rect 25556 6740 25562 6752
rect 25593 6749 25605 6752
rect 25639 6749 25651 6783
rect 25869 6783 25927 6789
rect 25869 6780 25881 6783
rect 25593 6743 25651 6749
rect 25700 6752 25881 6780
rect 25700 6712 25728 6752
rect 25869 6749 25881 6752
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 27062 6740 27068 6792
rect 27120 6780 27126 6792
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 27120 6752 27169 6780
rect 27120 6740 27126 6752
rect 27157 6749 27169 6752
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 27249 6783 27307 6789
rect 27249 6749 27261 6783
rect 27295 6780 27307 6783
rect 27632 6780 27660 6888
rect 27798 6876 27804 6888
rect 27856 6876 27862 6928
rect 27982 6876 27988 6928
rect 28040 6916 28046 6928
rect 28537 6919 28595 6925
rect 28537 6916 28549 6919
rect 28040 6888 28549 6916
rect 28040 6876 28046 6888
rect 28537 6885 28549 6888
rect 28583 6885 28595 6919
rect 28537 6879 28595 6885
rect 30929 6919 30987 6925
rect 30929 6885 30941 6919
rect 30975 6916 30987 6919
rect 31312 6916 31340 6944
rect 30975 6888 31340 6916
rect 32784 6888 33272 6916
rect 30975 6885 30987 6888
rect 30929 6879 30987 6885
rect 29270 6848 29276 6860
rect 28000 6820 29276 6848
rect 27890 6789 27896 6792
rect 27295 6752 27660 6780
rect 27709 6783 27767 6789
rect 27295 6749 27307 6752
rect 27249 6743 27307 6749
rect 27709 6749 27721 6783
rect 27755 6749 27767 6783
rect 27709 6743 27767 6749
rect 27857 6783 27896 6789
rect 27857 6749 27869 6783
rect 27857 6743 27896 6749
rect 23308 6684 25728 6712
rect 25777 6715 25835 6721
rect 25777 6681 25789 6715
rect 25823 6712 25835 6715
rect 27264 6712 27292 6743
rect 25823 6684 27292 6712
rect 27433 6715 27491 6721
rect 25823 6681 25835 6684
rect 25777 6675 25835 6681
rect 27433 6681 27445 6715
rect 27479 6712 27491 6715
rect 27724 6712 27752 6743
rect 27890 6740 27896 6743
rect 27948 6740 27954 6792
rect 28000 6789 28028 6820
rect 29270 6808 29276 6820
rect 29328 6808 29334 6860
rect 30466 6808 30472 6860
rect 30524 6808 30530 6860
rect 30576 6820 31064 6848
rect 30576 6792 30604 6820
rect 27985 6783 28043 6789
rect 27985 6749 27997 6783
rect 28031 6749 28043 6783
rect 27985 6743 28043 6749
rect 28166 6740 28172 6792
rect 28224 6789 28230 6792
rect 28224 6743 28232 6789
rect 28350 6780 28356 6792
rect 28276 6752 28356 6780
rect 28224 6740 28230 6743
rect 27479 6684 27752 6712
rect 28077 6715 28135 6721
rect 27479 6681 27491 6684
rect 27433 6675 27491 6681
rect 28077 6681 28089 6715
rect 28123 6712 28135 6715
rect 28276 6712 28304 6752
rect 28350 6740 28356 6752
rect 28408 6740 28414 6792
rect 28442 6740 28448 6792
rect 28500 6780 28506 6792
rect 28721 6783 28779 6789
rect 28721 6780 28733 6783
rect 28500 6752 28733 6780
rect 28500 6740 28506 6752
rect 28721 6749 28733 6752
rect 28767 6749 28779 6783
rect 28721 6743 28779 6749
rect 28905 6783 28963 6789
rect 28905 6749 28917 6783
rect 28951 6749 28963 6783
rect 28905 6743 28963 6749
rect 28997 6783 29055 6789
rect 28997 6749 29009 6783
rect 29043 6749 29055 6783
rect 28997 6743 29055 6749
rect 28920 6712 28948 6743
rect 28123 6684 28304 6712
rect 28368 6684 28948 6712
rect 28123 6681 28135 6684
rect 28077 6675 28135 6681
rect 17800 6616 18000 6644
rect 15013 6607 15071 6613
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18690 6644 18696 6656
rect 18104 6616 18696 6644
rect 18104 6604 18110 6616
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 21358 6604 21364 6656
rect 21416 6604 21422 6656
rect 22554 6604 22560 6656
rect 22612 6604 22618 6656
rect 22830 6604 22836 6656
rect 22888 6604 22894 6656
rect 25501 6647 25559 6653
rect 25501 6613 25513 6647
rect 25547 6644 25559 6647
rect 25590 6644 25596 6656
rect 25547 6616 25596 6644
rect 25547 6613 25559 6616
rect 25501 6607 25559 6613
rect 25590 6604 25596 6616
rect 25648 6604 25654 6656
rect 28368 6653 28396 6684
rect 28353 6647 28411 6653
rect 28353 6613 28365 6647
rect 28399 6613 28411 6647
rect 28353 6607 28411 6613
rect 28626 6604 28632 6656
rect 28684 6644 28690 6656
rect 29012 6644 29040 6743
rect 29178 6740 29184 6792
rect 29236 6780 29242 6792
rect 30193 6783 30251 6789
rect 30193 6780 30205 6783
rect 29236 6752 30205 6780
rect 29236 6740 29242 6752
rect 30193 6749 30205 6752
rect 30239 6749 30251 6783
rect 30193 6743 30251 6749
rect 30558 6740 30564 6792
rect 30616 6740 30622 6792
rect 30650 6740 30656 6792
rect 30708 6740 30714 6792
rect 31036 6789 31064 6820
rect 31202 6808 31208 6860
rect 31260 6808 31266 6860
rect 32490 6808 32496 6860
rect 32548 6808 32554 6860
rect 32784 6857 32812 6888
rect 32769 6851 32827 6857
rect 32769 6848 32781 6851
rect 32600 6820 32781 6848
rect 31021 6783 31079 6789
rect 31021 6749 31033 6783
rect 31067 6749 31079 6783
rect 31021 6743 31079 6749
rect 31113 6783 31171 6789
rect 31113 6749 31125 6783
rect 31159 6780 31171 6783
rect 31220 6780 31248 6808
rect 31159 6752 31248 6780
rect 31159 6749 31171 6752
rect 31113 6743 31171 6749
rect 31938 6740 31944 6792
rect 31996 6780 32002 6792
rect 32600 6780 32628 6820
rect 32769 6817 32781 6820
rect 32815 6817 32827 6851
rect 32769 6811 32827 6817
rect 32861 6851 32919 6857
rect 32861 6817 32873 6851
rect 32907 6848 32919 6851
rect 33244 6848 33272 6888
rect 32907 6820 33180 6848
rect 33244 6820 33364 6848
rect 32907 6817 32919 6820
rect 32861 6811 32919 6817
rect 33152 6789 33180 6820
rect 31996 6752 32628 6780
rect 32677 6783 32735 6789
rect 31996 6740 32002 6752
rect 32677 6749 32689 6783
rect 32723 6749 32735 6783
rect 32677 6743 32735 6749
rect 32953 6783 33011 6789
rect 32953 6749 32965 6783
rect 32999 6774 33011 6783
rect 33137 6783 33195 6789
rect 32999 6749 33088 6774
rect 32953 6746 33088 6749
rect 32953 6743 33011 6746
rect 30668 6712 30696 6740
rect 30668 6684 31156 6712
rect 31128 6656 31156 6684
rect 32582 6672 32588 6724
rect 32640 6712 32646 6724
rect 32692 6712 32720 6743
rect 32640 6684 32720 6712
rect 32640 6672 32646 6684
rect 28684 6616 29040 6644
rect 28684 6604 28690 6616
rect 31110 6604 31116 6656
rect 31168 6604 31174 6656
rect 31202 6604 31208 6656
rect 31260 6644 31266 6656
rect 33060 6644 33088 6746
rect 33137 6749 33149 6783
rect 33183 6780 33195 6783
rect 33226 6780 33232 6792
rect 33183 6752 33232 6780
rect 33183 6749 33195 6752
rect 33137 6743 33195 6749
rect 33226 6740 33232 6752
rect 33284 6740 33290 6792
rect 33336 6789 33364 6820
rect 33321 6783 33379 6789
rect 33321 6749 33333 6783
rect 33367 6749 33379 6783
rect 33321 6743 33379 6749
rect 33413 6783 33471 6789
rect 33413 6749 33425 6783
rect 33459 6749 33471 6783
rect 33413 6743 33471 6749
rect 33428 6712 33456 6743
rect 33152 6684 33456 6712
rect 33152 6656 33180 6684
rect 31260 6616 33088 6644
rect 31260 6604 31266 6616
rect 33134 6604 33140 6656
rect 33192 6604 33198 6656
rect 1104 6554 38272 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38272 6554
rect 1104 6480 38272 6502
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6512 6412 6837 6440
rect 6512 6400 6518 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 8018 6400 8024 6452
rect 8076 6400 8082 6452
rect 8202 6400 8208 6452
rect 8260 6400 8266 6452
rect 8294 6400 8300 6452
rect 8352 6400 8358 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 9030 6440 9036 6452
rect 8444 6412 9036 6440
rect 8444 6400 8450 6412
rect 9030 6400 9036 6412
rect 9088 6440 9094 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 9088 6412 9229 6440
rect 9088 6400 9094 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9217 6403 9275 6409
rect 13170 6400 13176 6452
rect 13228 6400 13234 6452
rect 18046 6400 18052 6452
rect 18104 6400 18110 6452
rect 18414 6400 18420 6452
rect 18472 6400 18478 6452
rect 18506 6400 18512 6452
rect 18564 6440 18570 6452
rect 18877 6443 18935 6449
rect 18564 6412 18736 6440
rect 18564 6400 18570 6412
rect 8036 6372 8064 6400
rect 8220 6372 8248 6400
rect 7024 6344 8064 6372
rect 8128 6344 8248 6372
rect 7024 6313 7052 6344
rect 8128 6313 8156 6344
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 7944 6168 7972 6267
rect 8202 6264 8208 6316
rect 8260 6264 8266 6316
rect 8312 6304 8340 6400
rect 11885 6375 11943 6381
rect 9330 6344 9720 6372
rect 9330 6316 9358 6344
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8312 6276 8585 6304
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9692 6313 9720 6344
rect 11885 6341 11897 6375
rect 11931 6372 11943 6375
rect 12066 6372 12072 6384
rect 11931 6344 12072 6372
rect 11931 6341 11943 6344
rect 11885 6335 11943 6341
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 12158 6332 12164 6384
rect 12216 6372 12222 6384
rect 12253 6375 12311 6381
rect 12253 6372 12265 6375
rect 12216 6344 12265 6372
rect 12216 6332 12222 6344
rect 12253 6341 12265 6344
rect 12299 6341 12311 6375
rect 12253 6335 12311 6341
rect 12621 6375 12679 6381
rect 12621 6341 12633 6375
rect 12667 6372 12679 6375
rect 12802 6372 12808 6384
rect 12667 6344 12808 6372
rect 12667 6341 12679 6344
rect 12621 6335 12679 6341
rect 12802 6332 12808 6344
rect 12860 6332 12866 6384
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9421 6276 9505 6304
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 8386 6236 8392 6248
rect 8067 6208 8392 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 9214 6236 9220 6248
rect 8527 6208 9220 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 8110 6168 8116 6180
rect 7944 6140 8116 6168
rect 8110 6128 8116 6140
rect 8168 6128 8174 6180
rect 8294 6128 8300 6180
rect 8352 6128 8358 6180
rect 8570 6128 8576 6180
rect 8628 6128 8634 6180
rect 9232 6168 9260 6196
rect 9421 6168 9449 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 11606 6264 11612 6316
rect 11664 6264 11670 6316
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6304 13507 6307
rect 13722 6304 13728 6316
rect 13495 6276 13728 6304
rect 13495 6273 13507 6276
rect 13449 6267 13507 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 18064 6304 18092 6400
rect 18432 6313 18460 6400
rect 18708 6313 18736 6412
rect 18877 6409 18889 6443
rect 18923 6440 18935 6443
rect 19334 6440 19340 6452
rect 18923 6412 19340 6440
rect 18923 6409 18935 6412
rect 18877 6403 18935 6409
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19426 6400 19432 6452
rect 19484 6400 19490 6452
rect 22370 6400 22376 6452
rect 22428 6400 22434 6452
rect 22922 6440 22928 6452
rect 22480 6412 22928 6440
rect 19061 6375 19119 6381
rect 19061 6341 19073 6375
rect 19107 6372 19119 6375
rect 19444 6372 19472 6400
rect 19107 6344 19472 6372
rect 19107 6341 19119 6344
rect 19061 6335 19119 6341
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 18064 6276 18245 6304
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18417 6307 18475 6313
rect 18417 6273 18429 6307
rect 18463 6273 18475 6307
rect 18417 6267 18475 6273
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 19150 6304 19156 6316
rect 18739 6276 19156 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6236 13139 6239
rect 13127 6208 13584 6236
rect 13127 6205 13139 6208
rect 13081 6199 13139 6205
rect 9232 6140 9449 6168
rect 8386 6060 8392 6112
rect 8444 6060 8450 6112
rect 8588 6100 8616 6128
rect 13556 6112 13584 6208
rect 13630 6196 13636 6248
rect 13688 6196 13694 6248
rect 18248 6236 18276 6267
rect 18524 6236 18552 6267
rect 19150 6264 19156 6276
rect 19208 6304 19214 6316
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 19208 6276 19257 6304
rect 19208 6264 19214 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 18248 6208 18552 6236
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 19352 6236 19380 6344
rect 21910 6264 21916 6316
rect 21968 6304 21974 6316
rect 22388 6313 22416 6400
rect 22480 6313 22508 6412
rect 22922 6400 22928 6412
rect 22980 6400 22986 6452
rect 23109 6443 23167 6449
rect 23109 6409 23121 6443
rect 23155 6440 23167 6443
rect 23198 6440 23204 6452
rect 23155 6412 23204 6440
rect 23155 6409 23167 6412
rect 23109 6403 23167 6409
rect 23198 6400 23204 6412
rect 23256 6400 23262 6452
rect 24118 6400 24124 6452
rect 24176 6440 24182 6452
rect 24679 6443 24737 6449
rect 24176 6412 24624 6440
rect 24176 6400 24182 6412
rect 24596 6372 24624 6412
rect 24679 6409 24691 6443
rect 24725 6440 24737 6443
rect 25130 6440 25136 6452
rect 24725 6412 25136 6440
rect 24725 6409 24737 6412
rect 24679 6403 24737 6409
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 28169 6443 28227 6449
rect 26620 6412 28120 6440
rect 24765 6375 24823 6381
rect 24765 6372 24777 6375
rect 22664 6344 24532 6372
rect 24596 6344 24777 6372
rect 22664 6313 22692 6344
rect 22189 6307 22247 6313
rect 22189 6304 22201 6307
rect 21968 6276 22201 6304
rect 21968 6264 21974 6276
rect 22189 6273 22201 6276
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6273 22431 6307
rect 22373 6267 22431 6273
rect 22465 6307 22523 6313
rect 22465 6273 22477 6307
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 22613 6307 22692 6313
rect 22613 6273 22625 6307
rect 22659 6276 22692 6307
rect 22659 6273 22671 6276
rect 22613 6267 22671 6273
rect 22738 6264 22744 6316
rect 22796 6264 22802 6316
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 22971 6307 23029 6313
rect 22971 6273 22983 6307
rect 23017 6304 23029 6307
rect 23106 6304 23112 6316
rect 23017 6276 23112 6304
rect 23017 6273 23029 6276
rect 22971 6267 23029 6273
rect 18656 6208 19380 6236
rect 22848 6236 22876 6267
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 24394 6264 24400 6316
rect 24452 6264 24458 6316
rect 23842 6236 23848 6248
rect 22848 6208 23848 6236
rect 18656 6196 18662 6208
rect 15194 6128 15200 6180
rect 15252 6168 15258 6180
rect 15746 6168 15752 6180
rect 15252 6140 15752 6168
rect 15252 6128 15258 6140
rect 15746 6128 15752 6140
rect 15804 6128 15810 6180
rect 9309 6103 9367 6109
rect 9309 6100 9321 6103
rect 8588 6072 9321 6100
rect 9309 6069 9321 6072
rect 9355 6069 9367 6103
rect 9309 6063 9367 6069
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9456 6072 9781 6100
rect 9456 6060 9462 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 9769 6063 9827 6069
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 15102 6100 15108 6112
rect 14056 6072 15108 6100
rect 14056 6060 14062 6072
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 18322 6060 18328 6112
rect 18380 6060 18386 6112
rect 18708 6109 18736 6208
rect 23842 6196 23848 6208
rect 23900 6236 23906 6248
rect 24412 6236 24440 6264
rect 23900 6208 24440 6236
rect 24504 6236 24532 6344
rect 24765 6341 24777 6344
rect 24811 6341 24823 6375
rect 24765 6335 24823 6341
rect 25590 6332 25596 6384
rect 25648 6372 25654 6384
rect 26510 6372 26516 6384
rect 25648 6344 26516 6372
rect 25648 6332 25654 6344
rect 26510 6332 26516 6344
rect 26568 6332 26574 6384
rect 24578 6264 24584 6316
rect 24636 6264 24642 6316
rect 24857 6307 24915 6313
rect 24857 6273 24869 6307
rect 24903 6304 24915 6307
rect 24946 6304 24952 6316
rect 24903 6276 24952 6304
rect 24903 6273 24915 6276
rect 24857 6267 24915 6273
rect 24946 6264 24952 6276
rect 25004 6264 25010 6316
rect 26620 6236 26648 6412
rect 26786 6332 26792 6384
rect 26844 6372 26850 6384
rect 28092 6372 28120 6412
rect 28169 6409 28181 6443
rect 28215 6440 28227 6443
rect 28442 6440 28448 6452
rect 28215 6412 28448 6440
rect 28215 6409 28227 6412
rect 28169 6403 28227 6409
rect 28442 6400 28448 6412
rect 28500 6400 28506 6452
rect 31202 6440 31208 6452
rect 30024 6412 31208 6440
rect 28902 6372 28908 6384
rect 26844 6344 28028 6372
rect 28092 6344 28396 6372
rect 26844 6332 26850 6344
rect 28000 6313 28028 6344
rect 27801 6307 27859 6313
rect 27801 6273 27813 6307
rect 27847 6304 27859 6307
rect 27985 6307 28043 6313
rect 27847 6276 27936 6304
rect 27847 6273 27859 6276
rect 27801 6267 27859 6273
rect 27908 6248 27936 6276
rect 27985 6273 27997 6307
rect 28031 6273 28043 6307
rect 27985 6267 28043 6273
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 24504 6208 26648 6236
rect 23900 6196 23906 6208
rect 27890 6196 27896 6248
rect 27948 6196 27954 6248
rect 28092 6236 28120 6267
rect 28000 6208 28120 6236
rect 28368 6236 28396 6344
rect 28460 6344 28908 6372
rect 28460 6316 28488 6344
rect 28902 6332 28908 6344
rect 28960 6372 28966 6384
rect 30024 6372 30052 6412
rect 31202 6400 31208 6412
rect 31260 6400 31266 6452
rect 31938 6400 31944 6452
rect 31996 6400 32002 6452
rect 32122 6400 32128 6452
rect 32180 6400 32186 6452
rect 31573 6375 31631 6381
rect 31573 6372 31585 6375
rect 28960 6344 30052 6372
rect 30116 6344 31585 6372
rect 28960 6332 28966 6344
rect 30116 6316 30144 6344
rect 31573 6341 31585 6344
rect 31619 6341 31631 6375
rect 31573 6335 31631 6341
rect 31754 6332 31760 6384
rect 31812 6372 31818 6384
rect 32030 6372 32036 6384
rect 31812 6344 32036 6372
rect 31812 6332 31818 6344
rect 32030 6332 32036 6344
rect 32088 6332 32094 6384
rect 33134 6372 33140 6384
rect 32600 6344 33140 6372
rect 28442 6264 28448 6316
rect 28500 6264 28506 6316
rect 30098 6264 30104 6316
rect 30156 6264 30162 6316
rect 30285 6307 30343 6313
rect 30285 6273 30297 6307
rect 30331 6304 30343 6307
rect 30374 6304 30380 6316
rect 30331 6276 30380 6304
rect 30331 6273 30343 6276
rect 30285 6267 30343 6273
rect 30374 6264 30380 6276
rect 30432 6264 30438 6316
rect 32048 6304 32076 6332
rect 32600 6316 32628 6344
rect 33134 6332 33140 6344
rect 33192 6332 33198 6384
rect 32401 6307 32459 6313
rect 32401 6304 32413 6307
rect 32048 6276 32413 6304
rect 32401 6273 32413 6276
rect 32447 6273 32459 6307
rect 32401 6267 32459 6273
rect 32490 6264 32496 6316
rect 32548 6264 32554 6316
rect 32582 6264 32588 6316
rect 32640 6264 32646 6316
rect 32769 6307 32827 6313
rect 32769 6273 32781 6307
rect 32815 6273 32827 6307
rect 32769 6267 32827 6273
rect 29638 6236 29644 6248
rect 28368 6208 29644 6236
rect 27614 6168 27620 6180
rect 22848 6140 27620 6168
rect 22848 6112 22876 6140
rect 27614 6128 27620 6140
rect 27672 6128 27678 6180
rect 27801 6171 27859 6177
rect 27801 6137 27813 6171
rect 27847 6168 27859 6171
rect 28000 6168 28028 6208
rect 29638 6196 29644 6208
rect 29696 6236 29702 6248
rect 29696 6208 31754 6236
rect 29696 6196 29702 6208
rect 27847 6140 28028 6168
rect 27847 6137 27859 6140
rect 27801 6131 27859 6137
rect 28718 6128 28724 6180
rect 28776 6168 28782 6180
rect 30285 6171 30343 6177
rect 30285 6168 30297 6171
rect 28776 6140 30297 6168
rect 28776 6128 28782 6140
rect 30285 6137 30297 6140
rect 30331 6137 30343 6171
rect 31726 6168 31754 6208
rect 32030 6196 32036 6248
rect 32088 6236 32094 6248
rect 32600 6236 32628 6264
rect 32088 6208 32628 6236
rect 32088 6196 32094 6208
rect 32784 6168 32812 6267
rect 31726 6140 32812 6168
rect 30285 6131 30343 6137
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6069 18751 6103
rect 18693 6063 18751 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19429 6103 19487 6109
rect 19429 6100 19441 6103
rect 19392 6072 19441 6100
rect 19392 6060 19398 6072
rect 19429 6069 19441 6072
rect 19475 6069 19487 6103
rect 19429 6063 19487 6069
rect 22281 6103 22339 6109
rect 22281 6069 22293 6103
rect 22327 6100 22339 6103
rect 22554 6100 22560 6112
rect 22327 6072 22560 6100
rect 22327 6069 22339 6072
rect 22281 6063 22339 6069
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 22830 6060 22836 6112
rect 22888 6060 22894 6112
rect 26510 6060 26516 6112
rect 26568 6100 26574 6112
rect 33318 6100 33324 6112
rect 26568 6072 33324 6100
rect 26568 6060 26574 6072
rect 33318 6060 33324 6072
rect 33376 6060 33382 6112
rect 1104 6010 38272 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38272 6010
rect 1104 5936 38272 5958
rect 7926 5896 7932 5908
rect 7484 5868 7932 5896
rect 7484 5701 7512 5868
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 9398 5896 9404 5908
rect 9049 5868 9404 5896
rect 7653 5831 7711 5837
rect 7653 5797 7665 5831
rect 7699 5828 7711 5831
rect 8588 5828 8616 5856
rect 7699 5800 8616 5828
rect 7699 5797 7711 5800
rect 7653 5791 7711 5797
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8665 5763 8723 5769
rect 8665 5760 8677 5763
rect 7791 5732 8677 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 8665 5729 8677 5732
rect 8711 5729 8723 5763
rect 9049 5760 9077 5868
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 9508 5868 9720 5896
rect 9214 5788 9220 5840
rect 9272 5788 9278 5840
rect 8665 5723 8723 5729
rect 8956 5732 9077 5760
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5692 8171 5695
rect 8202 5692 8208 5704
rect 8159 5664 8208 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 8956 5701 8984 5732
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9232 5692 9260 5788
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 9088 5664 9133 5692
rect 9232 5664 9321 5692
rect 9088 5652 9094 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9398 5652 9404 5704
rect 9456 5701 9462 5704
rect 9456 5692 9464 5701
rect 9508 5692 9536 5868
rect 9585 5831 9643 5837
rect 9585 5797 9597 5831
rect 9631 5797 9643 5831
rect 9692 5828 9720 5868
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 11664 5868 12633 5896
rect 11664 5856 11670 5868
rect 12621 5865 12633 5868
rect 12667 5865 12679 5899
rect 12621 5859 12679 5865
rect 13078 5856 13084 5908
rect 13136 5856 13142 5908
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 15562 5896 15568 5908
rect 13228 5868 13492 5896
rect 13228 5856 13234 5868
rect 12710 5828 12716 5840
rect 9692 5800 12716 5828
rect 9585 5791 9643 5797
rect 9600 5760 9628 5791
rect 12710 5788 12716 5800
rect 12768 5828 12774 5840
rect 13357 5831 13415 5837
rect 13357 5828 13369 5831
rect 12768 5800 13369 5828
rect 12768 5788 12774 5800
rect 13357 5797 13369 5800
rect 13403 5797 13415 5831
rect 13357 5791 13415 5797
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9600 5732 9689 5760
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 13464 5760 13492 5868
rect 14660 5868 15568 5896
rect 9677 5723 9735 5729
rect 13004 5732 13492 5760
rect 9456 5664 9536 5692
rect 9456 5655 9464 5664
rect 9456 5652 9462 5655
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 9824 5664 10425 5692
rect 9824 5652 9830 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 12158 5652 12164 5704
rect 12216 5692 12222 5704
rect 13004 5701 13032 5732
rect 13538 5720 13544 5772
rect 13596 5760 13602 5772
rect 13596 5732 14412 5760
rect 13596 5720 13602 5732
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 12216 5664 12265 5692
rect 12216 5652 12222 5664
rect 12253 5661 12265 5664
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5661 13047 5695
rect 12989 5655 13047 5661
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 13998 5692 14004 5704
rect 13771 5664 14004 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 8404 5624 8432 5652
rect 9217 5627 9275 5633
rect 9217 5624 9229 5627
rect 8404 5596 9229 5624
rect 9217 5593 9229 5596
rect 9263 5593 9275 5627
rect 12452 5624 12480 5655
rect 9217 5587 9275 5593
rect 12268 5596 12480 5624
rect 13188 5624 13216 5655
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 13188 5596 13921 5624
rect 12268 5568 12296 5596
rect 7282 5516 7288 5568
rect 7340 5516 7346 5568
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10321 5559 10379 5565
rect 10321 5556 10333 5559
rect 10100 5528 10333 5556
rect 10100 5516 10106 5528
rect 10321 5525 10333 5528
rect 10367 5525 10379 5559
rect 10321 5519 10379 5525
rect 11698 5516 11704 5568
rect 11756 5516 11762 5568
rect 12250 5516 12256 5568
rect 12308 5516 12314 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 13188 5556 13216 5596
rect 13909 5593 13921 5596
rect 13955 5593 13967 5627
rect 13909 5587 13967 5593
rect 12860 5528 13216 5556
rect 14384 5556 14412 5732
rect 14660 5701 14688 5868
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 19978 5856 19984 5908
rect 20036 5856 20042 5908
rect 20625 5899 20683 5905
rect 20625 5865 20637 5899
rect 20671 5896 20683 5899
rect 22738 5896 22744 5908
rect 20671 5868 22744 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 22738 5856 22744 5868
rect 22796 5856 22802 5908
rect 24213 5899 24271 5905
rect 24213 5865 24225 5899
rect 24259 5896 24271 5899
rect 24578 5896 24584 5908
rect 24259 5868 24584 5896
rect 24259 5865 24271 5868
rect 24213 5859 24271 5865
rect 24578 5856 24584 5868
rect 24636 5856 24642 5908
rect 27709 5899 27767 5905
rect 27709 5865 27721 5899
rect 27755 5896 27767 5899
rect 28166 5896 28172 5908
rect 27755 5868 28172 5896
rect 27755 5865 27767 5868
rect 27709 5859 27767 5865
rect 28166 5856 28172 5868
rect 28224 5856 28230 5908
rect 28350 5856 28356 5908
rect 28408 5896 28414 5908
rect 29362 5896 29368 5908
rect 28408 5868 29368 5896
rect 28408 5856 28414 5868
rect 29362 5856 29368 5868
rect 29420 5856 29426 5908
rect 29472 5868 30052 5896
rect 15197 5831 15255 5837
rect 15197 5797 15209 5831
rect 15243 5828 15255 5831
rect 19996 5828 20024 5856
rect 29472 5840 29500 5868
rect 30024 5840 30052 5868
rect 30098 5856 30104 5908
rect 30156 5856 30162 5908
rect 31110 5856 31116 5908
rect 31168 5856 31174 5908
rect 32030 5856 32036 5908
rect 32088 5856 32094 5908
rect 32490 5856 32496 5908
rect 32548 5856 32554 5908
rect 15243 5800 15792 5828
rect 15243 5797 15255 5800
rect 15197 5791 15255 5797
rect 15102 5720 15108 5772
rect 15160 5760 15166 5772
rect 15764 5769 15792 5800
rect 19812 5800 20024 5828
rect 22940 5800 25636 5828
rect 15749 5763 15807 5769
rect 15160 5732 15332 5760
rect 15160 5720 15166 5732
rect 15304 5701 15332 5732
rect 15749 5729 15761 5763
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 19812 5701 19840 5800
rect 22940 5772 22968 5800
rect 19889 5763 19947 5769
rect 19889 5729 19901 5763
rect 19935 5760 19947 5763
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 19935 5732 20177 5760
rect 19935 5729 19947 5732
rect 19889 5723 19947 5729
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 22649 5763 22707 5769
rect 22649 5729 22661 5763
rect 22695 5760 22707 5763
rect 22922 5760 22928 5772
rect 22695 5732 22928 5760
rect 22695 5729 22707 5732
rect 22649 5723 22707 5729
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 23382 5760 23388 5772
rect 23216 5732 23388 5760
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 14829 5627 14887 5633
rect 14829 5624 14841 5627
rect 14516 5596 14841 5624
rect 14516 5584 14522 5596
rect 14829 5593 14841 5596
rect 14875 5593 14887 5627
rect 14829 5587 14887 5593
rect 14921 5627 14979 5633
rect 14921 5593 14933 5627
rect 14967 5593 14979 5627
rect 15028 5624 15056 5655
rect 15381 5627 15439 5633
rect 15381 5624 15393 5627
rect 15028 5596 15393 5624
rect 14921 5587 14979 5593
rect 15381 5593 15393 5596
rect 15427 5593 15439 5627
rect 15381 5587 15439 5593
rect 14936 5556 14964 5587
rect 15470 5584 15476 5636
rect 15528 5584 15534 5636
rect 19996 5624 20024 5655
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20257 5695 20315 5701
rect 20257 5692 20269 5695
rect 20128 5664 20269 5692
rect 20128 5652 20134 5664
rect 20257 5661 20269 5664
rect 20303 5661 20315 5695
rect 20257 5655 20315 5661
rect 22554 5652 22560 5704
rect 22612 5652 22618 5704
rect 23216 5701 23244 5732
rect 23382 5720 23388 5732
rect 23440 5760 23446 5772
rect 25608 5760 25636 5800
rect 27982 5788 27988 5840
rect 28040 5828 28046 5840
rect 28040 5800 28396 5828
rect 28040 5788 28046 5800
rect 28368 5760 28396 5800
rect 29454 5788 29460 5840
rect 29512 5788 29518 5840
rect 29914 5788 29920 5840
rect 29972 5788 29978 5840
rect 30006 5788 30012 5840
rect 30064 5828 30070 5840
rect 30469 5831 30527 5837
rect 30469 5828 30481 5831
rect 30064 5800 30481 5828
rect 30064 5788 30070 5800
rect 30469 5797 30481 5800
rect 30515 5797 30527 5831
rect 30469 5791 30527 5797
rect 23440 5732 23704 5760
rect 23440 5720 23446 5732
rect 23676 5701 23704 5732
rect 24136 5732 25360 5760
rect 25608 5732 28028 5760
rect 24136 5704 24164 5732
rect 22741 5695 22799 5701
rect 22741 5661 22753 5695
rect 22787 5692 22799 5695
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 22787 5664 23213 5692
rect 22787 5661 22799 5664
rect 22741 5655 22799 5661
rect 23201 5661 23213 5664
rect 23247 5661 23259 5695
rect 23201 5655 23259 5661
rect 23293 5695 23351 5701
rect 23293 5661 23305 5695
rect 23339 5661 23351 5695
rect 23293 5655 23351 5661
rect 23661 5695 23719 5701
rect 23661 5661 23673 5695
rect 23707 5661 23719 5695
rect 23661 5655 23719 5661
rect 20162 5624 20168 5636
rect 19996 5596 20168 5624
rect 20162 5584 20168 5596
rect 20220 5624 20226 5636
rect 20806 5624 20812 5636
rect 20220 5596 20812 5624
rect 20220 5584 20226 5596
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 22572 5624 22600 5652
rect 23308 5624 23336 5655
rect 23842 5652 23848 5704
rect 23900 5652 23906 5704
rect 23934 5652 23940 5704
rect 23992 5652 23998 5704
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5661 24087 5695
rect 24029 5655 24087 5661
rect 22572 5596 23336 5624
rect 24044 5624 24072 5655
rect 24118 5652 24124 5704
rect 24176 5652 24182 5704
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 24872 5624 24900 5655
rect 24946 5652 24952 5704
rect 25004 5692 25010 5704
rect 25332 5701 25360 5732
rect 25133 5695 25191 5701
rect 25133 5692 25145 5695
rect 25004 5664 25145 5692
rect 25004 5652 25010 5664
rect 25133 5661 25145 5664
rect 25179 5661 25191 5695
rect 25133 5655 25191 5661
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5661 25375 5695
rect 25317 5655 25375 5661
rect 25682 5652 25688 5704
rect 25740 5652 25746 5704
rect 27614 5652 27620 5704
rect 27672 5692 27678 5704
rect 27893 5695 27951 5701
rect 27893 5692 27905 5695
rect 27672 5664 27905 5692
rect 27672 5652 27678 5664
rect 27893 5661 27905 5664
rect 27939 5661 27951 5695
rect 27893 5655 27951 5661
rect 25700 5624 25728 5652
rect 24044 5596 24808 5624
rect 24872 5596 25728 5624
rect 28000 5624 28028 5732
rect 28092 5732 28304 5760
rect 28368 5732 32168 5760
rect 28092 5704 28120 5732
rect 28074 5652 28080 5704
rect 28132 5652 28138 5704
rect 28276 5701 28304 5732
rect 28169 5695 28227 5701
rect 28169 5661 28181 5695
rect 28215 5661 28227 5695
rect 28169 5655 28227 5661
rect 28261 5695 28319 5701
rect 28261 5661 28273 5695
rect 28307 5661 28319 5695
rect 28261 5655 28319 5661
rect 28445 5695 28503 5701
rect 28445 5661 28457 5695
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 28184 5624 28212 5655
rect 28460 5624 28488 5655
rect 29454 5652 29460 5704
rect 29512 5692 29518 5704
rect 29641 5695 29699 5701
rect 29641 5692 29653 5695
rect 29512 5664 29653 5692
rect 29512 5652 29518 5664
rect 29641 5661 29653 5664
rect 29687 5661 29699 5695
rect 29641 5655 29699 5661
rect 29914 5652 29920 5704
rect 29972 5692 29978 5704
rect 30193 5695 30251 5701
rect 30193 5692 30205 5695
rect 29972 5664 30205 5692
rect 29972 5652 29978 5664
rect 30193 5661 30205 5664
rect 30239 5661 30251 5695
rect 30193 5655 30251 5661
rect 30834 5652 30840 5704
rect 30892 5692 30898 5704
rect 30929 5695 30987 5701
rect 30929 5692 30941 5695
rect 30892 5664 30941 5692
rect 30892 5652 30898 5664
rect 30929 5661 30941 5664
rect 30975 5661 30987 5695
rect 30929 5655 30987 5661
rect 31938 5652 31944 5704
rect 31996 5652 32002 5704
rect 32140 5701 32168 5732
rect 32125 5695 32183 5701
rect 32125 5661 32137 5695
rect 32171 5692 32183 5695
rect 32508 5692 32536 5856
rect 32171 5664 32536 5692
rect 32171 5661 32183 5664
rect 32125 5655 32183 5661
rect 28000 5596 28488 5624
rect 15488 5556 15516 5584
rect 14384 5528 15516 5556
rect 12860 5516 12866 5528
rect 16390 5516 16396 5568
rect 16448 5516 16454 5568
rect 22830 5516 22836 5568
rect 22888 5516 22894 5568
rect 23474 5516 23480 5568
rect 23532 5516 23538 5568
rect 24670 5516 24676 5568
rect 24728 5516 24734 5568
rect 24780 5556 24808 5596
rect 30742 5584 30748 5636
rect 30800 5584 30806 5636
rect 27430 5556 27436 5568
rect 24780 5528 27436 5556
rect 27430 5516 27436 5528
rect 27488 5516 27494 5568
rect 29730 5516 29736 5568
rect 29788 5556 29794 5568
rect 30374 5556 30380 5568
rect 29788 5528 30380 5556
rect 29788 5516 29794 5528
rect 30374 5516 30380 5528
rect 30432 5556 30438 5568
rect 30653 5559 30711 5565
rect 30653 5556 30665 5559
rect 30432 5528 30665 5556
rect 30432 5516 30438 5528
rect 30653 5525 30665 5528
rect 30699 5525 30711 5559
rect 30653 5519 30711 5525
rect 1104 5466 38272 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38272 5466
rect 1104 5392 38272 5414
rect 7282 5352 7288 5364
rect 6656 5324 7288 5352
rect 6656 5293 6684 5324
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 8113 5355 8171 5361
rect 7524 5324 7788 5352
rect 7524 5312 7530 5324
rect 6641 5287 6699 5293
rect 6641 5253 6653 5287
rect 6687 5253 6699 5287
rect 6641 5247 6699 5253
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6144 5188 6377 5216
rect 6144 5176 6150 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 7760 5202 7788 5324
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 8202 5352 8208 5364
rect 8159 5324 8208 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 9401 5355 9459 5361
rect 9401 5352 9413 5355
rect 9088 5324 9413 5352
rect 9088 5312 9094 5324
rect 9401 5321 9413 5324
rect 9447 5321 9459 5355
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 9401 5315 9459 5321
rect 9646 5324 12173 5352
rect 9125 5287 9183 5293
rect 8680 5256 9076 5284
rect 8680 5228 8708 5256
rect 8389 5219 8447 5225
rect 6365 5179 6423 5185
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 8478 5216 8484 5228
rect 8435 5188 8484 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 8662 5176 8668 5228
rect 8720 5176 8726 5228
rect 9048 5225 9076 5256
rect 9125 5253 9137 5287
rect 9171 5284 9183 5287
rect 9646 5284 9674 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12526 5352 12532 5364
rect 12483 5324 12532 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 9171 5256 9674 5284
rect 9769 5287 9827 5293
rect 9171 5253 9183 5256
rect 9125 5247 9183 5253
rect 9769 5253 9781 5287
rect 9815 5284 9827 5287
rect 10042 5284 10048 5296
rect 9815 5256 10048 5284
rect 9815 5253 9827 5256
rect 9769 5247 9827 5253
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 12452 5284 12480 5315
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 13630 5352 13636 5364
rect 12728 5324 13636 5352
rect 11072 5256 12480 5284
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8905 5219 8963 5225
rect 8905 5185 8917 5219
rect 8951 5185 8963 5219
rect 8905 5179 8963 5185
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 9263 5219 9321 5225
rect 9263 5185 9275 5219
rect 9309 5216 9321 5219
rect 9398 5216 9404 5228
rect 9309 5188 9404 5216
rect 9309 5185 9321 5188
rect 9263 5179 9321 5185
rect 8496 5148 8524 5176
rect 8772 5148 8800 5179
rect 8496 5120 8800 5148
rect 8920 5148 8948 5179
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9490 5176 9496 5228
rect 9548 5176 9554 5228
rect 10870 5176 10876 5228
rect 10928 5176 10934 5228
rect 11072 5216 11100 5256
rect 12250 5216 12256 5228
rect 10980 5188 11100 5216
rect 11256 5188 12256 5216
rect 10980 5148 11008 5188
rect 8920 5120 11008 5148
rect 9306 5040 9312 5092
rect 9364 5040 9370 5092
rect 8202 4972 8208 5024
rect 8260 4972 8266 5024
rect 9324 5012 9352 5040
rect 11256 5021 11284 5188
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 12728 5225 12756 5324
rect 13630 5312 13636 5324
rect 13688 5352 13694 5364
rect 13725 5355 13783 5361
rect 13725 5352 13737 5355
rect 13688 5324 13737 5352
rect 13688 5312 13694 5324
rect 13725 5321 13737 5324
rect 13771 5321 13783 5355
rect 13725 5315 13783 5321
rect 14458 5312 14464 5364
rect 14516 5312 14522 5364
rect 15286 5352 15292 5364
rect 14660 5324 15292 5352
rect 13078 5244 13084 5296
rect 13136 5284 13142 5296
rect 13136 5256 14044 5284
rect 13136 5244 13142 5256
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 12158 5148 12164 5160
rect 11572 5120 12164 5148
rect 11572 5108 11578 5120
rect 12158 5108 12164 5120
rect 12216 5148 12222 5160
rect 12452 5148 12480 5179
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 13817 5219 13875 5225
rect 13817 5216 13829 5219
rect 13780 5188 13829 5216
rect 13780 5176 13786 5188
rect 13817 5185 13829 5188
rect 13863 5185 13875 5219
rect 13817 5179 13875 5185
rect 14016 5157 14044 5256
rect 14660 5225 14688 5324
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15470 5312 15476 5364
rect 15528 5352 15534 5364
rect 16439 5355 16497 5361
rect 16439 5352 16451 5355
rect 15528 5324 16451 5352
rect 15528 5312 15534 5324
rect 16439 5321 16451 5324
rect 16485 5321 16497 5355
rect 16439 5315 16497 5321
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 28166 5352 28172 5364
rect 19392 5324 20116 5352
rect 19392 5312 19398 5324
rect 16574 5284 16580 5296
rect 16054 5256 16580 5284
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 15102 5216 15108 5228
rect 14645 5179 14703 5185
rect 14752 5188 15108 5216
rect 12216 5120 12480 5148
rect 14001 5151 14059 5157
rect 12216 5108 12222 5120
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14384 5148 14412 5179
rect 14752 5148 14780 5188
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 16390 5176 16396 5228
rect 16448 5176 16454 5228
rect 14047 5120 14780 5148
rect 15013 5151 15071 5157
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 15013 5117 15025 5151
rect 15059 5148 15071 5151
rect 16408 5148 16436 5176
rect 15059 5120 16436 5148
rect 15059 5117 15071 5120
rect 15013 5111 15071 5117
rect 13446 5040 13452 5092
rect 13504 5080 13510 5092
rect 13504 5052 13768 5080
rect 13504 5040 13510 5052
rect 11241 5015 11299 5021
rect 11241 5012 11253 5015
rect 9324 4984 11253 5012
rect 11241 4981 11253 4984
rect 11287 4981 11299 5015
rect 11241 4975 11299 4981
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 13630 5012 13636 5024
rect 13403 4984 13636 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13740 5012 13768 5052
rect 16500 5012 16528 5256
rect 16574 5244 16580 5256
rect 16632 5244 16638 5296
rect 18322 5244 18328 5296
rect 18380 5284 18386 5296
rect 19242 5284 19248 5296
rect 18380 5256 19248 5284
rect 18380 5244 18386 5256
rect 19242 5244 19248 5256
rect 19300 5284 19306 5296
rect 19705 5287 19763 5293
rect 19300 5256 19472 5284
rect 19300 5244 19306 5256
rect 19334 5176 19340 5228
rect 19392 5176 19398 5228
rect 19444 5225 19472 5256
rect 19705 5253 19717 5287
rect 19751 5284 19763 5287
rect 19978 5284 19984 5296
rect 19751 5256 19984 5284
rect 19751 5253 19763 5256
rect 19705 5247 19763 5253
rect 19978 5244 19984 5256
rect 20036 5244 20042 5296
rect 20088 5225 20116 5324
rect 22066 5324 28172 5352
rect 20162 5244 20168 5296
rect 20220 5244 20226 5296
rect 20809 5287 20867 5293
rect 20809 5253 20821 5287
rect 20855 5284 20867 5287
rect 21453 5287 21511 5293
rect 21453 5284 21465 5287
rect 20855 5256 21465 5284
rect 20855 5253 20867 5256
rect 20809 5247 20867 5253
rect 21453 5253 21465 5256
rect 21499 5284 21511 5287
rect 22066 5284 22094 5324
rect 28166 5312 28172 5324
rect 28224 5312 28230 5364
rect 30101 5355 30159 5361
rect 29656 5324 30052 5352
rect 23474 5284 23480 5296
rect 21499 5256 22094 5284
rect 22756 5256 23480 5284
rect 21499 5253 21511 5256
rect 21453 5247 21511 5253
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5216 19487 5219
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19475 5188 19901 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 20073 5219 20131 5225
rect 20073 5185 20085 5219
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 19797 5151 19855 5157
rect 19797 5117 19809 5151
rect 19843 5148 19855 5151
rect 20180 5148 20208 5244
rect 20254 5176 20260 5228
rect 20312 5216 20318 5228
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 20312 5188 20545 5216
rect 20312 5176 20318 5188
rect 20533 5185 20545 5188
rect 20579 5185 20591 5219
rect 20533 5179 20591 5185
rect 21266 5176 21272 5228
rect 21324 5176 21330 5228
rect 22756 5225 22784 5256
rect 23474 5244 23480 5256
rect 23532 5244 23538 5296
rect 23584 5256 23796 5284
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 23198 5176 23204 5228
rect 23256 5176 23262 5228
rect 23382 5176 23388 5228
rect 23440 5216 23446 5228
rect 23584 5216 23612 5256
rect 23768 5225 23796 5256
rect 24302 5244 24308 5296
rect 24360 5244 24366 5296
rect 23440 5188 23612 5216
rect 23753 5219 23811 5225
rect 23440 5176 23446 5188
rect 23753 5185 23765 5219
rect 23799 5185 23811 5219
rect 23753 5179 23811 5185
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23900 5188 23949 5216
rect 23900 5176 23906 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 29546 5176 29552 5228
rect 29604 5216 29610 5228
rect 29656 5225 29684 5324
rect 29641 5219 29699 5225
rect 29641 5216 29653 5219
rect 29604 5188 29653 5216
rect 29604 5176 29610 5188
rect 29641 5185 29653 5188
rect 29687 5185 29699 5219
rect 29641 5179 29699 5185
rect 29730 5176 29736 5228
rect 29788 5176 29794 5228
rect 29917 5219 29975 5225
rect 29917 5185 29929 5219
rect 29963 5185 29975 5219
rect 30024 5222 30052 5324
rect 30101 5321 30113 5355
rect 30147 5352 30159 5355
rect 30834 5352 30840 5364
rect 30147 5324 30840 5352
rect 30147 5321 30159 5324
rect 30101 5315 30159 5321
rect 30834 5312 30840 5324
rect 30892 5312 30898 5364
rect 31573 5355 31631 5361
rect 31573 5321 31585 5355
rect 31619 5352 31631 5355
rect 31938 5352 31944 5364
rect 31619 5324 31944 5352
rect 31619 5321 31631 5324
rect 31573 5315 31631 5321
rect 31938 5312 31944 5324
rect 31996 5312 32002 5364
rect 31754 5244 31760 5296
rect 31812 5244 31818 5296
rect 30024 5216 30144 5222
rect 30285 5219 30343 5225
rect 30285 5216 30297 5219
rect 30024 5194 30297 5216
rect 30116 5188 30297 5194
rect 29917 5179 29975 5185
rect 30285 5185 30297 5188
rect 30331 5185 30343 5219
rect 30285 5179 30343 5185
rect 30561 5219 30619 5225
rect 30561 5185 30573 5219
rect 30607 5185 30619 5219
rect 30561 5179 30619 5185
rect 19843 5120 20208 5148
rect 19843 5117 19855 5120
rect 19797 5111 19855 5117
rect 20346 5108 20352 5160
rect 20404 5108 20410 5160
rect 20901 5151 20959 5157
rect 20901 5117 20913 5151
rect 20947 5117 20959 5151
rect 20901 5111 20959 5117
rect 22833 5151 22891 5157
rect 22833 5117 22845 5151
rect 22879 5148 22891 5151
rect 23017 5151 23075 5157
rect 23017 5148 23029 5151
rect 22879 5120 23029 5148
rect 22879 5117 22891 5120
rect 22833 5111 22891 5117
rect 23017 5117 23029 5120
rect 23063 5117 23075 5151
rect 23017 5111 23075 5117
rect 20070 5040 20076 5092
rect 20128 5080 20134 5092
rect 20916 5080 20944 5111
rect 29822 5108 29828 5160
rect 29880 5108 29886 5160
rect 24946 5080 24952 5092
rect 20128 5052 20944 5080
rect 22066 5052 24952 5080
rect 20128 5040 20134 5052
rect 13740 4984 16528 5012
rect 19150 4972 19156 5024
rect 19208 4972 19214 5024
rect 19610 4972 19616 5024
rect 19668 5012 19674 5024
rect 20622 5012 20628 5024
rect 19668 4984 20628 5012
rect 19668 4972 19674 4984
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 21637 5015 21695 5021
rect 21637 4981 21649 5015
rect 21683 5012 21695 5015
rect 22066 5012 22094 5052
rect 24946 5040 24952 5052
rect 25004 5040 25010 5092
rect 28166 5040 28172 5092
rect 28224 5080 28230 5092
rect 29921 5080 29949 5179
rect 30190 5108 30196 5160
rect 30248 5148 30254 5160
rect 30576 5148 30604 5179
rect 30650 5176 30656 5228
rect 30708 5216 30714 5228
rect 30745 5219 30803 5225
rect 30745 5216 30757 5219
rect 30708 5188 30757 5216
rect 30708 5176 30714 5188
rect 30745 5185 30757 5188
rect 30791 5216 30803 5219
rect 31205 5219 31263 5225
rect 31205 5216 31217 5219
rect 30791 5188 31217 5216
rect 30791 5185 30803 5188
rect 30745 5179 30803 5185
rect 31205 5185 31217 5188
rect 31251 5216 31263 5219
rect 31772 5216 31800 5244
rect 31251 5188 31800 5216
rect 31251 5185 31263 5188
rect 31205 5179 31263 5185
rect 31113 5151 31171 5157
rect 31113 5148 31125 5151
rect 30248 5120 31125 5148
rect 30248 5108 30254 5120
rect 31113 5117 31125 5120
rect 31159 5117 31171 5151
rect 31113 5111 31171 5117
rect 30208 5080 30236 5108
rect 28224 5052 29776 5080
rect 29921 5052 30236 5080
rect 28224 5040 28230 5052
rect 21683 4984 22094 5012
rect 21683 4981 21695 4984
rect 21637 4975 21695 4981
rect 23934 4972 23940 5024
rect 23992 5012 23998 5024
rect 25130 5012 25136 5024
rect 23992 4984 25136 5012
rect 23992 4972 23998 4984
rect 25130 4972 25136 4984
rect 25188 5012 25194 5024
rect 25682 5012 25688 5024
rect 25188 4984 25688 5012
rect 25188 4972 25194 4984
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 29454 4972 29460 5024
rect 29512 4972 29518 5024
rect 29748 5012 29776 5052
rect 30374 5040 30380 5092
rect 30432 5040 30438 5092
rect 30469 5083 30527 5089
rect 30469 5049 30481 5083
rect 30515 5049 30527 5083
rect 30469 5043 30527 5049
rect 29822 5012 29828 5024
rect 29748 4984 29828 5012
rect 29822 4972 29828 4984
rect 29880 5012 29886 5024
rect 30484 5012 30512 5043
rect 29880 4984 30512 5012
rect 29880 4972 29886 4984
rect 1104 4922 38272 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38272 4922
rect 1104 4848 38272 4870
rect 6720 4811 6778 4817
rect 6720 4777 6732 4811
rect 6766 4808 6778 4811
rect 8202 4808 8208 4820
rect 6766 4780 8208 4808
rect 6766 4777 6778 4780
rect 6720 4771 6778 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8662 4768 8668 4820
rect 8720 4808 8726 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 8720 4780 9321 4808
rect 8720 4768 8726 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9750 4811 9808 4817
rect 9750 4808 9762 4811
rect 9309 4771 9367 4777
rect 9508 4780 9762 4808
rect 9030 4700 9036 4752
rect 9088 4740 9094 4752
rect 9508 4740 9536 4780
rect 9750 4777 9762 4780
rect 9796 4777 9808 4811
rect 9750 4771 9808 4777
rect 13538 4768 13544 4820
rect 13596 4808 13602 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13596 4780 13645 4808
rect 13596 4768 13602 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 13872 4780 15424 4808
rect 13872 4768 13878 4780
rect 9088 4712 9536 4740
rect 13725 4743 13783 4749
rect 9088 4700 9094 4712
rect 13725 4709 13737 4743
rect 13771 4740 13783 4743
rect 15396 4740 15424 4780
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 16577 4811 16635 4817
rect 16577 4808 16589 4811
rect 15620 4780 16589 4808
rect 15620 4768 15626 4780
rect 16577 4777 16589 4780
rect 16623 4777 16635 4811
rect 16577 4771 16635 4777
rect 19150 4768 19156 4820
rect 19208 4768 19214 4820
rect 19981 4811 20039 4817
rect 19981 4777 19993 4811
rect 20027 4808 20039 4811
rect 20070 4808 20076 4820
rect 20027 4780 20076 4808
rect 20027 4777 20039 4780
rect 19981 4771 20039 4777
rect 20070 4768 20076 4780
rect 20128 4768 20134 4820
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 20312 4780 20361 4808
rect 20312 4768 20318 4780
rect 20349 4777 20361 4780
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 20533 4811 20591 4817
rect 20533 4777 20545 4811
rect 20579 4808 20591 4811
rect 21266 4808 21272 4820
rect 20579 4780 21272 4808
rect 20579 4777 20591 4780
rect 20533 4771 20591 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 24581 4811 24639 4817
rect 24581 4808 24593 4811
rect 23256 4780 24593 4808
rect 23256 4768 23262 4780
rect 24581 4777 24593 4780
rect 24627 4777 24639 4811
rect 24581 4771 24639 4777
rect 24670 4768 24676 4820
rect 24728 4768 24734 4820
rect 25314 4768 25320 4820
rect 25372 4808 25378 4820
rect 25590 4808 25596 4820
rect 25372 4780 25596 4808
rect 25372 4768 25378 4780
rect 25590 4768 25596 4780
rect 25648 4768 25654 4820
rect 25682 4768 25688 4820
rect 25740 4808 25746 4820
rect 25866 4808 25872 4820
rect 25740 4780 25872 4808
rect 25740 4768 25746 4780
rect 25866 4768 25872 4780
rect 25924 4808 25930 4820
rect 26053 4811 26111 4817
rect 26053 4808 26065 4811
rect 25924 4780 26065 4808
rect 25924 4768 25930 4780
rect 26053 4777 26065 4780
rect 26099 4777 26111 4811
rect 26053 4771 26111 4777
rect 26418 4768 26424 4820
rect 26476 4768 26482 4820
rect 27706 4808 27712 4820
rect 27080 4780 27712 4808
rect 15841 4743 15899 4749
rect 15841 4740 15853 4743
rect 13771 4712 14228 4740
rect 15396 4712 15853 4740
rect 13771 4709 13783 4712
rect 13725 4703 13783 4709
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 6236 4644 6469 4672
rect 6236 4632 6242 4644
rect 6457 4641 6469 4644
rect 6503 4672 6515 4675
rect 9490 4672 9496 4684
rect 6503 4644 9496 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 9490 4632 9496 4644
rect 9548 4672 9554 4684
rect 11698 4672 11704 4684
rect 9548 4644 11704 4672
rect 9548 4632 9554 4644
rect 11698 4632 11704 4644
rect 11756 4672 11762 4684
rect 11885 4675 11943 4681
rect 11885 4672 11897 4675
rect 11756 4644 11897 4672
rect 11756 4632 11762 4644
rect 11885 4641 11897 4644
rect 11931 4672 11943 4675
rect 14200 4672 14228 4712
rect 15841 4709 15853 4712
rect 15887 4740 15899 4743
rect 19168 4740 19196 4768
rect 23937 4743 23995 4749
rect 15887 4712 15976 4740
rect 19168 4712 23888 4740
rect 15887 4709 15899 4712
rect 15841 4703 15899 4709
rect 15948 4681 15976 4712
rect 14369 4675 14427 4681
rect 14369 4672 14381 4675
rect 11931 4644 14136 4672
rect 14200 4644 14381 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 2590 4604 2596 4616
rect 1535 4576 2596 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9306 4604 9312 4616
rect 8987 4576 9312 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 13446 4604 13452 4616
rect 10928 4576 11652 4604
rect 13294 4590 13452 4604
rect 10928 4564 10934 4576
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 934 4428 940 4480
rect 992 4468 998 4480
rect 1581 4471 1639 4477
rect 1581 4468 1593 4471
rect 992 4440 1593 4468
rect 992 4428 998 4440
rect 1581 4437 1593 4440
rect 1627 4437 1639 4471
rect 1581 4431 1639 4437
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 8312 4468 8340 4564
rect 9125 4539 9183 4545
rect 9125 4505 9137 4539
rect 9171 4536 9183 4539
rect 9214 4536 9220 4548
rect 9171 4508 9220 4536
rect 9171 4505 9183 4508
rect 9125 4499 9183 4505
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 8251 4440 8340 4468
rect 9232 4468 9260 4496
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 9232 4440 11253 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 11241 4437 11253 4440
rect 11287 4468 11299 4471
rect 11514 4468 11520 4480
rect 11287 4440 11520 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 11624 4468 11652 4576
rect 13280 4576 13452 4590
rect 12161 4539 12219 4545
rect 12161 4505 12173 4539
rect 12207 4536 12219 4539
rect 12434 4536 12440 4548
rect 12207 4508 12440 4536
rect 12207 4505 12219 4508
rect 12161 4499 12219 4505
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 13280 4468 13308 4576
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 14108 4613 14136 4644
rect 14369 4641 14381 4644
rect 14415 4641 14427 4675
rect 14369 4635 14427 4641
rect 15933 4675 15991 4681
rect 15933 4641 15945 4675
rect 15979 4641 15991 4675
rect 15933 4635 15991 4641
rect 19334 4632 19340 4684
rect 19392 4632 19398 4684
rect 19610 4632 19616 4684
rect 19668 4632 19674 4684
rect 20438 4672 20444 4684
rect 19720 4644 20444 4672
rect 13909 4607 13967 4613
rect 13909 4604 13921 4607
rect 13688 4576 13921 4604
rect 13688 4564 13694 4576
rect 13909 4573 13921 4576
rect 13955 4573 13967 4607
rect 13909 4567 13967 4573
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 11624 4440 13308 4468
rect 14108 4468 14136 4567
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19352 4604 19380 4632
rect 19720 4613 19748 4644
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 21358 4632 21364 4684
rect 21416 4672 21422 4684
rect 23293 4675 23351 4681
rect 21416 4644 22968 4672
rect 21416 4632 21422 4644
rect 22940 4616 22968 4644
rect 23293 4641 23305 4675
rect 23339 4672 23351 4675
rect 23382 4672 23388 4684
rect 23339 4644 23388 4672
rect 23339 4641 23351 4644
rect 23293 4635 23351 4641
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19352 4576 19441 4604
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 22649 4607 22707 4613
rect 19705 4567 19763 4573
rect 20088 4576 22094 4604
rect 15010 4496 15016 4548
rect 15068 4496 15074 4548
rect 20088 4536 20116 4576
rect 19444 4508 20116 4536
rect 20165 4539 20223 4545
rect 15286 4468 15292 4480
rect 14108 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 19444 4477 19472 4508
rect 20165 4505 20177 4539
rect 20211 4505 20223 4539
rect 20165 4499 20223 4505
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4437 19487 4471
rect 19429 4431 19487 4437
rect 20070 4428 20076 4480
rect 20128 4468 20134 4480
rect 20180 4468 20208 4499
rect 20346 4496 20352 4548
rect 20404 4545 20410 4548
rect 20404 4539 20423 4545
rect 20411 4505 20423 4539
rect 20404 4499 20423 4505
rect 20404 4496 20410 4499
rect 20128 4440 20208 4468
rect 22066 4468 22094 4576
rect 22649 4573 22661 4607
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 22664 4536 22692 4567
rect 22922 4564 22928 4616
rect 22980 4564 22986 4616
rect 23860 4604 23888 4712
rect 23937 4709 23949 4743
rect 23983 4709 23995 4743
rect 23937 4703 23995 4709
rect 23952 4672 23980 4703
rect 24688 4681 24716 4768
rect 25222 4700 25228 4752
rect 25280 4740 25286 4752
rect 27080 4740 27108 4780
rect 27706 4768 27712 4780
rect 27764 4808 27770 4820
rect 28442 4808 28448 4820
rect 27764 4780 28448 4808
rect 27764 4768 27770 4780
rect 28442 4768 28448 4780
rect 28500 4768 28506 4820
rect 29454 4768 29460 4820
rect 29512 4768 29518 4820
rect 30006 4768 30012 4820
rect 30064 4768 30070 4820
rect 30190 4768 30196 4820
rect 30248 4808 30254 4820
rect 30285 4811 30343 4817
rect 30285 4808 30297 4811
rect 30248 4780 30297 4808
rect 30248 4768 30254 4780
rect 30285 4777 30297 4780
rect 30331 4777 30343 4811
rect 30285 4771 30343 4777
rect 30377 4811 30435 4817
rect 30377 4777 30389 4811
rect 30423 4808 30435 4811
rect 30742 4808 30748 4820
rect 30423 4780 30748 4808
rect 30423 4777 30435 4780
rect 30377 4771 30435 4777
rect 30742 4768 30748 4780
rect 30800 4768 30806 4820
rect 25280 4712 27108 4740
rect 27157 4743 27215 4749
rect 25280 4700 25286 4712
rect 27157 4709 27169 4743
rect 27203 4740 27215 4743
rect 28074 4740 28080 4752
rect 27203 4712 28080 4740
rect 27203 4709 27215 4712
rect 27157 4703 27215 4709
rect 28074 4700 28080 4712
rect 28132 4700 28138 4752
rect 28718 4700 28724 4752
rect 28776 4700 28782 4752
rect 24673 4675 24731 4681
rect 23952 4644 24440 4672
rect 24412 4613 24440 4644
rect 24673 4641 24685 4675
rect 24719 4641 24731 4675
rect 24673 4635 24731 4641
rect 24765 4675 24823 4681
rect 24765 4641 24777 4675
rect 24811 4641 24823 4675
rect 26881 4675 26939 4681
rect 24765 4635 24823 4641
rect 24964 4644 25912 4672
rect 24213 4607 24271 4613
rect 24213 4604 24225 4607
rect 23860 4576 24225 4604
rect 24213 4573 24225 4576
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 24397 4607 24455 4613
rect 24397 4573 24409 4607
rect 24443 4573 24455 4607
rect 24397 4567 24455 4573
rect 24489 4607 24547 4613
rect 24489 4573 24501 4607
rect 24535 4604 24547 4607
rect 24780 4604 24808 4635
rect 24964 4613 24992 4644
rect 24535 4576 24808 4604
rect 24949 4607 25007 4613
rect 24535 4573 24547 4576
rect 24489 4567 24547 4573
rect 24949 4573 24961 4607
rect 24995 4573 25007 4607
rect 24949 4567 25007 4573
rect 25041 4607 25099 4613
rect 25041 4573 25053 4607
rect 25087 4573 25099 4607
rect 25041 4567 25099 4573
rect 25133 4607 25191 4613
rect 25133 4573 25145 4607
rect 25179 4573 25191 4607
rect 25133 4567 25191 4573
rect 23937 4539 23995 4545
rect 23937 4536 23949 4539
rect 22664 4508 23949 4536
rect 23937 4505 23949 4508
rect 23983 4536 23995 4539
rect 24026 4536 24032 4548
rect 23983 4508 24032 4536
rect 23983 4505 23995 4508
rect 23937 4499 23995 4505
rect 24026 4496 24032 4508
rect 24084 4496 24090 4548
rect 24228 4536 24256 4567
rect 24964 4536 24992 4567
rect 24228 4508 24992 4536
rect 24121 4471 24179 4477
rect 24121 4468 24133 4471
rect 22066 4440 24133 4468
rect 20128 4428 20134 4440
rect 24121 4437 24133 4440
rect 24167 4468 24179 4471
rect 25056 4468 25084 4567
rect 25148 4536 25176 4567
rect 25222 4564 25228 4616
rect 25280 4564 25286 4616
rect 25498 4604 25504 4616
rect 25332 4576 25504 4604
rect 25332 4536 25360 4576
rect 25498 4564 25504 4576
rect 25556 4564 25562 4616
rect 25590 4564 25596 4616
rect 25648 4564 25654 4616
rect 25884 4613 25912 4644
rect 26881 4641 26893 4675
rect 26927 4672 26939 4675
rect 27062 4672 27068 4684
rect 26927 4644 27068 4672
rect 26927 4641 26939 4644
rect 26881 4635 26939 4641
rect 27062 4632 27068 4644
rect 27120 4672 27126 4684
rect 27120 4644 27660 4672
rect 27120 4632 27126 4644
rect 25869 4607 25927 4613
rect 25869 4573 25881 4607
rect 25915 4573 25927 4607
rect 25869 4567 25927 4573
rect 25958 4564 25964 4616
rect 26016 4564 26022 4616
rect 26786 4564 26792 4616
rect 26844 4564 26850 4616
rect 27632 4613 27660 4644
rect 28534 4632 28540 4684
rect 28592 4632 28598 4684
rect 27617 4607 27675 4613
rect 27617 4573 27629 4607
rect 27663 4604 27675 4607
rect 28629 4607 28687 4613
rect 28629 4604 28641 4607
rect 27663 4576 28641 4604
rect 27663 4573 27675 4576
rect 27617 4567 27675 4573
rect 28629 4573 28641 4576
rect 28675 4604 28687 4607
rect 28736 4604 28764 4700
rect 29270 4632 29276 4684
rect 29328 4632 29334 4684
rect 29472 4672 29500 4768
rect 29472 4644 30420 4672
rect 28675 4576 28764 4604
rect 29825 4607 29883 4613
rect 28675 4573 28687 4576
rect 28629 4567 28687 4573
rect 29825 4573 29837 4607
rect 29871 4604 29883 4607
rect 29914 4604 29920 4616
rect 29871 4576 29920 4604
rect 29871 4573 29883 4576
rect 29825 4567 29883 4573
rect 29914 4564 29920 4576
rect 29972 4564 29978 4616
rect 30392 4613 30420 4644
rect 30377 4607 30435 4613
rect 30377 4573 30389 4607
rect 30423 4573 30435 4607
rect 30377 4567 30435 4573
rect 30561 4607 30619 4613
rect 30561 4573 30573 4607
rect 30607 4604 30619 4607
rect 30650 4604 30656 4616
rect 30607 4576 30656 4604
rect 30607 4573 30619 4576
rect 30561 4567 30619 4573
rect 30650 4564 30656 4576
rect 30708 4564 30714 4616
rect 25148 4508 25360 4536
rect 25409 4539 25467 4545
rect 25409 4505 25421 4539
rect 25455 4536 25467 4539
rect 26510 4536 26516 4548
rect 25455 4508 26516 4536
rect 25455 4505 25467 4508
rect 25409 4499 25467 4505
rect 26510 4496 26516 4508
rect 26568 4536 26574 4548
rect 26878 4536 26884 4548
rect 26568 4508 26884 4536
rect 26568 4496 26574 4508
rect 26878 4496 26884 4508
rect 26936 4496 26942 4548
rect 27430 4496 27436 4548
rect 27488 4496 27494 4548
rect 25777 4471 25835 4477
rect 25777 4468 25789 4471
rect 24167 4440 25789 4468
rect 24167 4437 24179 4440
rect 24121 4431 24179 4437
rect 25777 4437 25789 4440
rect 25823 4437 25835 4471
rect 25777 4431 25835 4437
rect 27801 4471 27859 4477
rect 27801 4437 27813 4471
rect 27847 4468 27859 4471
rect 27890 4468 27896 4480
rect 27847 4440 27896 4468
rect 27847 4437 27859 4440
rect 27801 4431 27859 4437
rect 27890 4428 27896 4440
rect 27948 4428 27954 4480
rect 1104 4378 38272 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38272 4378
rect 1104 4304 38272 4326
rect 8570 4224 8576 4276
rect 8628 4264 8634 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8628 4236 9045 4264
rect 8628 4224 8634 4236
rect 9033 4233 9045 4236
rect 9079 4233 9091 4267
rect 9033 4227 9091 4233
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 12621 4267 12679 4273
rect 12621 4264 12633 4267
rect 12492 4236 12633 4264
rect 12492 4224 12498 4236
rect 12621 4233 12633 4236
rect 12667 4233 12679 4267
rect 12621 4227 12679 4233
rect 12989 4267 13047 4273
rect 12989 4233 13001 4267
rect 13035 4264 13047 4267
rect 13262 4264 13268 4276
rect 13035 4236 13268 4264
rect 13035 4233 13047 4236
rect 12989 4227 13047 4233
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 25130 4224 25136 4276
rect 25188 4224 25194 4276
rect 25314 4224 25320 4276
rect 25372 4264 25378 4276
rect 25409 4267 25467 4273
rect 25409 4264 25421 4267
rect 25372 4236 25421 4264
rect 25372 4224 25378 4236
rect 25409 4233 25421 4236
rect 25455 4233 25467 4267
rect 25409 4227 25467 4233
rect 25777 4267 25835 4273
rect 25777 4233 25789 4267
rect 25823 4264 25835 4267
rect 26329 4267 26387 4273
rect 25823 4236 26234 4264
rect 25823 4233 25835 4236
rect 25777 4227 25835 4233
rect 13078 4156 13084 4208
rect 13136 4156 13142 4208
rect 24026 4196 24032 4208
rect 20640 4168 22508 4196
rect 23414 4168 24032 4196
rect 13078 4153 13136 4156
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8352 4100 8401 4128
rect 8352 4088 8358 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 12802 4088 12808 4140
rect 12860 4088 12866 4140
rect 13078 4119 13090 4153
rect 13124 4119 13136 4153
rect 20640 4140 20668 4168
rect 13078 4113 13136 4119
rect 20438 4088 20444 4140
rect 20496 4088 20502 4140
rect 20622 4088 20628 4140
rect 20680 4088 20686 4140
rect 22480 4137 22508 4168
rect 24026 4156 24032 4168
rect 24084 4156 24090 4208
rect 25148 4196 25176 4224
rect 25148 4168 25452 4196
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4097 21971 4131
rect 21913 4091 21971 4097
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4128 22523 4131
rect 25317 4131 25375 4137
rect 25317 4128 25329 4131
rect 22511 4100 25329 4128
rect 22511 4097 22523 4100
rect 22465 4091 22523 4097
rect 25317 4097 25329 4100
rect 25363 4097 25375 4131
rect 25424 4128 25452 4168
rect 25866 4156 25872 4208
rect 25924 4156 25930 4208
rect 25608 4137 25728 4138
rect 25495 4131 25553 4137
rect 25495 4128 25507 4131
rect 25424 4100 25507 4128
rect 25317 4091 25375 4097
rect 25495 4097 25507 4100
rect 25541 4097 25553 4131
rect 25495 4091 25553 4097
rect 25593 4131 25728 4137
rect 25593 4097 25605 4131
rect 25639 4110 25728 4131
rect 25639 4097 25651 4110
rect 25593 4091 25651 4097
rect 20456 4060 20484 4088
rect 21928 4060 21956 4091
rect 20456 4032 21956 4060
rect 25332 4060 25360 4091
rect 25700 4060 25728 4110
rect 25785 4121 25843 4127
rect 25785 4087 25797 4121
rect 25831 4118 25843 4121
rect 25884 4118 25912 4156
rect 25831 4090 25912 4118
rect 26053 4131 26111 4137
rect 26053 4097 26065 4131
rect 26099 4097 26111 4131
rect 26053 4091 26111 4097
rect 25831 4087 25843 4090
rect 25785 4081 25843 4087
rect 25958 4060 25964 4072
rect 25332 4052 25728 4060
rect 25884 4052 25964 4060
rect 25332 4032 25964 4052
rect 25700 4024 25912 4032
rect 25958 4020 25964 4032
rect 26016 4020 26022 4072
rect 24026 3952 24032 4004
rect 24084 3992 24090 4004
rect 25498 3992 25504 4004
rect 24084 3964 25504 3992
rect 24084 3952 24090 3964
rect 25498 3952 25504 3964
rect 25556 3992 25562 4004
rect 26068 3992 26096 4091
rect 25556 3964 26096 3992
rect 26206 3992 26234 4236
rect 26329 4233 26341 4267
rect 26375 4264 26387 4267
rect 26786 4264 26792 4276
rect 26375 4236 26792 4264
rect 26375 4233 26387 4236
rect 26329 4227 26387 4233
rect 26786 4224 26792 4236
rect 26844 4224 26850 4276
rect 26973 4267 27031 4273
rect 26973 4233 26985 4267
rect 27019 4264 27031 4267
rect 27062 4264 27068 4276
rect 27019 4236 27068 4264
rect 27019 4233 27031 4236
rect 26973 4227 27031 4233
rect 27062 4224 27068 4236
rect 27120 4224 27126 4276
rect 27430 4224 27436 4276
rect 27488 4224 27494 4276
rect 27890 4224 27896 4276
rect 27948 4224 27954 4276
rect 28074 4224 28080 4276
rect 28132 4264 28138 4276
rect 28132 4236 28488 4264
rect 28132 4224 28138 4236
rect 26418 4156 26424 4208
rect 26476 4156 26482 4208
rect 26510 4156 26516 4208
rect 26568 4196 26574 4208
rect 26697 4199 26755 4205
rect 26568 4168 26648 4196
rect 26568 4156 26574 4168
rect 26329 4063 26387 4069
rect 26329 4029 26341 4063
rect 26375 4060 26387 4063
rect 26436 4060 26464 4156
rect 26620 4137 26648 4168
rect 26697 4165 26709 4199
rect 26743 4196 26755 4199
rect 27448 4196 27476 4224
rect 26743 4168 27476 4196
rect 26743 4165 26755 4168
rect 26697 4159 26755 4165
rect 27706 4156 27712 4208
rect 27764 4196 27770 4208
rect 27801 4199 27859 4205
rect 27801 4196 27813 4199
rect 27764 4168 27813 4196
rect 27764 4156 27770 4168
rect 27801 4165 27813 4168
rect 27847 4165 27859 4199
rect 27908 4196 27936 4224
rect 28460 4196 28488 4236
rect 28534 4224 28540 4276
rect 28592 4224 28598 4276
rect 27908 4168 28120 4196
rect 28460 4168 28672 4196
rect 27801 4159 27859 4165
rect 26605 4131 26663 4137
rect 26605 4097 26617 4131
rect 26651 4097 26663 4131
rect 26605 4091 26663 4097
rect 26789 4131 26847 4137
rect 26789 4097 26801 4131
rect 26835 4128 26847 4131
rect 27341 4131 27399 4137
rect 27341 4128 27353 4131
rect 26835 4100 27353 4128
rect 26835 4097 26847 4100
rect 26789 4091 26847 4097
rect 27341 4097 27353 4100
rect 27387 4097 27399 4131
rect 27341 4091 27399 4097
rect 27617 4131 27675 4137
rect 27617 4097 27629 4131
rect 27663 4128 27675 4131
rect 27982 4128 27988 4140
rect 27663 4100 27988 4128
rect 27663 4097 27675 4100
rect 27617 4091 27675 4097
rect 26375 4032 26464 4060
rect 26375 4029 26387 4032
rect 26329 4023 26387 4029
rect 26804 3992 26832 4091
rect 27982 4088 27988 4100
rect 28040 4088 28046 4140
rect 28092 4137 28120 4168
rect 28077 4131 28135 4137
rect 28077 4097 28089 4131
rect 28123 4097 28135 4131
rect 28077 4091 28135 4097
rect 28166 4088 28172 4140
rect 28224 4128 28230 4140
rect 28644 4137 28672 4168
rect 28445 4131 28503 4137
rect 28445 4128 28457 4131
rect 28224 4100 28457 4128
rect 28224 4088 28230 4100
rect 28445 4097 28457 4100
rect 28491 4097 28503 4131
rect 28445 4091 28503 4097
rect 28629 4131 28687 4137
rect 28629 4097 28641 4131
rect 28675 4128 28687 4131
rect 29546 4128 29552 4140
rect 28675 4100 29552 4128
rect 28675 4097 28687 4100
rect 28629 4091 28687 4097
rect 29546 4088 29552 4100
rect 29604 4088 29610 4140
rect 26878 4020 26884 4072
rect 26936 4060 26942 4072
rect 27433 4063 27491 4069
rect 27433 4060 27445 4063
rect 26936 4032 27445 4060
rect 26936 4020 26942 4032
rect 27433 4029 27445 4032
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 26206 3964 26832 3992
rect 25556 3952 25562 3964
rect 27338 3952 27344 4004
rect 27396 3952 27402 4004
rect 22922 3884 22928 3936
rect 22980 3924 22986 3936
rect 26145 3927 26203 3933
rect 26145 3924 26157 3927
rect 22980 3896 26157 3924
rect 22980 3884 22986 3896
rect 26145 3893 26157 3896
rect 26191 3924 26203 3927
rect 27356 3924 27384 3952
rect 26191 3896 27384 3924
rect 27801 3927 27859 3933
rect 26191 3893 26203 3896
rect 26145 3887 26203 3893
rect 27801 3893 27813 3927
rect 27847 3924 27859 3927
rect 28626 3924 28632 3936
rect 27847 3896 28632 3924
rect 27847 3893 27859 3896
rect 27801 3887 27859 3893
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 1104 3834 38272 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38272 3834
rect 1104 3760 38272 3782
rect 1104 3290 38272 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38272 3290
rect 1104 3216 38272 3238
rect 16482 3136 16488 3188
rect 16540 3136 16546 3188
rect 17678 3136 17684 3188
rect 17736 3136 17742 3188
rect 36906 3136 36912 3188
rect 36964 3136 36970 3188
rect 11790 3000 11796 3052
rect 11848 3000 11854 3052
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3040 16451 3043
rect 16500 3040 16528 3136
rect 16439 3012 16528 3040
rect 17589 3043 17647 3049
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 17589 3009 17601 3043
rect 17635 3040 17647 3043
rect 17696 3040 17724 3136
rect 17635 3012 17724 3040
rect 24581 3043 24639 3049
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 24581 3009 24593 3043
rect 24627 3040 24639 3043
rect 25406 3040 25412 3052
rect 24627 3012 25412 3040
rect 24627 3009 24639 3012
rect 24581 3003 24639 3009
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 36924 3040 36952 3136
rect 37093 3043 37151 3049
rect 37093 3040 37105 3043
rect 36924 3012 37105 3040
rect 37093 3009 37105 3012
rect 37139 3009 37151 3043
rect 37093 3003 37151 3009
rect 37553 3043 37611 3049
rect 37553 3009 37565 3043
rect 37599 3009 37611 3043
rect 37553 3003 37611 3009
rect 37568 2972 37596 3003
rect 36924 2944 37596 2972
rect 36924 2913 36952 2944
rect 36909 2907 36967 2913
rect 36909 2873 36921 2907
rect 36955 2873 36967 2907
rect 36909 2867 36967 2873
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 8260 2808 11621 2836
rect 8260 2796 8266 2808
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 11609 2799 11667 2805
rect 12986 2796 12992 2848
rect 13044 2796 13050 2848
rect 16206 2796 16212 2848
rect 16264 2796 16270 2848
rect 17402 2796 17408 2848
rect 17460 2796 17466 2848
rect 21910 2796 21916 2848
rect 21968 2836 21974 2848
rect 24397 2839 24455 2845
rect 24397 2836 24409 2839
rect 21968 2808 24409 2836
rect 21968 2796 21974 2808
rect 24397 2805 24409 2808
rect 24443 2805 24455 2839
rect 24397 2799 24455 2805
rect 37182 2796 37188 2848
rect 37240 2836 37246 2848
rect 37645 2839 37703 2845
rect 37645 2836 37657 2839
rect 37240 2808 37657 2836
rect 37240 2796 37246 2808
rect 37645 2805 37657 2808
rect 37691 2805 37703 2839
rect 37645 2799 37703 2805
rect 1104 2746 38272 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38272 2746
rect 1104 2672 38272 2694
rect 8662 2592 8668 2644
rect 8720 2592 8726 2644
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 37645 2567 37703 2573
rect 37645 2564 37657 2567
rect 26206 2536 37657 2564
rect 10226 2456 10232 2508
rect 10284 2496 10290 2508
rect 26206 2496 26234 2536
rect 37645 2533 37657 2536
rect 37691 2533 37703 2567
rect 37645 2527 37703 2533
rect 10284 2468 26234 2496
rect 10284 2456 10290 2468
rect 1486 2388 1492 2440
rect 1544 2388 1550 2440
rect 2130 2388 2136 2440
rect 2188 2388 2194 2440
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 8202 2428 8208 2440
rect 6687 2400 8208 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 9640 2400 11284 2428
rect 9640 2388 9646 2400
rect 11146 2320 11152 2372
rect 11204 2320 11210 2372
rect 11256 2360 11284 2400
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 13044 2400 13093 2428
rect 13044 2388 13050 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 16206 2428 16212 2440
rect 15059 2400 16212 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 16206 2388 16212 2400
rect 16264 2388 16270 2440
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17460 2400 17601 2428
rect 17460 2388 17466 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 21910 2428 21916 2440
rect 19567 2400 21916 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 21910 2388 21916 2400
rect 21968 2388 21974 2440
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 27065 2363 27123 2369
rect 27065 2360 27077 2363
rect 11256 2332 27077 2360
rect 27065 2329 27077 2332
rect 27111 2329 27123 2363
rect 27065 2323 27123 2329
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 72 2264 1593 2292
rect 72 2252 78 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 2004 2264 2237 2292
rect 2004 2252 2010 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 3970 2252 3976 2304
rect 4028 2292 4034 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 4028 2264 4169 2292
rect 4028 2252 4034 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 6880 2264 6929 2292
rect 6880 2252 6886 2264
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 6917 2255 6975 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 15068 2264 15301 2292
rect 15068 2252 15074 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26476 2264 27169 2292
rect 26476 2252 26482 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 1104 2202 38272 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38272 2202
rect 1104 2128 38272 2150
<< via1 >>
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 20 39040 72 39092
rect 4528 39040 4580 39092
rect 9036 39040 9088 39092
rect 11060 39040 11112 39092
rect 12900 39040 12952 39092
rect 9128 38972 9180 39024
rect 17408 39040 17460 39092
rect 21916 39040 21968 39092
rect 26424 39040 26476 39092
rect 32864 39040 32916 39092
rect 15476 38972 15528 39024
rect 16028 38972 16080 39024
rect 3792 38904 3844 38956
rect 4804 38947 4856 38956
rect 4804 38913 4813 38947
rect 4813 38913 4847 38947
rect 4847 38913 4856 38947
rect 4804 38904 4856 38913
rect 9312 38947 9364 38956
rect 9312 38913 9321 38947
rect 9321 38913 9355 38947
rect 9355 38913 9364 38947
rect 9312 38904 9364 38913
rect 11612 38947 11664 38956
rect 11612 38913 11621 38947
rect 11621 38913 11655 38947
rect 11655 38913 11664 38947
rect 11612 38904 11664 38913
rect 11980 38904 12032 38956
rect 12716 38947 12768 38956
rect 12716 38913 12725 38947
rect 12725 38913 12759 38947
rect 12759 38913 12768 38947
rect 12716 38904 12768 38913
rect 12992 38947 13044 38956
rect 12992 38913 13001 38947
rect 13001 38913 13035 38947
rect 13035 38913 13044 38947
rect 12992 38904 13044 38913
rect 24400 38972 24452 39024
rect 30932 38972 30984 39024
rect 35900 38972 35952 39024
rect 19984 38904 20036 38956
rect 22100 38947 22152 38956
rect 22100 38913 22109 38947
rect 22109 38913 22143 38947
rect 22143 38913 22152 38947
rect 22100 38904 22152 38913
rect 24768 38947 24820 38956
rect 24768 38913 24777 38947
rect 24777 38913 24811 38947
rect 24811 38913 24820 38947
rect 24768 38904 24820 38913
rect 25044 38904 25096 38956
rect 27068 38947 27120 38956
rect 27068 38913 27077 38947
rect 27077 38913 27111 38947
rect 27111 38913 27120 38947
rect 27068 38904 27120 38913
rect 33048 38947 33100 38956
rect 33048 38913 33057 38947
rect 33057 38913 33091 38947
rect 33091 38913 33100 38947
rect 33048 38904 33100 38913
rect 35624 38947 35676 38956
rect 35624 38913 35633 38947
rect 35633 38913 35667 38947
rect 35667 38913 35676 38947
rect 35624 38904 35676 38913
rect 37372 38904 37424 38956
rect 11244 38836 11296 38888
rect 26148 38879 26200 38888
rect 26148 38845 26157 38879
rect 26157 38845 26191 38879
rect 26191 38845 26200 38879
rect 26148 38836 26200 38845
rect 10232 38768 10284 38820
rect 12348 38743 12400 38752
rect 12348 38709 12357 38743
rect 12357 38709 12391 38743
rect 12391 38709 12400 38743
rect 12348 38700 12400 38709
rect 12440 38700 12492 38752
rect 16028 38768 16080 38820
rect 24952 38700 25004 38752
rect 31208 38743 31260 38752
rect 31208 38709 31217 38743
rect 31217 38709 31251 38743
rect 31251 38709 31260 38743
rect 31208 38700 31260 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 4804 38496 4856 38548
rect 9312 38539 9364 38548
rect 9312 38505 9321 38539
rect 9321 38505 9355 38539
rect 9355 38505 9364 38539
rect 9312 38496 9364 38505
rect 12440 38496 12492 38548
rect 17500 38496 17552 38548
rect 22652 38496 22704 38548
rect 24400 38539 24452 38548
rect 24400 38505 24409 38539
rect 24409 38505 24443 38539
rect 24443 38505 24452 38539
rect 24400 38496 24452 38505
rect 12348 38360 12400 38412
rect 14464 38360 14516 38412
rect 20904 38360 20956 38412
rect 5172 38335 5224 38344
rect 5172 38301 5181 38335
rect 5181 38301 5215 38335
rect 5215 38301 5224 38335
rect 5172 38292 5224 38301
rect 9496 38335 9548 38344
rect 9496 38301 9505 38335
rect 9505 38301 9539 38335
rect 9539 38301 9548 38335
rect 9496 38292 9548 38301
rect 20168 38335 20220 38344
rect 20168 38301 20177 38335
rect 20177 38301 20211 38335
rect 20211 38301 20220 38335
rect 20168 38292 20220 38301
rect 24400 38360 24452 38412
rect 10416 38267 10468 38276
rect 10416 38233 10425 38267
rect 10425 38233 10459 38267
rect 10459 38233 10468 38267
rect 10416 38224 10468 38233
rect 7104 38156 7156 38208
rect 8576 38199 8628 38208
rect 8576 38165 8585 38199
rect 8585 38165 8619 38199
rect 8619 38165 8628 38199
rect 8576 38156 8628 38165
rect 10600 38156 10652 38208
rect 11888 38199 11940 38208
rect 11888 38165 11897 38199
rect 11897 38165 11931 38199
rect 11931 38165 11940 38199
rect 11888 38156 11940 38165
rect 11980 38156 12032 38208
rect 14004 38224 14056 38276
rect 22560 38335 22612 38344
rect 22560 38301 22569 38335
rect 22569 38301 22603 38335
rect 22603 38301 22612 38335
rect 25044 38496 25096 38548
rect 24952 38360 25004 38412
rect 26148 38360 26200 38412
rect 27896 38496 27948 38548
rect 30288 38496 30340 38548
rect 33048 38496 33100 38548
rect 35624 38496 35676 38548
rect 37924 38496 37976 38548
rect 27344 38360 27396 38412
rect 27620 38360 27672 38412
rect 22560 38292 22612 38301
rect 13728 38156 13780 38208
rect 16212 38156 16264 38208
rect 18696 38156 18748 38208
rect 19892 38156 19944 38208
rect 24860 38224 24912 38276
rect 24952 38267 25004 38276
rect 24952 38233 24961 38267
rect 24961 38233 24995 38267
rect 24995 38233 25004 38267
rect 24952 38224 25004 38233
rect 22284 38199 22336 38208
rect 22284 38165 22293 38199
rect 22293 38165 22327 38199
rect 22327 38165 22336 38199
rect 22284 38156 22336 38165
rect 24768 38156 24820 38208
rect 26424 38199 26476 38208
rect 26424 38165 26433 38199
rect 26433 38165 26467 38199
rect 26467 38165 26476 38199
rect 26424 38156 26476 38165
rect 27252 38267 27304 38276
rect 27252 38233 27261 38267
rect 27261 38233 27295 38267
rect 27295 38233 27304 38267
rect 27252 38224 27304 38233
rect 27344 38224 27396 38276
rect 27620 38156 27672 38208
rect 31208 38292 31260 38344
rect 29828 38267 29880 38276
rect 29828 38233 29837 38267
rect 29837 38233 29871 38267
rect 29871 38233 29880 38267
rect 29828 38224 29880 38233
rect 30288 38224 30340 38276
rect 32036 38292 32088 38344
rect 34520 38292 34572 38344
rect 29276 38156 29328 38208
rect 31944 38199 31996 38208
rect 31944 38165 31953 38199
rect 31953 38165 31987 38199
rect 31987 38165 31996 38199
rect 31944 38156 31996 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 8576 37952 8628 38004
rect 10416 37952 10468 38004
rect 10784 37952 10836 38004
rect 10600 37884 10652 37936
rect 8668 37791 8720 37800
rect 8668 37757 8677 37791
rect 8677 37757 8711 37791
rect 8711 37757 8720 37791
rect 8668 37748 8720 37757
rect 11152 37791 11204 37800
rect 11152 37757 11161 37791
rect 11161 37757 11195 37791
rect 11195 37757 11204 37791
rect 11152 37748 11204 37757
rect 11612 37952 11664 38004
rect 12716 37952 12768 38004
rect 13728 37952 13780 38004
rect 13084 37884 13136 37936
rect 11704 37859 11756 37868
rect 11704 37825 11713 37859
rect 11713 37825 11747 37859
rect 11747 37825 11756 37859
rect 11704 37816 11756 37825
rect 14464 37952 14516 38004
rect 14556 37952 14608 38004
rect 14280 37859 14332 37868
rect 14280 37825 14289 37859
rect 14289 37825 14323 37859
rect 14323 37825 14332 37859
rect 14280 37816 14332 37825
rect 14372 37816 14424 37868
rect 11888 37680 11940 37732
rect 12348 37680 12400 37732
rect 17500 37927 17552 37936
rect 17500 37893 17509 37927
rect 17509 37893 17543 37927
rect 17543 37893 17552 37927
rect 17500 37884 17552 37893
rect 17684 37952 17736 38004
rect 17868 37995 17920 38004
rect 17868 37961 17877 37995
rect 17877 37961 17911 37995
rect 17911 37961 17920 37995
rect 17868 37952 17920 37961
rect 18696 37952 18748 38004
rect 18788 37952 18840 38004
rect 14832 37816 14884 37868
rect 15752 37816 15804 37868
rect 15936 37859 15988 37868
rect 15936 37825 15945 37859
rect 15945 37825 15979 37859
rect 15979 37825 15988 37859
rect 15936 37816 15988 37825
rect 16028 37859 16080 37868
rect 16028 37825 16037 37859
rect 16037 37825 16071 37859
rect 16071 37825 16080 37859
rect 16028 37816 16080 37825
rect 18144 37816 18196 37868
rect 18512 37816 18564 37868
rect 18880 37816 18932 37868
rect 19064 37859 19116 37868
rect 19064 37825 19073 37859
rect 19073 37825 19107 37859
rect 19107 37825 19116 37859
rect 19064 37816 19116 37825
rect 19156 37859 19208 37868
rect 19156 37825 19165 37859
rect 19165 37825 19199 37859
rect 19199 37825 19208 37859
rect 19156 37816 19208 37825
rect 20168 37952 20220 38004
rect 22192 37952 22244 38004
rect 22652 37952 22704 38004
rect 23940 37952 23992 38004
rect 24952 37952 25004 38004
rect 19984 37884 20036 37936
rect 20168 37816 20220 37868
rect 22284 37884 22336 37936
rect 26424 37952 26476 38004
rect 27252 37952 27304 38004
rect 22008 37859 22060 37868
rect 22008 37825 22017 37859
rect 22017 37825 22051 37859
rect 22051 37825 22060 37859
rect 22008 37816 22060 37825
rect 22468 37816 22520 37868
rect 22652 37816 22704 37868
rect 22836 37859 22888 37868
rect 22836 37825 22845 37859
rect 22845 37825 22879 37859
rect 22879 37825 22888 37859
rect 22836 37816 22888 37825
rect 22928 37859 22980 37868
rect 22928 37825 22937 37859
rect 22937 37825 22971 37859
rect 22971 37825 22980 37859
rect 22928 37816 22980 37825
rect 20904 37791 20956 37800
rect 20904 37757 20913 37791
rect 20913 37757 20947 37791
rect 20947 37757 20956 37791
rect 20904 37748 20956 37757
rect 20996 37791 21048 37800
rect 20996 37757 21005 37791
rect 21005 37757 21039 37791
rect 21039 37757 21048 37791
rect 20996 37748 21048 37757
rect 29276 37995 29328 38004
rect 29276 37961 29285 37995
rect 29285 37961 29319 37995
rect 29319 37961 29328 37995
rect 29276 37952 29328 37961
rect 29828 37952 29880 38004
rect 21548 37680 21600 37732
rect 22836 37680 22888 37732
rect 24952 37859 25004 37868
rect 24952 37825 24961 37859
rect 24961 37825 24995 37859
rect 24995 37825 25004 37859
rect 24952 37816 25004 37825
rect 25228 37859 25280 37868
rect 25228 37825 25237 37859
rect 25237 37825 25271 37859
rect 25271 37825 25280 37859
rect 25228 37816 25280 37825
rect 25412 37859 25464 37868
rect 25412 37825 25421 37859
rect 25421 37825 25455 37859
rect 25455 37825 25464 37859
rect 25412 37816 25464 37825
rect 25228 37680 25280 37732
rect 26976 37748 27028 37800
rect 27344 37816 27396 37868
rect 27988 37859 28040 37868
rect 27988 37825 27997 37859
rect 27997 37825 28031 37859
rect 28031 37825 28040 37859
rect 27988 37816 28040 37825
rect 27528 37791 27580 37800
rect 10140 37655 10192 37664
rect 10140 37621 10149 37655
rect 10149 37621 10183 37655
rect 10183 37621 10192 37655
rect 10140 37612 10192 37621
rect 15200 37612 15252 37664
rect 19340 37655 19392 37664
rect 19340 37621 19349 37655
rect 19349 37621 19383 37655
rect 19383 37621 19392 37655
rect 19340 37612 19392 37621
rect 19800 37655 19852 37664
rect 19800 37621 19809 37655
rect 19809 37621 19843 37655
rect 19843 37621 19852 37655
rect 19800 37612 19852 37621
rect 22100 37612 22152 37664
rect 22376 37655 22428 37664
rect 22376 37621 22385 37655
rect 22385 37621 22419 37655
rect 22419 37621 22428 37655
rect 22376 37612 22428 37621
rect 23112 37655 23164 37664
rect 23112 37621 23121 37655
rect 23121 37621 23155 37655
rect 23155 37621 23164 37655
rect 23112 37612 23164 37621
rect 24768 37612 24820 37664
rect 25412 37612 25464 37664
rect 26240 37612 26292 37664
rect 27528 37757 27537 37791
rect 27537 37757 27571 37791
rect 27571 37757 27580 37791
rect 27528 37748 27580 37757
rect 27804 37748 27856 37800
rect 29184 37859 29236 37868
rect 29184 37825 29193 37859
rect 29193 37825 29227 37859
rect 29227 37825 29236 37859
rect 29184 37816 29236 37825
rect 31944 37952 31996 38004
rect 30288 37884 30340 37936
rect 32312 37859 32364 37868
rect 32312 37825 32321 37859
rect 32321 37825 32355 37859
rect 32355 37825 32364 37859
rect 32312 37816 32364 37825
rect 27528 37612 27580 37664
rect 32036 37680 32088 37732
rect 31760 37655 31812 37664
rect 31760 37621 31769 37655
rect 31769 37621 31803 37655
rect 31803 37621 31812 37655
rect 31760 37612 31812 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 8668 37408 8720 37460
rect 16028 37408 16080 37460
rect 17868 37408 17920 37460
rect 23112 37408 23164 37460
rect 24860 37408 24912 37460
rect 11152 37340 11204 37392
rect 13268 37340 13320 37392
rect 15936 37340 15988 37392
rect 6460 37272 6512 37324
rect 10048 37315 10100 37324
rect 10048 37281 10057 37315
rect 10057 37281 10091 37315
rect 10091 37281 10100 37315
rect 10048 37272 10100 37281
rect 10140 37272 10192 37324
rect 18236 37340 18288 37392
rect 19064 37340 19116 37392
rect 25044 37340 25096 37392
rect 27068 37340 27120 37392
rect 940 37136 992 37188
rect 14280 37247 14332 37256
rect 14280 37213 14289 37247
rect 14289 37213 14323 37247
rect 14323 37213 14332 37247
rect 14280 37204 14332 37213
rect 18052 37272 18104 37324
rect 19340 37272 19392 37324
rect 19800 37204 19852 37256
rect 21548 37204 21600 37256
rect 21824 37204 21876 37256
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 22100 37247 22152 37256
rect 22100 37213 22109 37247
rect 22109 37213 22143 37247
rect 22143 37213 22152 37247
rect 22100 37204 22152 37213
rect 24676 37272 24728 37324
rect 26976 37315 27028 37324
rect 26976 37281 26985 37315
rect 26985 37281 27019 37315
rect 27019 37281 27028 37315
rect 26976 37272 27028 37281
rect 15108 37179 15160 37188
rect 15108 37145 15117 37179
rect 15117 37145 15151 37179
rect 15151 37145 15160 37179
rect 15108 37136 15160 37145
rect 19432 37179 19484 37188
rect 19432 37145 19441 37179
rect 19441 37145 19475 37179
rect 19475 37145 19484 37179
rect 19432 37136 19484 37145
rect 22376 37204 22428 37256
rect 22652 37247 22704 37256
rect 22652 37213 22662 37247
rect 22662 37213 22696 37247
rect 22696 37213 22704 37247
rect 22652 37204 22704 37213
rect 23112 37204 23164 37256
rect 11796 37068 11848 37120
rect 15936 37068 15988 37120
rect 18788 37068 18840 37120
rect 19156 37068 19208 37120
rect 22836 37179 22888 37188
rect 22836 37145 22845 37179
rect 22845 37145 22879 37179
rect 22879 37145 22888 37179
rect 22836 37136 22888 37145
rect 22928 37179 22980 37188
rect 22928 37145 22937 37179
rect 22937 37145 22971 37179
rect 22971 37145 22980 37179
rect 22928 37136 22980 37145
rect 23848 37247 23900 37256
rect 23848 37213 23857 37247
rect 23857 37213 23891 37247
rect 23891 37213 23900 37247
rect 23848 37204 23900 37213
rect 25228 37204 25280 37256
rect 27804 37272 27856 37324
rect 29184 37272 29236 37324
rect 31208 37315 31260 37324
rect 31208 37281 31217 37315
rect 31217 37281 31251 37315
rect 31251 37281 31260 37315
rect 31208 37272 31260 37281
rect 31300 37315 31352 37324
rect 31300 37281 31309 37315
rect 31309 37281 31343 37315
rect 31343 37281 31352 37315
rect 31300 37272 31352 37281
rect 20076 37068 20128 37120
rect 23572 37179 23624 37188
rect 23572 37145 23581 37179
rect 23581 37145 23615 37179
rect 23615 37145 23624 37179
rect 23572 37136 23624 37145
rect 34520 37204 34572 37256
rect 23204 37111 23256 37120
rect 23204 37077 23213 37111
rect 23213 37077 23247 37111
rect 23247 37077 23256 37111
rect 23204 37068 23256 37077
rect 23664 37068 23716 37120
rect 25872 37068 25924 37120
rect 32312 37136 32364 37188
rect 37280 37179 37332 37188
rect 37280 37145 37289 37179
rect 37289 37145 37323 37179
rect 37323 37145 37332 37179
rect 37280 37136 37332 37145
rect 31116 37111 31168 37120
rect 31116 37077 31125 37111
rect 31125 37077 31159 37111
rect 31159 37077 31168 37111
rect 31116 37068 31168 37077
rect 31208 37068 31260 37120
rect 33140 37068 33192 37120
rect 37832 37111 37884 37120
rect 37832 37077 37841 37111
rect 37841 37077 37875 37111
rect 37875 37077 37884 37111
rect 37832 37068 37884 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 18236 36864 18288 36916
rect 22652 36864 22704 36916
rect 23848 36864 23900 36916
rect 24400 36864 24452 36916
rect 28264 36864 28316 36916
rect 31760 36864 31812 36916
rect 18880 36796 18932 36848
rect 21456 36796 21508 36848
rect 21916 36796 21968 36848
rect 15844 36728 15896 36780
rect 16212 36771 16264 36780
rect 16212 36737 16221 36771
rect 16221 36737 16255 36771
rect 16255 36737 16264 36771
rect 16212 36728 16264 36737
rect 16304 36771 16356 36780
rect 16304 36737 16318 36771
rect 16318 36737 16352 36771
rect 16352 36737 16356 36771
rect 16304 36728 16356 36737
rect 20168 36728 20220 36780
rect 24952 36796 25004 36848
rect 7104 36660 7156 36712
rect 17224 36660 17276 36712
rect 20444 36660 20496 36712
rect 25320 36728 25372 36780
rect 25964 36728 26016 36780
rect 26148 36728 26200 36780
rect 29736 36796 29788 36848
rect 31116 36796 31168 36848
rect 32956 36771 33008 36780
rect 32956 36737 32965 36771
rect 32965 36737 32999 36771
rect 32999 36737 33008 36771
rect 32956 36728 33008 36737
rect 28724 36660 28776 36712
rect 11796 36592 11848 36644
rect 22928 36592 22980 36644
rect 24584 36592 24636 36644
rect 26792 36592 26844 36644
rect 30012 36592 30064 36644
rect 7012 36524 7064 36576
rect 15292 36524 15344 36576
rect 16212 36524 16264 36576
rect 18512 36524 18564 36576
rect 19892 36524 19944 36576
rect 20352 36524 20404 36576
rect 20904 36524 20956 36576
rect 21916 36524 21968 36576
rect 25688 36524 25740 36576
rect 25780 36567 25832 36576
rect 25780 36533 25789 36567
rect 25789 36533 25823 36567
rect 25823 36533 25832 36567
rect 25780 36524 25832 36533
rect 27436 36524 27488 36576
rect 32772 36567 32824 36576
rect 32772 36533 32781 36567
rect 32781 36533 32815 36567
rect 32815 36533 32824 36567
rect 32772 36524 32824 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 7012 36320 7064 36372
rect 17500 36320 17552 36372
rect 18328 36320 18380 36372
rect 18420 36320 18472 36372
rect 19432 36320 19484 36372
rect 22468 36320 22520 36372
rect 23296 36320 23348 36372
rect 23572 36320 23624 36372
rect 25044 36320 25096 36372
rect 26240 36320 26292 36372
rect 26424 36320 26476 36372
rect 26792 36320 26844 36372
rect 10692 36227 10744 36236
rect 10692 36193 10701 36227
rect 10701 36193 10735 36227
rect 10735 36193 10744 36227
rect 10692 36184 10744 36193
rect 8944 36159 8996 36168
rect 8944 36125 8953 36159
rect 8953 36125 8987 36159
rect 8987 36125 8996 36159
rect 8944 36116 8996 36125
rect 5540 36048 5592 36100
rect 6828 36048 6880 36100
rect 7196 36091 7248 36100
rect 7196 36057 7205 36091
rect 7205 36057 7239 36091
rect 7239 36057 7248 36091
rect 7196 36048 7248 36057
rect 8484 36048 8536 36100
rect 5356 35980 5408 36032
rect 6736 36023 6788 36032
rect 6736 35989 6745 36023
rect 6745 35989 6779 36023
rect 6779 35989 6788 36023
rect 6736 35980 6788 35989
rect 8668 36023 8720 36032
rect 8668 35989 8677 36023
rect 8677 35989 8711 36023
rect 8711 35989 8720 36023
rect 8668 35980 8720 35989
rect 9220 36091 9272 36100
rect 9220 36057 9229 36091
rect 9229 36057 9263 36091
rect 9263 36057 9272 36091
rect 9220 36048 9272 36057
rect 10600 36116 10652 36168
rect 12348 36116 12400 36168
rect 12624 36159 12676 36168
rect 12624 36125 12633 36159
rect 12633 36125 12667 36159
rect 12667 36125 12676 36159
rect 12624 36116 12676 36125
rect 12808 36116 12860 36168
rect 13636 36159 13688 36168
rect 13636 36125 13645 36159
rect 13645 36125 13679 36159
rect 13679 36125 13688 36159
rect 13636 36116 13688 36125
rect 17132 36184 17184 36236
rect 15200 36159 15252 36168
rect 15200 36125 15209 36159
rect 15209 36125 15243 36159
rect 15243 36125 15252 36159
rect 15200 36116 15252 36125
rect 15292 36159 15344 36168
rect 15292 36125 15301 36159
rect 15301 36125 15335 36159
rect 15335 36125 15344 36159
rect 15292 36116 15344 36125
rect 15568 36159 15620 36168
rect 15568 36125 15577 36159
rect 15577 36125 15611 36159
rect 15611 36125 15620 36159
rect 15568 36116 15620 36125
rect 17776 36252 17828 36304
rect 18604 36252 18656 36304
rect 18328 36184 18380 36236
rect 18696 36184 18748 36236
rect 17684 36159 17736 36168
rect 17684 36125 17693 36159
rect 17693 36125 17727 36159
rect 17727 36125 17736 36159
rect 17684 36116 17736 36125
rect 17776 36159 17828 36168
rect 17776 36125 17785 36159
rect 17785 36125 17819 36159
rect 17819 36125 17828 36159
rect 17776 36116 17828 36125
rect 18144 36116 18196 36168
rect 12440 36091 12492 36100
rect 12440 36057 12449 36091
rect 12449 36057 12483 36091
rect 12483 36057 12492 36091
rect 12440 36048 12492 36057
rect 14740 36048 14792 36100
rect 18512 36159 18564 36168
rect 18512 36125 18522 36159
rect 18522 36125 18556 36159
rect 18556 36125 18564 36159
rect 18512 36116 18564 36125
rect 18788 36159 18840 36168
rect 18788 36125 18797 36159
rect 18797 36125 18831 36159
rect 18831 36125 18840 36159
rect 18788 36116 18840 36125
rect 18880 36159 18932 36168
rect 18880 36125 18894 36159
rect 18894 36125 18928 36159
rect 18928 36125 18932 36159
rect 18880 36116 18932 36125
rect 12992 36023 13044 36032
rect 12992 35989 13001 36023
rect 13001 35989 13035 36023
rect 13035 35989 13044 36023
rect 12992 35980 13044 35989
rect 17408 35980 17460 36032
rect 18604 36048 18656 36100
rect 19340 36048 19392 36100
rect 19892 36116 19944 36168
rect 20352 36159 20404 36168
rect 20352 36125 20361 36159
rect 20361 36125 20395 36159
rect 20395 36125 20404 36159
rect 20352 36116 20404 36125
rect 20444 36116 20496 36168
rect 22100 36184 22152 36236
rect 20720 36159 20772 36168
rect 20720 36125 20729 36159
rect 20729 36125 20763 36159
rect 20763 36125 20772 36159
rect 20720 36116 20772 36125
rect 20352 35980 20404 36032
rect 22468 36116 22520 36168
rect 22652 36184 22704 36236
rect 22744 36116 22796 36168
rect 26056 36252 26108 36304
rect 21640 35980 21692 36032
rect 24124 36116 24176 36168
rect 24952 36116 25004 36168
rect 25320 36184 25372 36236
rect 25504 36159 25556 36168
rect 25504 36125 25513 36159
rect 25513 36125 25547 36159
rect 25547 36125 25556 36159
rect 25504 36116 25556 36125
rect 25964 36159 26016 36168
rect 25964 36125 25973 36159
rect 25973 36125 26007 36159
rect 26007 36125 26016 36159
rect 25964 36116 26016 36125
rect 26332 36159 26384 36168
rect 26332 36125 26341 36159
rect 26341 36125 26375 36159
rect 26375 36125 26384 36159
rect 26332 36116 26384 36125
rect 26424 36159 26476 36168
rect 26424 36125 26434 36159
rect 26434 36125 26468 36159
rect 26468 36125 26476 36159
rect 26424 36116 26476 36125
rect 25320 36048 25372 36100
rect 25136 35980 25188 36032
rect 25596 35980 25648 36032
rect 26056 36048 26108 36100
rect 26240 36048 26292 36100
rect 26516 36048 26568 36100
rect 29092 36320 29144 36372
rect 29368 36320 29420 36372
rect 27436 36252 27488 36304
rect 27804 36184 27856 36236
rect 29460 36252 29512 36304
rect 27436 36159 27488 36168
rect 27436 36125 27445 36159
rect 27445 36125 27479 36159
rect 27479 36125 27488 36159
rect 27436 36116 27488 36125
rect 26976 36023 27028 36032
rect 26976 35989 26985 36023
rect 26985 35989 27019 36023
rect 27019 35989 27028 36023
rect 26976 35980 27028 35989
rect 28264 36048 28316 36100
rect 28724 35980 28776 36032
rect 29276 36116 29328 36168
rect 29368 36116 29420 36168
rect 29736 36116 29788 36168
rect 30012 36159 30064 36168
rect 32772 36227 32824 36236
rect 32772 36193 32781 36227
rect 32781 36193 32815 36227
rect 32815 36193 32824 36227
rect 32772 36184 32824 36193
rect 30012 36125 30026 36159
rect 30026 36125 30060 36159
rect 30060 36125 30064 36159
rect 30012 36116 30064 36125
rect 30932 36159 30984 36168
rect 30932 36125 30941 36159
rect 30941 36125 30975 36159
rect 30975 36125 30984 36159
rect 30932 36116 30984 36125
rect 29368 35980 29420 36032
rect 30380 36023 30432 36032
rect 30380 35989 30389 36023
rect 30389 35989 30423 36023
rect 30423 35989 30432 36023
rect 30380 35980 30432 35989
rect 30748 36023 30800 36032
rect 30748 35989 30757 36023
rect 30757 35989 30791 36023
rect 30791 35989 30800 36023
rect 30748 35980 30800 35989
rect 32680 36048 32732 36100
rect 32772 35980 32824 36032
rect 34244 36023 34296 36032
rect 34244 35989 34253 36023
rect 34253 35989 34287 36023
rect 34287 35989 34296 36023
rect 34244 35980 34296 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 5540 35819 5592 35828
rect 5540 35785 5549 35819
rect 5549 35785 5583 35819
rect 5583 35785 5592 35819
rect 5540 35776 5592 35785
rect 7196 35776 7248 35828
rect 5632 35708 5684 35760
rect 6460 35708 6512 35760
rect 5724 35683 5776 35692
rect 5724 35649 5733 35683
rect 5733 35649 5767 35683
rect 5767 35649 5776 35683
rect 5724 35640 5776 35649
rect 8668 35776 8720 35828
rect 8944 35776 8996 35828
rect 9220 35776 9272 35828
rect 10692 35776 10744 35828
rect 13636 35776 13688 35828
rect 15568 35776 15620 35828
rect 17132 35776 17184 35828
rect 18696 35776 18748 35828
rect 6828 35572 6880 35624
rect 8484 35708 8536 35760
rect 11980 35751 12032 35760
rect 11980 35717 11989 35751
rect 11989 35717 12023 35751
rect 12023 35717 12032 35751
rect 11980 35708 12032 35717
rect 20904 35708 20956 35760
rect 22744 35776 22796 35828
rect 21640 35708 21692 35760
rect 21916 35708 21968 35760
rect 8944 35572 8996 35624
rect 9956 35640 10008 35692
rect 10784 35504 10836 35556
rect 8208 35436 8260 35488
rect 10600 35479 10652 35488
rect 10600 35445 10609 35479
rect 10609 35445 10643 35479
rect 10643 35445 10652 35479
rect 10600 35436 10652 35445
rect 11796 35640 11848 35692
rect 12808 35640 12860 35692
rect 12992 35683 13044 35692
rect 12992 35649 13002 35683
rect 13002 35649 13036 35683
rect 13036 35649 13044 35683
rect 12992 35640 13044 35649
rect 13176 35640 13228 35692
rect 13268 35683 13320 35692
rect 13268 35649 13277 35683
rect 13277 35649 13311 35683
rect 13311 35649 13320 35683
rect 13268 35640 13320 35649
rect 13360 35683 13412 35692
rect 13360 35649 13374 35683
rect 13374 35649 13408 35683
rect 13408 35649 13412 35683
rect 13360 35640 13412 35649
rect 14188 35640 14240 35692
rect 18604 35640 18656 35692
rect 21732 35640 21784 35692
rect 21824 35640 21876 35692
rect 22192 35640 22244 35692
rect 12256 35572 12308 35624
rect 22376 35683 22428 35692
rect 22376 35649 22385 35683
rect 22385 35649 22419 35683
rect 22419 35649 22428 35683
rect 22376 35640 22428 35649
rect 22560 35640 22612 35692
rect 22836 35683 22888 35692
rect 22836 35649 22846 35683
rect 22846 35649 22880 35683
rect 22880 35649 22888 35683
rect 22836 35640 22888 35649
rect 25780 35776 25832 35828
rect 27436 35776 27488 35828
rect 25596 35708 25648 35760
rect 26148 35708 26200 35760
rect 23572 35572 23624 35624
rect 25780 35683 25832 35692
rect 25780 35649 25789 35683
rect 25789 35649 25823 35683
rect 25823 35649 25832 35683
rect 25780 35640 25832 35649
rect 26056 35640 26108 35692
rect 26240 35640 26292 35692
rect 27344 35640 27396 35692
rect 27436 35572 27488 35624
rect 27804 35572 27856 35624
rect 29184 35640 29236 35692
rect 29460 35683 29512 35692
rect 29460 35649 29469 35683
rect 29469 35649 29503 35683
rect 29503 35649 29512 35683
rect 29460 35640 29512 35649
rect 29552 35640 29604 35692
rect 23112 35504 23164 35556
rect 24032 35504 24084 35556
rect 25320 35504 25372 35556
rect 25504 35504 25556 35556
rect 29000 35504 29052 35556
rect 12716 35436 12768 35488
rect 13360 35436 13412 35488
rect 21824 35436 21876 35488
rect 22376 35436 22428 35488
rect 22652 35479 22704 35488
rect 22652 35445 22661 35479
rect 22661 35445 22695 35479
rect 22695 35445 22704 35479
rect 22652 35436 22704 35445
rect 22744 35436 22796 35488
rect 23388 35479 23440 35488
rect 23388 35445 23397 35479
rect 23397 35445 23431 35479
rect 23431 35445 23440 35479
rect 23388 35436 23440 35445
rect 24584 35436 24636 35488
rect 26516 35436 26568 35488
rect 29276 35479 29328 35488
rect 29276 35445 29285 35479
rect 29285 35445 29319 35479
rect 29319 35445 29328 35479
rect 29276 35436 29328 35445
rect 29368 35436 29420 35488
rect 30380 35708 30432 35760
rect 30472 35708 30524 35760
rect 30840 35708 30892 35760
rect 30748 35572 30800 35624
rect 30840 35572 30892 35624
rect 32680 35776 32732 35828
rect 32956 35776 33008 35828
rect 33140 35819 33192 35828
rect 33140 35785 33149 35819
rect 33149 35785 33183 35819
rect 33183 35785 33192 35819
rect 33140 35776 33192 35785
rect 34244 35776 34296 35828
rect 33324 35615 33376 35624
rect 33324 35581 33333 35615
rect 33333 35581 33367 35615
rect 33367 35581 33376 35615
rect 33324 35572 33376 35581
rect 31852 35479 31904 35488
rect 31852 35445 31861 35479
rect 31861 35445 31895 35479
rect 31895 35445 31904 35479
rect 31852 35436 31904 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5724 35232 5776 35284
rect 8668 35232 8720 35284
rect 11888 35232 11940 35284
rect 11980 35275 12032 35284
rect 11980 35241 11989 35275
rect 11989 35241 12023 35275
rect 12023 35241 12032 35275
rect 11980 35232 12032 35241
rect 12072 35232 12124 35284
rect 17500 35164 17552 35216
rect 6552 35139 6604 35148
rect 6552 35105 6561 35139
rect 6561 35105 6595 35139
rect 6595 35105 6604 35139
rect 6552 35096 6604 35105
rect 10600 35096 10652 35148
rect 17408 35096 17460 35148
rect 20720 35164 20772 35216
rect 20904 35164 20956 35216
rect 5448 35028 5500 35080
rect 9956 35071 10008 35080
rect 9956 35037 9965 35071
rect 9965 35037 9999 35071
rect 9999 35037 10008 35071
rect 9956 35028 10008 35037
rect 14372 35028 14424 35080
rect 14832 35028 14884 35080
rect 6736 34960 6788 35012
rect 19340 35028 19392 35080
rect 19432 35071 19484 35080
rect 19432 35037 19441 35071
rect 19441 35037 19475 35071
rect 19475 35037 19484 35071
rect 19432 35028 19484 35037
rect 19984 35028 20036 35080
rect 20904 35028 20956 35080
rect 20996 35071 21048 35080
rect 20996 35037 21005 35071
rect 21005 35037 21039 35071
rect 21039 35037 21048 35071
rect 20996 35028 21048 35037
rect 22192 35232 22244 35284
rect 22652 35232 22704 35284
rect 27252 35232 27304 35284
rect 28264 35232 28316 35284
rect 30472 35232 30524 35284
rect 30932 35232 30984 35284
rect 4528 34935 4580 34944
rect 4528 34901 4537 34935
rect 4537 34901 4571 34935
rect 4571 34901 4580 34935
rect 4528 34892 4580 34901
rect 6460 34935 6512 34944
rect 6460 34901 6469 34935
rect 6469 34901 6503 34935
rect 6503 34901 6512 34935
rect 6460 34892 6512 34901
rect 8024 34935 8076 34944
rect 8024 34901 8033 34935
rect 8033 34901 8067 34935
rect 8067 34901 8076 34935
rect 8024 34892 8076 34901
rect 9404 34892 9456 34944
rect 10232 34892 10284 34944
rect 10692 34892 10744 34944
rect 10876 34892 10928 34944
rect 11980 34892 12032 34944
rect 14464 34892 14516 34944
rect 14648 34935 14700 34944
rect 14648 34901 14657 34935
rect 14657 34901 14691 34935
rect 14691 34901 14700 34935
rect 14648 34892 14700 34901
rect 15384 34892 15436 34944
rect 18236 34892 18288 34944
rect 21180 34960 21232 35012
rect 21272 35003 21324 35012
rect 21272 34969 21281 35003
rect 21281 34969 21315 35003
rect 21315 34969 21324 35003
rect 21272 34960 21324 34969
rect 21456 35071 21508 35080
rect 21456 35037 21470 35071
rect 21470 35037 21504 35071
rect 21504 35037 21508 35071
rect 21456 35028 21508 35037
rect 21640 35028 21692 35080
rect 22284 35071 22336 35080
rect 22284 35037 22294 35071
rect 22294 35037 22328 35071
rect 22328 35037 22336 35071
rect 23388 35164 23440 35216
rect 25412 35207 25464 35216
rect 25412 35173 25421 35207
rect 25421 35173 25455 35207
rect 25455 35173 25464 35207
rect 25412 35164 25464 35173
rect 25596 35164 25648 35216
rect 22284 35028 22336 35037
rect 23112 35028 23164 35080
rect 24216 35096 24268 35148
rect 23388 35071 23440 35080
rect 23388 35037 23397 35071
rect 23397 35037 23431 35071
rect 23431 35037 23440 35071
rect 23388 35028 23440 35037
rect 22928 34960 22980 35012
rect 19984 34892 20036 34944
rect 20720 34892 20772 34944
rect 24860 35028 24912 35080
rect 25136 35071 25188 35080
rect 25136 35037 25145 35071
rect 25145 35037 25179 35071
rect 25179 35037 25188 35071
rect 25136 35028 25188 35037
rect 25780 35071 25832 35080
rect 25780 35037 25789 35071
rect 25789 35037 25823 35071
rect 25823 35037 25832 35071
rect 25780 35028 25832 35037
rect 28264 35096 28316 35148
rect 31300 35139 31352 35148
rect 31300 35105 31309 35139
rect 31309 35105 31343 35139
rect 31343 35105 31352 35139
rect 31300 35096 31352 35105
rect 33692 35096 33744 35148
rect 25596 34960 25648 35012
rect 26976 35028 27028 35080
rect 27436 35028 27488 35080
rect 27712 35071 27764 35080
rect 27712 35037 27721 35071
rect 27721 35037 27755 35071
rect 27755 35037 27764 35071
rect 27712 35028 27764 35037
rect 29460 35028 29512 35080
rect 31852 35028 31904 35080
rect 22284 34892 22336 34944
rect 22836 34935 22888 34944
rect 22836 34901 22845 34935
rect 22845 34901 22879 34935
rect 22879 34901 22888 34935
rect 22836 34892 22888 34901
rect 23112 34935 23164 34944
rect 23112 34901 23121 34935
rect 23121 34901 23155 34935
rect 23155 34901 23164 34935
rect 23112 34892 23164 34901
rect 23204 34892 23256 34944
rect 23388 34892 23440 34944
rect 23756 34892 23808 34944
rect 24768 34892 24820 34944
rect 24952 34892 25004 34944
rect 25044 34892 25096 34944
rect 29552 34960 29604 35012
rect 31116 34935 31168 34944
rect 31116 34901 31125 34935
rect 31125 34901 31159 34935
rect 31159 34901 31168 34935
rect 31116 34892 31168 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4528 34688 4580 34740
rect 6460 34688 6512 34740
rect 8944 34688 8996 34740
rect 9680 34688 9732 34740
rect 10876 34688 10928 34740
rect 6736 34552 6788 34604
rect 8024 34620 8076 34672
rect 9404 34620 9456 34672
rect 19432 34688 19484 34740
rect 20168 34688 20220 34740
rect 20996 34688 21048 34740
rect 22836 34688 22888 34740
rect 4620 34527 4672 34536
rect 4620 34493 4629 34527
rect 4629 34493 4663 34527
rect 4663 34493 4672 34527
rect 4620 34484 4672 34493
rect 9220 34552 9272 34604
rect 10692 34552 10744 34604
rect 10876 34552 10928 34604
rect 11888 34552 11940 34604
rect 16120 34620 16172 34672
rect 16764 34620 16816 34672
rect 17224 34663 17276 34672
rect 17224 34629 17233 34663
rect 17233 34629 17267 34663
rect 17267 34629 17276 34663
rect 17224 34620 17276 34629
rect 19800 34620 19852 34672
rect 20444 34663 20496 34672
rect 20444 34629 20453 34663
rect 20453 34629 20487 34663
rect 20487 34629 20496 34663
rect 20444 34620 20496 34629
rect 20536 34620 20588 34672
rect 20628 34663 20680 34672
rect 20628 34629 20653 34663
rect 20653 34629 20680 34663
rect 20628 34620 20680 34629
rect 21732 34620 21784 34672
rect 6644 34416 6696 34468
rect 7748 34484 7800 34536
rect 8116 34527 8168 34536
rect 8116 34493 8125 34527
rect 8125 34493 8159 34527
rect 8159 34493 8168 34527
rect 8116 34484 8168 34493
rect 12440 34595 12492 34604
rect 12440 34561 12449 34595
rect 12449 34561 12483 34595
rect 12483 34561 12492 34595
rect 12440 34552 12492 34561
rect 12900 34552 12952 34604
rect 13176 34552 13228 34604
rect 15108 34552 15160 34604
rect 17316 34552 17368 34604
rect 17684 34595 17736 34604
rect 17684 34561 17693 34595
rect 17693 34561 17727 34595
rect 17727 34561 17736 34595
rect 17684 34552 17736 34561
rect 17868 34552 17920 34604
rect 19432 34552 19484 34604
rect 12716 34416 12768 34468
rect 16948 34527 17000 34536
rect 16948 34493 16957 34527
rect 16957 34493 16991 34527
rect 16991 34493 17000 34527
rect 16948 34484 17000 34493
rect 16672 34416 16724 34468
rect 19984 34527 20036 34536
rect 19984 34493 19993 34527
rect 19993 34493 20027 34527
rect 20027 34493 20036 34527
rect 19984 34484 20036 34493
rect 20260 34595 20312 34604
rect 20260 34561 20305 34595
rect 20305 34561 20312 34595
rect 20260 34552 20312 34561
rect 20812 34552 20864 34604
rect 22192 34552 22244 34604
rect 22284 34595 22336 34604
rect 22284 34561 22293 34595
rect 22293 34561 22327 34595
rect 22327 34561 22336 34595
rect 22284 34552 22336 34561
rect 21640 34484 21692 34536
rect 6368 34391 6420 34400
rect 6368 34357 6377 34391
rect 6377 34357 6411 34391
rect 6411 34357 6420 34391
rect 6368 34348 6420 34357
rect 12532 34348 12584 34400
rect 16396 34348 16448 34400
rect 16856 34391 16908 34400
rect 16856 34357 16865 34391
rect 16865 34357 16899 34391
rect 16899 34357 16908 34391
rect 16856 34348 16908 34357
rect 22468 34416 22520 34468
rect 24952 34688 25004 34740
rect 25780 34688 25832 34740
rect 24584 34620 24636 34672
rect 23480 34595 23532 34604
rect 23480 34561 23489 34595
rect 23489 34561 23523 34595
rect 23523 34561 23532 34595
rect 23480 34552 23532 34561
rect 23572 34552 23624 34604
rect 25044 34552 25096 34604
rect 22928 34484 22980 34536
rect 23204 34484 23256 34536
rect 23388 34527 23440 34536
rect 23388 34493 23397 34527
rect 23397 34493 23431 34527
rect 23431 34493 23440 34527
rect 23388 34484 23440 34493
rect 24492 34484 24544 34536
rect 25228 34552 25280 34604
rect 25780 34552 25832 34604
rect 25964 34552 26016 34604
rect 26516 34595 26568 34604
rect 26516 34561 26525 34595
rect 26525 34561 26559 34595
rect 26559 34561 26568 34595
rect 26516 34552 26568 34561
rect 27252 34620 27304 34672
rect 27896 34620 27948 34672
rect 29092 34595 29144 34604
rect 29092 34561 29101 34595
rect 29101 34561 29135 34595
rect 29135 34561 29144 34595
rect 29092 34552 29144 34561
rect 29368 34663 29420 34672
rect 29368 34629 29377 34663
rect 29377 34629 29411 34663
rect 29411 34629 29420 34663
rect 29368 34620 29420 34629
rect 29920 34620 29972 34672
rect 29460 34595 29512 34604
rect 25504 34416 25556 34468
rect 27896 34484 27948 34536
rect 28540 34484 28592 34536
rect 29460 34561 29469 34595
rect 29469 34561 29503 34595
rect 29503 34561 29512 34595
rect 29460 34552 29512 34561
rect 30012 34552 30064 34604
rect 30380 34552 30432 34604
rect 20352 34348 20404 34400
rect 21824 34391 21876 34400
rect 21824 34357 21833 34391
rect 21833 34357 21867 34391
rect 21867 34357 21876 34391
rect 21824 34348 21876 34357
rect 22744 34348 22796 34400
rect 23204 34348 23256 34400
rect 25044 34348 25096 34400
rect 25596 34348 25648 34400
rect 25688 34391 25740 34400
rect 25688 34357 25697 34391
rect 25697 34357 25731 34391
rect 25731 34357 25740 34391
rect 25688 34348 25740 34357
rect 27252 34348 27304 34400
rect 31116 34484 31168 34536
rect 37556 34595 37608 34604
rect 37556 34561 37565 34595
rect 37565 34561 37599 34595
rect 37599 34561 37608 34595
rect 37556 34552 37608 34561
rect 31392 34527 31444 34536
rect 31392 34493 31401 34527
rect 31401 34493 31435 34527
rect 31435 34493 31444 34527
rect 31392 34484 31444 34493
rect 29184 34416 29236 34468
rect 33324 34484 33376 34536
rect 37924 34484 37976 34536
rect 29736 34391 29788 34400
rect 29736 34357 29745 34391
rect 29745 34357 29779 34391
rect 29779 34357 29788 34391
rect 29736 34348 29788 34357
rect 30656 34391 30708 34400
rect 30656 34357 30665 34391
rect 30665 34357 30699 34391
rect 30699 34357 30708 34391
rect 30656 34348 30708 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4620 34144 4672 34196
rect 8116 34144 8168 34196
rect 11980 34144 12032 34196
rect 12808 34144 12860 34196
rect 14648 34144 14700 34196
rect 16856 34144 16908 34196
rect 16948 34144 17000 34196
rect 20168 34144 20220 34196
rect 22468 34144 22520 34196
rect 26516 34144 26568 34196
rect 27436 34144 27488 34196
rect 30380 34144 30432 34196
rect 30656 34144 30708 34196
rect 12348 34119 12400 34128
rect 12348 34085 12357 34119
rect 12357 34085 12391 34119
rect 12391 34085 12400 34119
rect 12348 34076 12400 34085
rect 14280 34076 14332 34128
rect 7748 34008 7800 34060
rect 5448 33940 5500 33992
rect 6368 33940 6420 33992
rect 7104 33983 7156 33992
rect 7104 33949 7113 33983
rect 7113 33949 7147 33983
rect 7147 33949 7156 33983
rect 7104 33940 7156 33949
rect 8208 33872 8260 33924
rect 4528 33847 4580 33856
rect 4528 33813 4537 33847
rect 4537 33813 4571 33847
rect 4571 33813 4580 33847
rect 4528 33804 4580 33813
rect 7196 33847 7248 33856
rect 7196 33813 7205 33847
rect 7205 33813 7239 33847
rect 7239 33813 7248 33847
rect 7196 33804 7248 33813
rect 9956 34051 10008 34060
rect 9956 34017 9965 34051
rect 9965 34017 9999 34051
rect 9999 34017 10008 34051
rect 9956 34008 10008 34017
rect 9680 33983 9732 33992
rect 9680 33949 9689 33983
rect 9689 33949 9723 33983
rect 9723 33949 9732 33983
rect 9680 33940 9732 33949
rect 10232 33940 10284 33992
rect 12532 33940 12584 33992
rect 12624 33983 12676 33992
rect 12624 33949 12633 33983
rect 12633 33949 12667 33983
rect 12667 33949 12676 33983
rect 12624 33940 12676 33949
rect 14740 33983 14792 33992
rect 14740 33949 14749 33983
rect 14749 33949 14783 33983
rect 14783 33949 14792 33983
rect 14740 33940 14792 33949
rect 14924 33983 14976 33992
rect 14924 33949 14933 33983
rect 14933 33949 14967 33983
rect 14967 33949 14976 33983
rect 14924 33940 14976 33949
rect 15752 33940 15804 33992
rect 16028 33940 16080 33992
rect 16120 33940 16172 33992
rect 16488 33983 16540 33992
rect 16488 33949 16497 33983
rect 16497 33949 16531 33983
rect 16531 33949 16540 33983
rect 16488 33940 16540 33949
rect 15936 33872 15988 33924
rect 16672 33940 16724 33992
rect 16948 33940 17000 33992
rect 9772 33847 9824 33856
rect 9772 33813 9781 33847
rect 9781 33813 9815 33847
rect 9815 33813 9824 33847
rect 9772 33804 9824 33813
rect 9864 33804 9916 33856
rect 12532 33847 12584 33856
rect 12532 33813 12541 33847
rect 12541 33813 12575 33847
rect 12575 33813 12584 33847
rect 12532 33804 12584 33813
rect 13084 33804 13136 33856
rect 17132 33847 17184 33856
rect 17132 33813 17141 33847
rect 17141 33813 17175 33847
rect 17175 33813 17184 33847
rect 17132 33804 17184 33813
rect 17224 33804 17276 33856
rect 17316 33804 17368 33856
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18052 33940 18104 33949
rect 17868 33915 17920 33924
rect 17868 33881 17877 33915
rect 17877 33881 17911 33915
rect 17911 33881 17920 33915
rect 17868 33872 17920 33881
rect 17960 33915 18012 33924
rect 17960 33881 17969 33915
rect 17969 33881 18003 33915
rect 18003 33881 18012 33915
rect 17960 33872 18012 33881
rect 18512 33847 18564 33856
rect 18512 33813 18521 33847
rect 18521 33813 18555 33847
rect 18555 33813 18564 33847
rect 18512 33804 18564 33813
rect 19800 33940 19852 33992
rect 20444 33940 20496 33992
rect 21180 34008 21232 34060
rect 24308 34008 24360 34060
rect 24584 34051 24636 34060
rect 24584 34017 24593 34051
rect 24593 34017 24627 34051
rect 24627 34017 24636 34051
rect 24584 34008 24636 34017
rect 19340 33872 19392 33924
rect 20536 33915 20588 33924
rect 20536 33881 20545 33915
rect 20545 33881 20579 33915
rect 20579 33881 20588 33915
rect 20536 33872 20588 33881
rect 21732 33940 21784 33992
rect 22376 33940 22428 33992
rect 25412 33983 25464 33992
rect 25412 33949 25421 33983
rect 25421 33949 25455 33983
rect 25455 33949 25464 33983
rect 25412 33940 25464 33949
rect 27252 34008 27304 34060
rect 27528 34051 27580 34060
rect 27528 34017 27537 34051
rect 27537 34017 27571 34051
rect 27571 34017 27580 34051
rect 27528 34008 27580 34017
rect 28632 34008 28684 34060
rect 29552 34008 29604 34060
rect 25688 33983 25740 33992
rect 25688 33949 25697 33983
rect 25697 33949 25731 33983
rect 25731 33949 25740 33983
rect 25688 33940 25740 33949
rect 26056 33940 26108 33992
rect 24676 33872 24728 33924
rect 27712 33872 27764 33924
rect 29736 33940 29788 33992
rect 30380 33940 30432 33992
rect 31392 34144 31444 34196
rect 32864 34144 32916 34196
rect 33692 34008 33744 34060
rect 32680 33940 32732 33992
rect 32772 33940 32824 33992
rect 30472 33872 30524 33924
rect 33140 33872 33192 33924
rect 34612 33872 34664 33924
rect 21548 33804 21600 33856
rect 21916 33804 21968 33856
rect 22652 33804 22704 33856
rect 25044 33804 25096 33856
rect 25136 33847 25188 33856
rect 25136 33813 25145 33847
rect 25145 33813 25179 33847
rect 25179 33813 25188 33847
rect 25136 33804 25188 33813
rect 26516 33804 26568 33856
rect 27436 33804 27488 33856
rect 28356 33847 28408 33856
rect 28356 33813 28365 33847
rect 28365 33813 28399 33847
rect 28399 33813 28408 33847
rect 28356 33804 28408 33813
rect 28448 33804 28500 33856
rect 31392 33804 31444 33856
rect 33232 33804 33284 33856
rect 33324 33847 33376 33856
rect 33324 33813 33333 33847
rect 33333 33813 33367 33847
rect 33367 33813 33376 33847
rect 33324 33804 33376 33813
rect 34152 33804 34204 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4528 33600 4580 33652
rect 7196 33600 7248 33652
rect 9864 33600 9916 33652
rect 14924 33600 14976 33652
rect 6828 33532 6880 33584
rect 9220 33532 9272 33584
rect 10324 33532 10376 33584
rect 12532 33532 12584 33584
rect 14096 33532 14148 33584
rect 14464 33575 14516 33584
rect 14464 33541 14473 33575
rect 14473 33541 14507 33575
rect 14507 33541 14516 33575
rect 14464 33532 14516 33541
rect 16120 33532 16172 33584
rect 14372 33507 14424 33516
rect 14372 33473 14381 33507
rect 14381 33473 14415 33507
rect 14415 33473 14424 33507
rect 14372 33464 14424 33473
rect 14556 33507 14608 33516
rect 14556 33473 14565 33507
rect 14565 33473 14599 33507
rect 14599 33473 14608 33507
rect 14556 33464 14608 33473
rect 14648 33464 14700 33516
rect 4620 33439 4672 33448
rect 4620 33405 4629 33439
rect 4629 33405 4663 33439
rect 4663 33405 4672 33439
rect 4620 33396 4672 33405
rect 7288 33439 7340 33448
rect 7288 33405 7297 33439
rect 7297 33405 7331 33439
rect 7331 33405 7340 33439
rect 7288 33396 7340 33405
rect 9772 33439 9824 33448
rect 9772 33405 9781 33439
rect 9781 33405 9815 33439
rect 9815 33405 9824 33439
rect 9772 33396 9824 33405
rect 16856 33464 16908 33516
rect 18512 33600 18564 33652
rect 17408 33575 17460 33584
rect 17408 33541 17417 33575
rect 17417 33541 17451 33575
rect 17451 33541 17460 33575
rect 17408 33532 17460 33541
rect 17500 33575 17552 33584
rect 17500 33541 17509 33575
rect 17509 33541 17543 33575
rect 17543 33541 17552 33575
rect 17500 33532 17552 33541
rect 17776 33464 17828 33516
rect 24308 33600 24360 33652
rect 28356 33600 28408 33652
rect 9496 33328 9548 33380
rect 6184 33260 6236 33312
rect 8760 33303 8812 33312
rect 8760 33269 8769 33303
rect 8769 33269 8803 33303
rect 8803 33269 8812 33303
rect 8760 33260 8812 33269
rect 12532 33328 12584 33380
rect 17316 33396 17368 33448
rect 17408 33396 17460 33448
rect 17960 33328 18012 33380
rect 18788 33507 18840 33516
rect 18788 33473 18797 33507
rect 18797 33473 18831 33507
rect 18831 33473 18840 33507
rect 18788 33464 18840 33473
rect 21088 33532 21140 33584
rect 22008 33575 22060 33584
rect 22008 33541 22017 33575
rect 22017 33541 22051 33575
rect 22051 33541 22060 33575
rect 22008 33532 22060 33541
rect 22100 33575 22152 33584
rect 22100 33541 22109 33575
rect 22109 33541 22143 33575
rect 22143 33541 22152 33575
rect 22100 33532 22152 33541
rect 22744 33532 22796 33584
rect 23296 33532 23348 33584
rect 18880 33396 18932 33448
rect 19432 33396 19484 33448
rect 19892 33464 19944 33516
rect 20536 33464 20588 33516
rect 21456 33464 21508 33516
rect 23756 33464 23808 33516
rect 24952 33532 25004 33584
rect 19616 33439 19668 33448
rect 19616 33405 19625 33439
rect 19625 33405 19659 33439
rect 19659 33405 19668 33439
rect 19616 33396 19668 33405
rect 21732 33328 21784 33380
rect 23388 33396 23440 33448
rect 25688 33464 25740 33516
rect 28540 33532 28592 33584
rect 33324 33600 33376 33652
rect 37556 33600 37608 33652
rect 31668 33532 31720 33584
rect 33600 33532 33652 33584
rect 32864 33507 32916 33516
rect 32864 33473 32873 33507
rect 32873 33473 32907 33507
rect 32907 33473 32916 33507
rect 32864 33464 32916 33473
rect 34152 33464 34204 33516
rect 37556 33507 37608 33516
rect 37556 33473 37565 33507
rect 37565 33473 37599 33507
rect 37599 33473 37608 33507
rect 37556 33464 37608 33473
rect 26240 33396 26292 33448
rect 28448 33439 28500 33448
rect 28448 33405 28457 33439
rect 28457 33405 28491 33439
rect 28491 33405 28500 33439
rect 28448 33396 28500 33405
rect 11060 33260 11112 33312
rect 15936 33260 15988 33312
rect 18328 33260 18380 33312
rect 21364 33260 21416 33312
rect 22836 33260 22888 33312
rect 29736 33260 29788 33312
rect 30196 33260 30248 33312
rect 33324 33260 33376 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4620 33056 4672 33108
rect 7288 33056 7340 33108
rect 8116 33056 8168 33108
rect 6644 32920 6696 32972
rect 8116 32920 8168 32972
rect 9772 33099 9824 33108
rect 9772 33065 9781 33099
rect 9781 33065 9815 33099
rect 9815 33065 9824 33099
rect 9772 33056 9824 33065
rect 10048 33056 10100 33108
rect 10508 33056 10560 33108
rect 17132 33056 17184 33108
rect 17408 33056 17460 33108
rect 17684 33056 17736 33108
rect 18328 33099 18380 33108
rect 18328 33065 18337 33099
rect 18337 33065 18371 33099
rect 18371 33065 18380 33099
rect 18328 33056 18380 33065
rect 20168 33056 20220 33108
rect 6184 32759 6236 32768
rect 6184 32725 6193 32759
rect 6193 32725 6227 32759
rect 6227 32725 6236 32759
rect 6184 32716 6236 32725
rect 8760 32852 8812 32904
rect 8944 32852 8996 32904
rect 9496 32852 9548 32904
rect 9956 32895 10008 32904
rect 9956 32861 9965 32895
rect 9965 32861 9999 32895
rect 9999 32861 10008 32895
rect 9956 32852 10008 32861
rect 10048 32895 10100 32904
rect 10048 32861 10057 32895
rect 10057 32861 10091 32895
rect 10091 32861 10100 32895
rect 10048 32852 10100 32861
rect 8852 32784 8904 32836
rect 9404 32716 9456 32768
rect 10692 32784 10744 32836
rect 13084 32852 13136 32904
rect 15660 32920 15712 32972
rect 16304 32920 16356 32972
rect 17868 32920 17920 32972
rect 17960 32852 18012 32904
rect 18880 32920 18932 32972
rect 18972 32920 19024 32972
rect 18236 32852 18288 32904
rect 20444 32988 20496 33040
rect 22284 33056 22336 33108
rect 23848 33056 23900 33108
rect 28448 33056 28500 33108
rect 37556 33056 37608 33108
rect 21916 32988 21968 33040
rect 22744 32988 22796 33040
rect 20628 32852 20680 32904
rect 20996 32852 21048 32904
rect 13452 32784 13504 32836
rect 14464 32784 14516 32836
rect 16304 32784 16356 32836
rect 17224 32784 17276 32836
rect 12716 32716 12768 32768
rect 12808 32716 12860 32768
rect 16948 32759 17000 32768
rect 16948 32725 16957 32759
rect 16957 32725 16991 32759
rect 16991 32725 17000 32759
rect 16948 32716 17000 32725
rect 17592 32716 17644 32768
rect 17960 32716 18012 32768
rect 18696 32784 18748 32836
rect 19432 32827 19484 32836
rect 19432 32793 19441 32827
rect 19441 32793 19475 32827
rect 19475 32793 19484 32827
rect 19432 32784 19484 32793
rect 19892 32716 19944 32768
rect 20076 32716 20128 32768
rect 20628 32716 20680 32768
rect 21180 32716 21232 32768
rect 22008 32852 22060 32904
rect 22192 32895 22244 32904
rect 22192 32861 22201 32895
rect 22201 32861 22235 32895
rect 22235 32861 22244 32895
rect 22192 32852 22244 32861
rect 22652 32895 22704 32904
rect 22652 32861 22666 32895
rect 22666 32861 22700 32895
rect 22700 32861 22704 32895
rect 22652 32852 22704 32861
rect 22836 32852 22888 32904
rect 23020 32895 23072 32904
rect 23020 32861 23030 32895
rect 23030 32861 23064 32895
rect 23064 32861 23072 32895
rect 23020 32852 23072 32861
rect 21456 32759 21508 32768
rect 21456 32725 21465 32759
rect 21465 32725 21499 32759
rect 21499 32725 21508 32759
rect 21456 32716 21508 32725
rect 21824 32759 21876 32768
rect 21824 32725 21833 32759
rect 21833 32725 21867 32759
rect 21867 32725 21876 32759
rect 21824 32716 21876 32725
rect 22376 32784 22428 32836
rect 22744 32716 22796 32768
rect 23112 32716 23164 32768
rect 23296 32827 23348 32836
rect 23296 32793 23305 32827
rect 23305 32793 23339 32827
rect 23339 32793 23348 32827
rect 23296 32784 23348 32793
rect 23848 32852 23900 32904
rect 25412 32852 25464 32904
rect 25780 32895 25832 32904
rect 25780 32861 25789 32895
rect 25789 32861 25823 32895
rect 25823 32861 25832 32895
rect 25780 32852 25832 32861
rect 26056 32895 26108 32904
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 26148 32895 26200 32904
rect 26148 32861 26157 32895
rect 26157 32861 26191 32895
rect 26191 32861 26200 32895
rect 26148 32852 26200 32861
rect 24032 32784 24084 32836
rect 24308 32784 24360 32836
rect 26332 32852 26384 32904
rect 27068 32895 27120 32904
rect 27068 32861 27077 32895
rect 27077 32861 27111 32895
rect 27111 32861 27120 32895
rect 27068 32852 27120 32861
rect 31484 32988 31536 33040
rect 28632 32920 28684 32972
rect 28908 32920 28960 32972
rect 23480 32716 23532 32768
rect 25596 32759 25648 32768
rect 25596 32725 25605 32759
rect 25605 32725 25639 32759
rect 25639 32725 25648 32759
rect 25596 32716 25648 32725
rect 26424 32759 26476 32768
rect 26424 32725 26433 32759
rect 26433 32725 26467 32759
rect 26467 32725 26476 32759
rect 26424 32716 26476 32725
rect 27160 32759 27212 32768
rect 27160 32725 27169 32759
rect 27169 32725 27203 32759
rect 27203 32725 27212 32759
rect 27160 32716 27212 32725
rect 27896 32784 27948 32836
rect 29000 32852 29052 32904
rect 33416 32963 33468 32972
rect 33416 32929 33425 32963
rect 33425 32929 33459 32963
rect 33459 32929 33468 32963
rect 33416 32920 33468 32929
rect 33232 32895 33284 32904
rect 28448 32784 28500 32836
rect 33232 32861 33241 32895
rect 33241 32861 33275 32895
rect 33275 32861 33284 32895
rect 33232 32852 33284 32861
rect 30748 32784 30800 32836
rect 33968 32784 34020 32836
rect 34612 32784 34664 32836
rect 34796 32852 34848 32904
rect 29736 32716 29788 32768
rect 33692 32759 33744 32768
rect 33692 32725 33701 32759
rect 33701 32725 33735 32759
rect 33735 32725 33744 32759
rect 33692 32716 33744 32725
rect 34796 32759 34848 32768
rect 34796 32725 34805 32759
rect 34805 32725 34839 32759
rect 34839 32725 34848 32759
rect 34796 32716 34848 32725
rect 35072 32759 35124 32768
rect 35072 32725 35081 32759
rect 35081 32725 35115 32759
rect 35115 32725 35124 32759
rect 35072 32716 35124 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 8760 32512 8812 32564
rect 12348 32512 12400 32564
rect 6184 32444 6236 32496
rect 5356 32376 5408 32428
rect 10048 32444 10100 32496
rect 11060 32444 11112 32496
rect 10692 32376 10744 32428
rect 11520 32376 11572 32428
rect 6736 32308 6788 32360
rect 11980 32376 12032 32428
rect 12348 32419 12400 32428
rect 12348 32385 12358 32419
rect 12358 32385 12392 32419
rect 12392 32385 12400 32419
rect 12348 32376 12400 32385
rect 12440 32308 12492 32360
rect 12900 32376 12952 32428
rect 15200 32376 15252 32428
rect 18236 32376 18288 32428
rect 18328 32376 18380 32428
rect 20720 32444 20772 32496
rect 21824 32512 21876 32564
rect 22192 32512 22244 32564
rect 22376 32512 22428 32564
rect 22652 32512 22704 32564
rect 23020 32512 23072 32564
rect 18696 32419 18748 32428
rect 18696 32385 18705 32419
rect 18705 32385 18739 32419
rect 18739 32385 18748 32419
rect 18696 32376 18748 32385
rect 18880 32376 18932 32428
rect 19156 32376 19208 32428
rect 19524 32376 19576 32428
rect 20076 32419 20128 32428
rect 20076 32385 20085 32419
rect 20085 32385 20119 32419
rect 20119 32385 20128 32419
rect 20076 32376 20128 32385
rect 12624 32240 12676 32292
rect 14464 32308 14516 32360
rect 20168 32308 20220 32360
rect 22008 32419 22060 32428
rect 22008 32385 22015 32419
rect 22015 32385 22060 32419
rect 22008 32376 22060 32385
rect 22100 32419 22152 32428
rect 22100 32385 22109 32419
rect 22109 32385 22143 32419
rect 22143 32385 22152 32419
rect 22100 32376 22152 32385
rect 20720 32240 20772 32292
rect 21732 32308 21784 32360
rect 23112 32444 23164 32496
rect 23388 32444 23440 32496
rect 23480 32444 23532 32496
rect 25596 32512 25648 32564
rect 26332 32512 26384 32564
rect 26424 32512 26476 32564
rect 22744 32376 22796 32428
rect 22928 32376 22980 32428
rect 22652 32308 22704 32360
rect 7472 32172 7524 32224
rect 10692 32215 10744 32224
rect 10692 32181 10701 32215
rect 10701 32181 10735 32215
rect 10735 32181 10744 32215
rect 10692 32172 10744 32181
rect 12900 32215 12952 32224
rect 12900 32181 12909 32215
rect 12909 32181 12943 32215
rect 12943 32181 12952 32215
rect 12900 32172 12952 32181
rect 13176 32172 13228 32224
rect 18236 32215 18288 32224
rect 18236 32181 18245 32215
rect 18245 32181 18279 32215
rect 18279 32181 18288 32215
rect 18236 32172 18288 32181
rect 19892 32172 19944 32224
rect 20168 32172 20220 32224
rect 22284 32240 22336 32292
rect 23020 32308 23072 32360
rect 23388 32351 23440 32360
rect 23388 32317 23397 32351
rect 23397 32317 23431 32351
rect 23431 32317 23440 32351
rect 23388 32308 23440 32317
rect 23848 32419 23900 32428
rect 23848 32385 23857 32419
rect 23857 32385 23891 32419
rect 23891 32385 23900 32419
rect 23848 32376 23900 32385
rect 23756 32308 23808 32360
rect 24124 32376 24176 32428
rect 24584 32376 24636 32428
rect 24952 32376 25004 32428
rect 25320 32376 25372 32428
rect 25688 32419 25740 32428
rect 25688 32385 25697 32419
rect 25697 32385 25731 32419
rect 25731 32385 25740 32419
rect 25688 32376 25740 32385
rect 26240 32444 26292 32496
rect 25044 32308 25096 32360
rect 25504 32308 25556 32360
rect 23940 32240 23992 32292
rect 24860 32240 24912 32292
rect 26148 32240 26200 32292
rect 21732 32172 21784 32224
rect 23480 32172 23532 32224
rect 23572 32172 23624 32224
rect 23848 32172 23900 32224
rect 26240 32172 26292 32224
rect 26516 32351 26568 32360
rect 26516 32317 26525 32351
rect 26525 32317 26559 32351
rect 26559 32317 26568 32351
rect 26516 32308 26568 32317
rect 26608 32351 26660 32360
rect 26608 32317 26617 32351
rect 26617 32317 26651 32351
rect 26651 32317 26660 32351
rect 26608 32308 26660 32317
rect 27160 32512 27212 32564
rect 29092 32512 29144 32564
rect 29644 32512 29696 32564
rect 28540 32444 28592 32496
rect 28632 32444 28684 32496
rect 30196 32444 30248 32496
rect 29644 32419 29696 32428
rect 29644 32385 29653 32419
rect 29653 32385 29687 32419
rect 29687 32385 29696 32419
rect 29644 32376 29696 32385
rect 29736 32419 29788 32428
rect 29736 32385 29746 32419
rect 29746 32385 29780 32419
rect 29780 32385 29788 32419
rect 29736 32376 29788 32385
rect 29000 32351 29052 32360
rect 29000 32317 29009 32351
rect 29009 32317 29043 32351
rect 29043 32317 29052 32351
rect 29000 32308 29052 32317
rect 30104 32419 30156 32428
rect 30104 32385 30118 32419
rect 30118 32385 30152 32419
rect 30152 32385 30156 32419
rect 30380 32512 30432 32564
rect 30748 32555 30800 32564
rect 30748 32521 30757 32555
rect 30757 32521 30791 32555
rect 30791 32521 30800 32555
rect 30748 32512 30800 32521
rect 30104 32376 30156 32385
rect 30840 32419 30892 32428
rect 30840 32385 30849 32419
rect 30849 32385 30883 32419
rect 30883 32385 30892 32419
rect 30840 32376 30892 32385
rect 30012 32308 30064 32360
rect 32496 32512 32548 32564
rect 31484 32444 31536 32496
rect 34796 32512 34848 32564
rect 35072 32512 35124 32564
rect 33232 32444 33284 32496
rect 30564 32240 30616 32292
rect 33968 32376 34020 32428
rect 31484 32172 31536 32224
rect 32128 32215 32180 32224
rect 32128 32181 32137 32215
rect 32137 32181 32171 32215
rect 32171 32181 32180 32215
rect 32128 32172 32180 32181
rect 33692 32308 33744 32360
rect 34244 32308 34296 32360
rect 36636 32351 36688 32360
rect 36636 32317 36645 32351
rect 36645 32317 36679 32351
rect 36679 32317 36688 32351
rect 36636 32308 36688 32317
rect 33968 32172 34020 32224
rect 34152 32172 34204 32224
rect 35900 32172 35952 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3884 31807 3936 31816
rect 3884 31773 3893 31807
rect 3893 31773 3927 31807
rect 3927 31773 3936 31807
rect 3884 31764 3936 31773
rect 6828 31968 6880 32020
rect 7840 31968 7892 32020
rect 8208 31968 8260 32020
rect 8024 31900 8076 31952
rect 9404 31900 9456 31952
rect 4160 31739 4212 31748
rect 4160 31705 4169 31739
rect 4169 31705 4203 31739
rect 4203 31705 4212 31739
rect 4160 31696 4212 31705
rect 5816 31807 5868 31816
rect 5816 31773 5825 31807
rect 5825 31773 5859 31807
rect 5859 31773 5868 31807
rect 5816 31764 5868 31773
rect 8944 31832 8996 31884
rect 11152 31968 11204 32020
rect 11704 31968 11756 32020
rect 12716 31968 12768 32020
rect 18604 32011 18656 32020
rect 18604 31977 18613 32011
rect 18613 31977 18647 32011
rect 18647 31977 18656 32011
rect 18604 31968 18656 31977
rect 20352 31968 20404 32020
rect 10232 31832 10284 31884
rect 12808 31764 12860 31816
rect 12900 31764 12952 31816
rect 10600 31739 10652 31748
rect 10600 31705 10609 31739
rect 10609 31705 10643 31739
rect 10643 31705 10652 31739
rect 10600 31696 10652 31705
rect 10876 31696 10928 31748
rect 14740 31832 14792 31884
rect 20628 31900 20680 31952
rect 20720 31900 20772 31952
rect 20904 31900 20956 31952
rect 21456 31900 21508 31952
rect 16856 31764 16908 31816
rect 17132 31764 17184 31816
rect 14280 31696 14332 31748
rect 14464 31696 14516 31748
rect 6736 31628 6788 31680
rect 7748 31671 7800 31680
rect 7748 31637 7757 31671
rect 7757 31637 7791 31671
rect 7791 31637 7800 31671
rect 7748 31628 7800 31637
rect 8668 31671 8720 31680
rect 8668 31637 8677 31671
rect 8677 31637 8711 31671
rect 8711 31637 8720 31671
rect 8668 31628 8720 31637
rect 9404 31628 9456 31680
rect 12072 31671 12124 31680
rect 12072 31637 12081 31671
rect 12081 31637 12115 31671
rect 12115 31637 12124 31671
rect 12072 31628 12124 31637
rect 14372 31628 14424 31680
rect 14648 31671 14700 31680
rect 14648 31637 14657 31671
rect 14657 31637 14691 31671
rect 14691 31637 14700 31671
rect 14648 31628 14700 31637
rect 14924 31671 14976 31680
rect 14924 31637 14933 31671
rect 14933 31637 14967 31671
rect 14967 31637 14976 31671
rect 14924 31628 14976 31637
rect 15476 31696 15528 31748
rect 16304 31696 16356 31748
rect 19064 31764 19116 31816
rect 19984 31764 20036 31816
rect 20352 31832 20404 31884
rect 20536 31832 20588 31884
rect 20812 31875 20864 31884
rect 20812 31841 20821 31875
rect 20821 31841 20855 31875
rect 20855 31841 20864 31875
rect 20812 31832 20864 31841
rect 21180 31832 21232 31884
rect 22560 31968 22612 32020
rect 23756 31968 23808 32020
rect 26056 31968 26108 32020
rect 26240 31968 26292 32020
rect 27160 31968 27212 32020
rect 27988 31968 28040 32020
rect 28356 31968 28408 32020
rect 30748 31968 30800 32020
rect 32128 31968 32180 32020
rect 32496 31968 32548 32020
rect 33600 31968 33652 32020
rect 34152 31968 34204 32020
rect 34244 32011 34296 32020
rect 34244 31977 34253 32011
rect 34253 31977 34287 32011
rect 34287 31977 34296 32011
rect 34244 31968 34296 31977
rect 22008 31832 22060 31884
rect 18972 31696 19024 31748
rect 18788 31628 18840 31680
rect 19800 31628 19852 31680
rect 20352 31628 20404 31680
rect 20996 31696 21048 31748
rect 21180 31628 21232 31680
rect 21272 31628 21324 31680
rect 21640 31628 21692 31680
rect 22192 31764 22244 31816
rect 22560 31764 22612 31816
rect 22744 31807 22796 31816
rect 22744 31773 22753 31807
rect 22753 31773 22787 31807
rect 22787 31773 22796 31807
rect 22744 31764 22796 31773
rect 30564 31900 30616 31952
rect 24952 31832 25004 31884
rect 23388 31764 23440 31816
rect 24584 31764 24636 31816
rect 22468 31628 22520 31680
rect 23020 31628 23072 31680
rect 23112 31628 23164 31680
rect 25228 31696 25280 31748
rect 25504 31696 25556 31748
rect 25872 31764 25924 31816
rect 26056 31764 26108 31816
rect 29000 31832 29052 31884
rect 31116 31875 31168 31884
rect 31116 31841 31125 31875
rect 31125 31841 31159 31875
rect 31159 31841 31168 31875
rect 31116 31832 31168 31841
rect 31852 31832 31904 31884
rect 33600 31832 33652 31884
rect 33968 31875 34020 31884
rect 33968 31841 33977 31875
rect 33977 31841 34011 31875
rect 34011 31841 34020 31875
rect 33968 31832 34020 31841
rect 30196 31807 30248 31816
rect 30196 31773 30205 31807
rect 30205 31773 30239 31807
rect 30239 31773 30248 31807
rect 30196 31764 30248 31773
rect 30380 31807 30432 31816
rect 30380 31773 30389 31807
rect 30389 31773 30423 31807
rect 30423 31773 30432 31807
rect 30380 31764 30432 31773
rect 30472 31764 30524 31816
rect 28632 31696 28684 31748
rect 29000 31628 29052 31680
rect 31760 31696 31812 31748
rect 36636 31628 36688 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 3884 31424 3936 31476
rect 4160 31424 4212 31476
rect 5816 31424 5868 31476
rect 6736 31467 6788 31476
rect 6736 31433 6745 31467
rect 6745 31433 6779 31467
rect 6779 31433 6788 31467
rect 6736 31424 6788 31433
rect 8116 31424 8168 31476
rect 11520 31467 11572 31476
rect 11520 31433 11529 31467
rect 11529 31433 11563 31467
rect 11563 31433 11572 31467
rect 11520 31424 11572 31433
rect 14280 31467 14332 31476
rect 14280 31433 14289 31467
rect 14289 31433 14323 31467
rect 14323 31433 14332 31467
rect 14280 31424 14332 31433
rect 7748 31399 7800 31408
rect 7748 31365 7757 31399
rect 7757 31365 7791 31399
rect 7791 31365 7800 31399
rect 7748 31356 7800 31365
rect 7840 31356 7892 31408
rect 16580 31356 16632 31408
rect 16948 31356 17000 31408
rect 5356 31288 5408 31340
rect 5540 31288 5592 31340
rect 6644 31288 6696 31340
rect 7472 31331 7524 31340
rect 7472 31297 7481 31331
rect 7481 31297 7515 31331
rect 7515 31297 7524 31331
rect 7472 31288 7524 31297
rect 6460 31220 6512 31272
rect 6828 31220 6880 31272
rect 9404 31263 9456 31272
rect 9404 31229 9413 31263
rect 9413 31229 9447 31263
rect 9447 31229 9456 31263
rect 9404 31220 9456 31229
rect 9680 31263 9732 31272
rect 9680 31229 9689 31263
rect 9689 31229 9723 31263
rect 9723 31229 9732 31263
rect 9680 31220 9732 31229
rect 10876 31220 10928 31272
rect 13728 31288 13780 31340
rect 15292 31288 15344 31340
rect 12072 31220 12124 31272
rect 12164 31263 12216 31272
rect 12164 31229 12173 31263
rect 12173 31229 12207 31263
rect 12207 31229 12216 31263
rect 12164 31220 12216 31229
rect 16580 31220 16632 31272
rect 16948 31220 17000 31272
rect 17592 31356 17644 31408
rect 18880 31356 18932 31408
rect 17500 31331 17552 31340
rect 17500 31297 17509 31331
rect 17509 31297 17543 31331
rect 17543 31297 17552 31331
rect 17500 31288 17552 31297
rect 18604 31331 18656 31340
rect 18604 31297 18613 31331
rect 18613 31297 18647 31331
rect 18647 31297 18656 31331
rect 18604 31288 18656 31297
rect 18696 31288 18748 31340
rect 19156 31331 19208 31340
rect 19156 31297 19165 31331
rect 19165 31297 19199 31331
rect 19199 31297 19208 31331
rect 19156 31288 19208 31297
rect 20536 31356 20588 31408
rect 20812 31424 20864 31476
rect 22008 31424 22060 31476
rect 22100 31356 22152 31408
rect 19892 31288 19944 31340
rect 20720 31288 20772 31340
rect 20904 31288 20956 31340
rect 21548 31288 21600 31340
rect 22928 31424 22980 31476
rect 23296 31424 23348 31476
rect 24216 31424 24268 31476
rect 28816 31424 28868 31476
rect 29000 31424 29052 31476
rect 22928 31331 22980 31340
rect 22928 31297 22937 31331
rect 22937 31297 22971 31331
rect 22971 31297 22980 31331
rect 22928 31288 22980 31297
rect 23020 31331 23072 31340
rect 23020 31297 23029 31331
rect 23029 31297 23063 31331
rect 23063 31297 23072 31331
rect 23020 31288 23072 31297
rect 23296 31288 23348 31340
rect 25688 31356 25740 31408
rect 25872 31356 25924 31408
rect 28632 31356 28684 31408
rect 30196 31424 30248 31476
rect 31300 31424 31352 31476
rect 31852 31424 31904 31476
rect 18144 31220 18196 31272
rect 20260 31220 20312 31272
rect 20628 31220 20680 31272
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 26148 31288 26200 31340
rect 27896 31331 27948 31340
rect 27896 31297 27905 31331
rect 27905 31297 27939 31331
rect 27939 31297 27948 31331
rect 27896 31288 27948 31297
rect 27988 31331 28040 31340
rect 27988 31297 27997 31331
rect 27997 31297 28031 31331
rect 28031 31297 28040 31331
rect 27988 31288 28040 31297
rect 28080 31331 28132 31340
rect 28080 31297 28089 31331
rect 28089 31297 28123 31331
rect 28123 31297 28132 31331
rect 28080 31288 28132 31297
rect 28264 31331 28316 31340
rect 28264 31297 28273 31331
rect 28273 31297 28307 31331
rect 28307 31297 28316 31331
rect 28264 31288 28316 31297
rect 28816 31288 28868 31340
rect 29000 31331 29052 31340
rect 29000 31297 29009 31331
rect 29009 31297 29043 31331
rect 29043 31297 29052 31331
rect 29000 31288 29052 31297
rect 29092 31331 29144 31340
rect 29092 31297 29101 31331
rect 29101 31297 29135 31331
rect 29135 31297 29144 31331
rect 29092 31288 29144 31297
rect 29276 31331 29328 31340
rect 29276 31297 29285 31331
rect 29285 31297 29319 31331
rect 29319 31297 29328 31331
rect 29276 31288 29328 31297
rect 23848 31220 23900 31272
rect 27068 31220 27120 31272
rect 29920 31288 29972 31340
rect 30564 31288 30616 31340
rect 31300 31331 31352 31340
rect 31300 31297 31309 31331
rect 31309 31297 31343 31331
rect 31343 31297 31352 31331
rect 31300 31288 31352 31297
rect 31576 31331 31628 31340
rect 31576 31297 31585 31331
rect 31585 31297 31619 31331
rect 31619 31297 31628 31331
rect 31576 31288 31628 31297
rect 32312 31331 32364 31340
rect 32312 31297 32321 31331
rect 32321 31297 32355 31331
rect 32355 31297 32364 31331
rect 32312 31288 32364 31297
rect 34612 31288 34664 31340
rect 9220 31127 9272 31136
rect 9220 31093 9229 31127
rect 9229 31093 9263 31127
rect 9263 31093 9272 31127
rect 9220 31084 9272 31093
rect 11060 31084 11112 31136
rect 11244 31084 11296 31136
rect 11520 31084 11572 31136
rect 13268 31084 13320 31136
rect 16212 31084 16264 31136
rect 17040 31127 17092 31136
rect 17040 31093 17049 31127
rect 17049 31093 17083 31127
rect 17083 31093 17092 31127
rect 17040 31084 17092 31093
rect 17408 31152 17460 31204
rect 17684 31127 17736 31136
rect 17684 31093 17693 31127
rect 17693 31093 17727 31127
rect 17727 31093 17736 31127
rect 17684 31084 17736 31093
rect 17960 31152 18012 31204
rect 18236 31084 18288 31136
rect 18420 31084 18472 31136
rect 19340 31084 19392 31136
rect 20628 31084 20680 31136
rect 20996 31084 21048 31136
rect 21456 31084 21508 31136
rect 22928 31084 22980 31136
rect 23204 31127 23256 31136
rect 23204 31093 23213 31127
rect 23213 31093 23247 31127
rect 23247 31093 23256 31127
rect 23204 31084 23256 31093
rect 24032 31084 24084 31136
rect 25228 31127 25280 31136
rect 25228 31093 25237 31127
rect 25237 31093 25271 31127
rect 25271 31093 25280 31127
rect 25228 31084 25280 31093
rect 25596 31127 25648 31136
rect 25596 31093 25605 31127
rect 25605 31093 25639 31127
rect 25639 31093 25648 31127
rect 25596 31084 25648 31093
rect 27712 31084 27764 31136
rect 28080 31084 28132 31136
rect 28816 31084 28868 31136
rect 29276 31084 29328 31136
rect 30472 31084 30524 31136
rect 32036 31084 32088 31136
rect 32404 31084 32456 31136
rect 34796 31084 34848 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 8024 30923 8076 30932
rect 8024 30889 8033 30923
rect 8033 30889 8067 30923
rect 8067 30889 8076 30923
rect 8024 30880 8076 30889
rect 8944 30923 8996 30932
rect 8944 30889 8953 30923
rect 8953 30889 8987 30923
rect 8987 30889 8996 30923
rect 8944 30880 8996 30889
rect 9680 30880 9732 30932
rect 12072 30880 12124 30932
rect 6828 30744 6880 30796
rect 6368 30540 6420 30592
rect 6644 30540 6696 30592
rect 7932 30608 7984 30660
rect 8208 30719 8260 30728
rect 8208 30685 8217 30719
rect 8217 30685 8251 30719
rect 8251 30685 8260 30719
rect 8208 30676 8260 30685
rect 8484 30608 8536 30660
rect 8668 30676 8720 30728
rect 8944 30676 8996 30728
rect 9220 30676 9272 30728
rect 10692 30744 10744 30796
rect 11244 30608 11296 30660
rect 12624 30719 12676 30728
rect 12624 30685 12633 30719
rect 12633 30685 12667 30719
rect 12667 30685 12676 30719
rect 12624 30676 12676 30685
rect 15476 30880 15528 30932
rect 16764 30880 16816 30932
rect 16948 30880 17000 30932
rect 19892 30880 19944 30932
rect 14832 30812 14884 30864
rect 13084 30676 13136 30728
rect 14924 30787 14976 30796
rect 14924 30753 14933 30787
rect 14933 30753 14967 30787
rect 14967 30753 14976 30787
rect 14924 30744 14976 30753
rect 16580 30787 16632 30796
rect 15016 30719 15068 30728
rect 15016 30685 15025 30719
rect 15025 30685 15059 30719
rect 15059 30685 15068 30719
rect 15016 30676 15068 30685
rect 15108 30676 15160 30728
rect 8760 30583 8812 30592
rect 8760 30549 8769 30583
rect 8769 30549 8803 30583
rect 8803 30549 8812 30583
rect 8760 30540 8812 30549
rect 9220 30540 9272 30592
rect 11060 30583 11112 30592
rect 11060 30549 11069 30583
rect 11069 30549 11103 30583
rect 11103 30549 11112 30583
rect 11060 30540 11112 30549
rect 13636 30540 13688 30592
rect 14556 30583 14608 30592
rect 14556 30549 14565 30583
rect 14565 30549 14599 30583
rect 14599 30549 14608 30583
rect 14556 30540 14608 30549
rect 14924 30540 14976 30592
rect 16580 30753 16589 30787
rect 16589 30753 16623 30787
rect 16623 30753 16632 30787
rect 16580 30744 16632 30753
rect 15660 30676 15712 30728
rect 16028 30676 16080 30728
rect 17040 30812 17092 30864
rect 17224 30812 17276 30864
rect 17592 30812 17644 30864
rect 17868 30812 17920 30864
rect 18972 30812 19024 30864
rect 20812 30812 20864 30864
rect 15476 30540 15528 30592
rect 16580 30540 16632 30592
rect 17224 30676 17276 30728
rect 16948 30651 17000 30660
rect 16948 30617 16957 30651
rect 16957 30617 16991 30651
rect 16991 30617 17000 30651
rect 16948 30608 17000 30617
rect 17316 30583 17368 30592
rect 17316 30549 17325 30583
rect 17325 30549 17359 30583
rect 17359 30549 17368 30583
rect 17316 30540 17368 30549
rect 18144 30676 18196 30728
rect 18696 30676 18748 30728
rect 18328 30608 18380 30660
rect 18512 30651 18564 30660
rect 18512 30617 18521 30651
rect 18521 30617 18555 30651
rect 18555 30617 18564 30651
rect 18512 30608 18564 30617
rect 19340 30719 19392 30728
rect 19340 30685 19349 30719
rect 19349 30685 19383 30719
rect 19383 30685 19392 30719
rect 19340 30676 19392 30685
rect 21180 30812 21232 30864
rect 21456 30812 21508 30864
rect 21732 30744 21784 30796
rect 23204 30880 23256 30932
rect 23480 30880 23532 30932
rect 23940 30880 23992 30932
rect 27988 30880 28040 30932
rect 29000 30880 29052 30932
rect 30196 30880 30248 30932
rect 34796 30880 34848 30932
rect 25596 30812 25648 30864
rect 29276 30812 29328 30864
rect 21272 30719 21324 30728
rect 21272 30685 21281 30719
rect 21281 30685 21315 30719
rect 21315 30685 21324 30719
rect 21272 30676 21324 30685
rect 21364 30719 21416 30728
rect 21364 30685 21373 30719
rect 21373 30685 21407 30719
rect 21407 30685 21416 30719
rect 21364 30676 21416 30685
rect 21456 30676 21508 30728
rect 21824 30676 21876 30728
rect 22376 30676 22428 30728
rect 22836 30676 22888 30728
rect 23664 30676 23716 30728
rect 23756 30719 23808 30728
rect 23756 30685 23765 30719
rect 23765 30685 23799 30719
rect 23799 30685 23808 30719
rect 23756 30676 23808 30685
rect 23940 30719 23992 30728
rect 23940 30685 23949 30719
rect 23949 30685 23983 30719
rect 23983 30685 23992 30719
rect 23940 30676 23992 30685
rect 18052 30540 18104 30592
rect 19340 30540 19392 30592
rect 22376 30540 22428 30592
rect 22928 30583 22980 30592
rect 22928 30549 22937 30583
rect 22937 30549 22971 30583
rect 22971 30549 22980 30583
rect 22928 30540 22980 30549
rect 23296 30583 23348 30592
rect 23296 30549 23305 30583
rect 23305 30549 23339 30583
rect 23339 30549 23348 30583
rect 23296 30540 23348 30549
rect 25320 30676 25372 30728
rect 25872 30787 25924 30796
rect 25872 30753 25881 30787
rect 25881 30753 25915 30787
rect 25915 30753 25924 30787
rect 25872 30744 25924 30753
rect 25596 30719 25648 30728
rect 25596 30685 25605 30719
rect 25605 30685 25639 30719
rect 25639 30685 25648 30719
rect 25596 30676 25648 30685
rect 27068 30719 27120 30728
rect 27068 30685 27077 30719
rect 27077 30685 27111 30719
rect 27111 30685 27120 30719
rect 27068 30676 27120 30685
rect 28816 30719 28868 30728
rect 28816 30685 28825 30719
rect 28825 30685 28859 30719
rect 28859 30685 28868 30719
rect 28816 30676 28868 30685
rect 29184 30719 29236 30728
rect 29184 30685 29193 30719
rect 29193 30685 29227 30719
rect 29227 30685 29236 30719
rect 29184 30676 29236 30685
rect 29000 30608 29052 30660
rect 34336 30719 34388 30728
rect 34336 30685 34345 30719
rect 34345 30685 34379 30719
rect 34379 30685 34388 30719
rect 34336 30676 34388 30685
rect 23664 30540 23716 30592
rect 26976 30540 27028 30592
rect 29092 30540 29144 30592
rect 32220 30583 32272 30592
rect 32220 30549 32229 30583
rect 32229 30549 32263 30583
rect 32263 30549 32272 30583
rect 32220 30540 32272 30549
rect 32496 30540 32548 30592
rect 33048 30540 33100 30592
rect 35992 30608 36044 30660
rect 34520 30540 34572 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 8024 30200 8076 30252
rect 8760 30336 8812 30388
rect 9312 30336 9364 30388
rect 8484 30311 8536 30320
rect 8484 30277 8493 30311
rect 8493 30277 8527 30311
rect 8527 30277 8536 30311
rect 8484 30268 8536 30277
rect 10968 30268 11020 30320
rect 6368 30175 6420 30184
rect 6368 30141 6377 30175
rect 6377 30141 6411 30175
rect 6411 30141 6420 30175
rect 6368 30132 6420 30141
rect 8944 30200 8996 30252
rect 9220 30200 9272 30252
rect 9956 30200 10008 30252
rect 8208 29996 8260 30048
rect 9772 30132 9824 30184
rect 10508 30200 10560 30252
rect 11980 30200 12032 30252
rect 14924 30336 14976 30388
rect 15016 30336 15068 30388
rect 17316 30336 17368 30388
rect 18420 30336 18472 30388
rect 18972 30336 19024 30388
rect 12440 30268 12492 30320
rect 12900 30268 12952 30320
rect 14740 30268 14792 30320
rect 14832 30311 14884 30320
rect 14832 30277 14841 30311
rect 14841 30277 14875 30311
rect 14875 30277 14884 30311
rect 14832 30268 14884 30277
rect 16672 30268 16724 30320
rect 13452 30200 13504 30252
rect 14372 30200 14424 30252
rect 15016 30243 15068 30252
rect 15016 30209 15025 30243
rect 15025 30209 15059 30243
rect 15059 30209 15068 30243
rect 15016 30200 15068 30209
rect 10968 30064 11020 30116
rect 14004 30064 14056 30116
rect 10508 29996 10560 30048
rect 12900 30039 12952 30048
rect 12900 30005 12909 30039
rect 12909 30005 12943 30039
rect 12943 30005 12952 30039
rect 12900 29996 12952 30005
rect 14740 30064 14792 30116
rect 15292 30200 15344 30252
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 16580 30132 16632 30184
rect 17224 30243 17276 30252
rect 17224 30209 17233 30243
rect 17233 30209 17267 30243
rect 17267 30209 17276 30243
rect 17224 30200 17276 30209
rect 17684 30200 17736 30252
rect 17960 30311 18012 30320
rect 17960 30277 17969 30311
rect 17969 30277 18003 30311
rect 18003 30277 18012 30311
rect 17960 30268 18012 30277
rect 18788 30268 18840 30320
rect 20076 30268 20128 30320
rect 20536 30268 20588 30320
rect 20628 30311 20680 30320
rect 20628 30277 20637 30311
rect 20637 30277 20671 30311
rect 20671 30277 20680 30311
rect 20628 30268 20680 30277
rect 20812 30268 20864 30320
rect 21088 30311 21140 30320
rect 21088 30277 21097 30311
rect 21097 30277 21131 30311
rect 21131 30277 21140 30311
rect 21088 30268 21140 30277
rect 21824 30336 21876 30388
rect 22744 30336 22796 30388
rect 25044 30336 25096 30388
rect 25688 30336 25740 30388
rect 26148 30336 26200 30388
rect 21272 30311 21324 30320
rect 21272 30277 21281 30311
rect 21281 30277 21315 30311
rect 21315 30277 21324 30311
rect 21272 30268 21324 30277
rect 21456 30268 21508 30320
rect 18236 30200 18288 30252
rect 18788 30132 18840 30184
rect 19892 30200 19944 30252
rect 20168 30243 20220 30252
rect 20168 30209 20177 30243
rect 20177 30209 20211 30243
rect 20211 30209 20220 30243
rect 20168 30200 20220 30209
rect 20260 30243 20312 30252
rect 20260 30209 20269 30243
rect 20269 30209 20303 30243
rect 20303 30209 20312 30243
rect 20260 30200 20312 30209
rect 20720 30200 20772 30252
rect 25504 30243 25556 30252
rect 25504 30209 25513 30243
rect 25513 30209 25547 30243
rect 25547 30209 25556 30243
rect 25504 30200 25556 30209
rect 25688 30243 25740 30252
rect 25688 30209 25697 30243
rect 25697 30209 25731 30243
rect 25731 30209 25740 30243
rect 25688 30200 25740 30209
rect 26056 30200 26108 30252
rect 26332 30132 26384 30184
rect 19156 30064 19208 30116
rect 19708 30064 19760 30116
rect 17960 29996 18012 30048
rect 18512 29996 18564 30048
rect 19800 30039 19852 30048
rect 19800 30005 19809 30039
rect 19809 30005 19843 30039
rect 19843 30005 19852 30039
rect 19800 29996 19852 30005
rect 20352 29996 20404 30048
rect 21272 30039 21324 30048
rect 21272 30005 21281 30039
rect 21281 30005 21315 30039
rect 21315 30005 21324 30039
rect 21272 29996 21324 30005
rect 21640 29996 21692 30048
rect 22652 30064 22704 30116
rect 23204 30064 23256 30116
rect 24308 30064 24360 30116
rect 24676 30107 24728 30116
rect 24676 30073 24685 30107
rect 24685 30073 24719 30107
rect 24719 30073 24728 30107
rect 24676 30064 24728 30073
rect 22928 29996 22980 30048
rect 23112 29996 23164 30048
rect 25872 30039 25924 30048
rect 25872 30005 25881 30039
rect 25881 30005 25915 30039
rect 25915 30005 25924 30039
rect 25872 29996 25924 30005
rect 26056 30039 26108 30048
rect 26056 30005 26065 30039
rect 26065 30005 26099 30039
rect 26099 30005 26108 30039
rect 26056 29996 26108 30005
rect 27160 30268 27212 30320
rect 28540 30268 28592 30320
rect 29276 30268 29328 30320
rect 32496 30336 32548 30388
rect 34336 30336 34388 30388
rect 30840 30268 30892 30320
rect 30748 30200 30800 30252
rect 33140 30268 33192 30320
rect 34520 30268 34572 30320
rect 26700 30175 26752 30184
rect 26700 30141 26709 30175
rect 26709 30141 26743 30175
rect 26743 30141 26752 30175
rect 26700 30132 26752 30141
rect 26884 30132 26936 30184
rect 26976 30175 27028 30184
rect 26976 30141 26985 30175
rect 26985 30141 27019 30175
rect 27019 30141 27028 30175
rect 26976 30132 27028 30141
rect 27252 30175 27304 30184
rect 27252 30141 27261 30175
rect 27261 30141 27295 30175
rect 27295 30141 27304 30175
rect 27252 30132 27304 30141
rect 27896 30132 27948 30184
rect 29092 30175 29144 30184
rect 29092 30141 29101 30175
rect 29101 30141 29135 30175
rect 29135 30141 29144 30175
rect 29092 30132 29144 30141
rect 29828 29996 29880 30048
rect 31024 30039 31076 30048
rect 31024 30005 31033 30039
rect 31033 30005 31067 30039
rect 31067 30005 31076 30039
rect 31024 29996 31076 30005
rect 32404 30175 32456 30184
rect 32404 30141 32413 30175
rect 32413 30141 32447 30175
rect 32447 30141 32456 30175
rect 32404 30132 32456 30141
rect 33784 30132 33836 30184
rect 34244 30132 34296 30184
rect 31668 29996 31720 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12532 29835 12584 29844
rect 12532 29801 12541 29835
rect 12541 29801 12575 29835
rect 12575 29801 12584 29835
rect 12532 29792 12584 29801
rect 12900 29792 12952 29844
rect 16948 29792 17000 29844
rect 17500 29792 17552 29844
rect 19708 29792 19760 29844
rect 20076 29835 20128 29844
rect 20076 29801 20085 29835
rect 20085 29801 20119 29835
rect 20119 29801 20128 29835
rect 20076 29792 20128 29801
rect 20168 29792 20220 29844
rect 20352 29792 20404 29844
rect 20720 29792 20772 29844
rect 25228 29792 25280 29844
rect 25780 29792 25832 29844
rect 25872 29792 25924 29844
rect 26056 29792 26108 29844
rect 26332 29792 26384 29844
rect 27252 29792 27304 29844
rect 28816 29792 28868 29844
rect 30748 29792 30800 29844
rect 8024 29724 8076 29776
rect 9128 29724 9180 29776
rect 5724 29631 5776 29640
rect 5724 29597 5733 29631
rect 5733 29597 5767 29631
rect 5767 29597 5776 29631
rect 5724 29588 5776 29597
rect 6644 29588 6696 29640
rect 6276 29563 6328 29572
rect 6276 29529 6285 29563
rect 6285 29529 6319 29563
rect 6319 29529 6328 29563
rect 6276 29520 6328 29529
rect 9128 29520 9180 29572
rect 10324 29520 10376 29572
rect 12348 29631 12400 29640
rect 12348 29597 12357 29631
rect 12357 29597 12391 29631
rect 12391 29597 12400 29631
rect 12348 29588 12400 29597
rect 15568 29656 15620 29708
rect 13636 29631 13688 29640
rect 13636 29597 13645 29631
rect 13645 29597 13679 29631
rect 13679 29597 13688 29631
rect 13636 29588 13688 29597
rect 13912 29631 13964 29640
rect 13912 29597 13921 29631
rect 13921 29597 13955 29631
rect 13955 29597 13964 29631
rect 13912 29588 13964 29597
rect 14556 29588 14608 29640
rect 15292 29631 15344 29640
rect 15292 29597 15301 29631
rect 15301 29597 15335 29631
rect 15335 29597 15344 29631
rect 15292 29588 15344 29597
rect 15752 29588 15804 29640
rect 15568 29520 15620 29572
rect 4528 29495 4580 29504
rect 4528 29461 4537 29495
rect 4537 29461 4571 29495
rect 4571 29461 4580 29495
rect 4528 29452 4580 29461
rect 7656 29495 7708 29504
rect 7656 29461 7665 29495
rect 7665 29461 7699 29495
rect 7699 29461 7708 29495
rect 7656 29452 7708 29461
rect 8484 29452 8536 29504
rect 9680 29495 9732 29504
rect 9680 29461 9689 29495
rect 9689 29461 9723 29495
rect 9723 29461 9732 29495
rect 9680 29452 9732 29461
rect 11980 29452 12032 29504
rect 12900 29452 12952 29504
rect 13360 29495 13412 29504
rect 13360 29461 13369 29495
rect 13369 29461 13403 29495
rect 13403 29461 13412 29495
rect 13360 29452 13412 29461
rect 16120 29588 16172 29640
rect 21824 29724 21876 29776
rect 22008 29724 22060 29776
rect 23296 29724 23348 29776
rect 18512 29656 18564 29708
rect 18788 29656 18840 29708
rect 19616 29656 19668 29708
rect 16580 29588 16632 29640
rect 17132 29588 17184 29640
rect 17960 29588 18012 29640
rect 16212 29520 16264 29572
rect 19156 29588 19208 29640
rect 19248 29520 19300 29572
rect 19984 29588 20036 29640
rect 20168 29656 20220 29708
rect 20260 29588 20312 29640
rect 20812 29656 20864 29708
rect 24216 29656 24268 29708
rect 20536 29520 20588 29572
rect 22008 29520 22060 29572
rect 22468 29563 22520 29572
rect 22468 29529 22477 29563
rect 22477 29529 22511 29563
rect 22511 29529 22520 29563
rect 22468 29520 22520 29529
rect 22928 29588 22980 29640
rect 23112 29588 23164 29640
rect 23848 29588 23900 29640
rect 25412 29588 25464 29640
rect 34520 29792 34572 29844
rect 26516 29656 26568 29708
rect 15936 29452 15988 29504
rect 16396 29452 16448 29504
rect 16672 29452 16724 29504
rect 17408 29452 17460 29504
rect 17960 29495 18012 29504
rect 17960 29461 17969 29495
rect 17969 29461 18003 29495
rect 18003 29461 18012 29495
rect 17960 29452 18012 29461
rect 18236 29452 18288 29504
rect 18512 29452 18564 29504
rect 19340 29452 19392 29504
rect 19616 29452 19668 29504
rect 21180 29452 21232 29504
rect 26516 29520 26568 29572
rect 28908 29699 28960 29708
rect 28908 29665 28917 29699
rect 28917 29665 28951 29699
rect 28951 29665 28960 29699
rect 28908 29656 28960 29665
rect 30104 29656 30156 29708
rect 29460 29588 29512 29640
rect 29828 29631 29880 29640
rect 29828 29597 29838 29631
rect 29838 29597 29872 29631
rect 29872 29597 29880 29631
rect 29828 29588 29880 29597
rect 30012 29563 30064 29572
rect 30012 29529 30021 29563
rect 30021 29529 30055 29563
rect 30055 29529 30064 29563
rect 30012 29520 30064 29529
rect 31024 29656 31076 29708
rect 30656 29631 30708 29640
rect 30656 29597 30665 29631
rect 30665 29597 30699 29631
rect 30699 29597 30708 29631
rect 30656 29588 30708 29597
rect 30380 29520 30432 29572
rect 22836 29495 22888 29504
rect 22836 29461 22845 29495
rect 22845 29461 22879 29495
rect 22879 29461 22888 29495
rect 22836 29452 22888 29461
rect 23664 29452 23716 29504
rect 25504 29452 25556 29504
rect 25780 29452 25832 29504
rect 27988 29452 28040 29504
rect 28908 29452 28960 29504
rect 31760 29588 31812 29640
rect 32220 29588 32272 29640
rect 32864 29520 32916 29572
rect 32956 29563 33008 29572
rect 32956 29529 32965 29563
rect 32965 29529 32999 29563
rect 32999 29529 33008 29563
rect 32956 29520 33008 29529
rect 34336 29699 34388 29708
rect 34336 29665 34345 29699
rect 34345 29665 34379 29699
rect 34379 29665 34388 29699
rect 34336 29656 34388 29665
rect 34704 29631 34756 29640
rect 34704 29597 34713 29631
rect 34713 29597 34747 29631
rect 34747 29597 34756 29631
rect 34704 29588 34756 29597
rect 32496 29452 32548 29504
rect 34244 29495 34296 29504
rect 34244 29461 34253 29495
rect 34253 29461 34287 29495
rect 34287 29461 34296 29495
rect 34244 29452 34296 29461
rect 34796 29495 34848 29504
rect 34796 29461 34805 29495
rect 34805 29461 34839 29495
rect 34839 29461 34848 29495
rect 34796 29452 34848 29461
rect 34980 29495 35032 29504
rect 34980 29461 34989 29495
rect 34989 29461 35023 29495
rect 35023 29461 35032 29495
rect 34980 29452 35032 29461
rect 36360 29452 36412 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4528 29248 4580 29300
rect 16304 29248 16356 29300
rect 17960 29248 18012 29300
rect 6276 29112 6328 29164
rect 6736 29155 6788 29164
rect 6736 29121 6745 29155
rect 6745 29121 6779 29155
rect 6779 29121 6788 29155
rect 6736 29112 6788 29121
rect 7656 29180 7708 29232
rect 9128 29180 9180 29232
rect 9680 29180 9732 29232
rect 10324 29180 10376 29232
rect 12256 29180 12308 29232
rect 14004 29180 14056 29232
rect 12348 29112 12400 29164
rect 6644 29044 6696 29096
rect 7380 29044 7432 29096
rect 7748 29087 7800 29096
rect 7748 29053 7757 29087
rect 7757 29053 7791 29087
rect 7791 29053 7800 29087
rect 7748 29044 7800 29053
rect 7840 29044 7892 29096
rect 11520 29087 11572 29096
rect 11520 29053 11529 29087
rect 11529 29053 11563 29087
rect 11563 29053 11572 29087
rect 11520 29044 11572 29053
rect 11888 29044 11940 29096
rect 12072 29044 12124 29096
rect 16212 29180 16264 29232
rect 14188 29112 14240 29164
rect 14924 29112 14976 29164
rect 13360 29019 13412 29028
rect 13360 28985 13369 29019
rect 13369 28985 13403 29019
rect 13403 28985 13412 29019
rect 13360 28976 13412 28985
rect 16212 28976 16264 29028
rect 16672 28976 16724 29028
rect 18052 29019 18104 29028
rect 18052 28985 18061 29019
rect 18061 28985 18095 29019
rect 18095 28985 18104 29019
rect 18052 28976 18104 28985
rect 18512 29112 18564 29164
rect 18788 29248 18840 29300
rect 19064 29248 19116 29300
rect 21916 29248 21968 29300
rect 22008 29248 22060 29300
rect 22468 29248 22520 29300
rect 22560 29248 22612 29300
rect 22836 29248 22888 29300
rect 23848 29248 23900 29300
rect 25412 29248 25464 29300
rect 19248 29180 19300 29232
rect 20720 29112 20772 29164
rect 21548 29112 21600 29164
rect 22008 29155 22060 29164
rect 22008 29121 22017 29155
rect 22017 29121 22051 29155
rect 22051 29121 22060 29155
rect 22008 29112 22060 29121
rect 22284 29155 22336 29164
rect 22284 29121 22293 29155
rect 22293 29121 22327 29155
rect 22327 29121 22336 29155
rect 22284 29112 22336 29121
rect 22376 29112 22428 29164
rect 22468 29155 22520 29164
rect 22468 29121 22477 29155
rect 22477 29121 22511 29155
rect 22511 29121 22520 29155
rect 22468 29112 22520 29121
rect 22560 29155 22612 29164
rect 22560 29121 22569 29155
rect 22569 29121 22603 29155
rect 22603 29121 22612 29155
rect 22560 29112 22612 29121
rect 22652 29155 22704 29164
rect 22652 29121 22661 29155
rect 22661 29121 22695 29155
rect 22695 29121 22704 29155
rect 22652 29112 22704 29121
rect 23572 29112 23624 29164
rect 23664 29155 23716 29164
rect 23664 29121 23673 29155
rect 23673 29121 23707 29155
rect 23707 29121 23716 29155
rect 23664 29112 23716 29121
rect 24032 29112 24084 29164
rect 19064 29044 19116 29096
rect 25412 29155 25464 29164
rect 25412 29121 25421 29155
rect 25421 29121 25455 29155
rect 25455 29121 25464 29155
rect 25412 29112 25464 29121
rect 25504 29155 25556 29164
rect 25504 29121 25513 29155
rect 25513 29121 25547 29155
rect 25547 29121 25556 29155
rect 25504 29112 25556 29121
rect 21272 28976 21324 29028
rect 22100 28976 22152 29028
rect 24216 28976 24268 29028
rect 25228 28976 25280 29028
rect 25320 28976 25372 29028
rect 28724 29248 28776 29300
rect 29920 29291 29972 29300
rect 29920 29257 29929 29291
rect 29929 29257 29963 29291
rect 29963 29257 29972 29291
rect 29920 29248 29972 29257
rect 30380 29248 30432 29300
rect 31024 29248 31076 29300
rect 31300 29248 31352 29300
rect 31668 29248 31720 29300
rect 32956 29248 33008 29300
rect 34704 29248 34756 29300
rect 34796 29248 34848 29300
rect 31760 29180 31812 29232
rect 31944 29180 31996 29232
rect 32496 29223 32548 29232
rect 32496 29189 32505 29223
rect 32505 29189 32539 29223
rect 32539 29189 32548 29223
rect 32496 29180 32548 29189
rect 31576 29155 31628 29164
rect 31576 29121 31585 29155
rect 31585 29121 31619 29155
rect 31619 29121 31628 29155
rect 31576 29112 31628 29121
rect 34888 29180 34940 29232
rect 36360 29223 36412 29232
rect 36360 29189 36369 29223
rect 36369 29189 36403 29223
rect 36403 29189 36412 29223
rect 36360 29180 36412 29189
rect 36636 29155 36688 29164
rect 36636 29121 36645 29155
rect 36645 29121 36679 29155
rect 36679 29121 36688 29155
rect 36636 29112 36688 29121
rect 36820 29155 36872 29164
rect 36820 29121 36829 29155
rect 36829 29121 36863 29155
rect 36863 29121 36872 29155
rect 36820 29112 36872 29121
rect 28908 29044 28960 29096
rect 32312 29044 32364 29096
rect 32772 29087 32824 29096
rect 32772 29053 32781 29087
rect 32781 29053 32815 29087
rect 32815 29053 32824 29087
rect 32772 29044 32824 29053
rect 33416 29044 33468 29096
rect 34980 29044 35032 29096
rect 4988 28908 5040 28960
rect 6368 28951 6420 28960
rect 6368 28917 6377 28951
rect 6377 28917 6411 28951
rect 6411 28917 6420 28951
rect 6368 28908 6420 28917
rect 9128 28908 9180 28960
rect 10232 28908 10284 28960
rect 10416 28908 10468 28960
rect 13084 28908 13136 28960
rect 13636 28908 13688 28960
rect 16028 28908 16080 28960
rect 17224 28908 17276 28960
rect 18512 28908 18564 28960
rect 20076 28908 20128 28960
rect 20628 28908 20680 28960
rect 22652 28908 22704 28960
rect 23480 28908 23532 28960
rect 27988 28976 28040 29028
rect 31944 28976 31996 29028
rect 37280 28976 37332 29028
rect 26700 28908 26752 28960
rect 27068 28951 27120 28960
rect 27068 28917 27077 28951
rect 27077 28917 27111 28951
rect 27111 28917 27120 28951
rect 27068 28908 27120 28917
rect 29000 28908 29052 28960
rect 29552 28908 29604 28960
rect 31484 28908 31536 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4988 28747 5040 28756
rect 4988 28713 4997 28747
rect 4997 28713 5031 28747
rect 5031 28713 5040 28747
rect 4988 28704 5040 28713
rect 7748 28704 7800 28756
rect 10232 28704 10284 28756
rect 12440 28704 12492 28756
rect 13084 28704 13136 28756
rect 15568 28704 15620 28756
rect 20720 28704 20772 28756
rect 7840 28636 7892 28688
rect 8392 28636 8444 28688
rect 10508 28636 10560 28688
rect 11152 28636 11204 28688
rect 19432 28636 19484 28688
rect 33692 28704 33744 28756
rect 6368 28568 6420 28620
rect 5356 28500 5408 28552
rect 8024 28568 8076 28620
rect 1768 28407 1820 28416
rect 1768 28373 1777 28407
rect 1777 28373 1811 28407
rect 1811 28373 1820 28407
rect 1768 28364 1820 28373
rect 4344 28407 4396 28416
rect 4344 28373 4353 28407
rect 4353 28373 4387 28407
rect 4387 28373 4396 28407
rect 4344 28364 4396 28373
rect 6920 28407 6972 28416
rect 6920 28373 6929 28407
rect 6929 28373 6963 28407
rect 6963 28373 6972 28407
rect 6920 28364 6972 28373
rect 8392 28543 8444 28552
rect 8392 28509 8401 28543
rect 8401 28509 8435 28543
rect 8435 28509 8444 28543
rect 8392 28500 8444 28509
rect 8944 28500 8996 28552
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 8852 28432 8904 28484
rect 10416 28543 10468 28552
rect 10416 28509 10425 28543
rect 10425 28509 10459 28543
rect 10459 28509 10468 28543
rect 10416 28500 10468 28509
rect 10508 28543 10560 28552
rect 10508 28509 10517 28543
rect 10517 28509 10551 28543
rect 10551 28509 10560 28543
rect 10508 28500 10560 28509
rect 10876 28500 10928 28552
rect 10968 28543 11020 28552
rect 10968 28509 10977 28543
rect 10977 28509 11011 28543
rect 11011 28509 11020 28543
rect 10968 28500 11020 28509
rect 10324 28475 10376 28484
rect 10324 28441 10333 28475
rect 10333 28441 10367 28475
rect 10367 28441 10376 28475
rect 10324 28432 10376 28441
rect 11428 28500 11480 28552
rect 14188 28568 14240 28620
rect 20352 28611 20404 28620
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 16856 28500 16908 28552
rect 17224 28543 17276 28552
rect 17224 28509 17233 28543
rect 17233 28509 17267 28543
rect 17267 28509 17276 28543
rect 17224 28500 17276 28509
rect 20352 28577 20361 28611
rect 20361 28577 20395 28611
rect 20395 28577 20404 28611
rect 20352 28568 20404 28577
rect 17960 28500 18012 28552
rect 19340 28500 19392 28552
rect 20260 28543 20312 28552
rect 20260 28509 20269 28543
rect 20269 28509 20303 28543
rect 20303 28509 20312 28543
rect 20260 28500 20312 28509
rect 11060 28364 11112 28416
rect 20352 28432 20404 28484
rect 20536 28543 20588 28552
rect 20536 28509 20545 28543
rect 20545 28509 20579 28543
rect 20579 28509 20588 28543
rect 20536 28500 20588 28509
rect 23388 28568 23440 28620
rect 22008 28432 22060 28484
rect 23020 28475 23072 28484
rect 23020 28441 23029 28475
rect 23029 28441 23063 28475
rect 23063 28441 23072 28475
rect 23020 28432 23072 28441
rect 11704 28407 11756 28416
rect 11704 28373 11713 28407
rect 11713 28373 11747 28407
rect 11747 28373 11756 28407
rect 11704 28364 11756 28373
rect 17868 28407 17920 28416
rect 17868 28373 17877 28407
rect 17877 28373 17911 28407
rect 17911 28373 17920 28407
rect 17868 28364 17920 28373
rect 19984 28364 20036 28416
rect 22652 28364 22704 28416
rect 23296 28432 23348 28484
rect 24216 28679 24268 28688
rect 24216 28645 24225 28679
rect 24225 28645 24259 28679
rect 24259 28645 24268 28679
rect 24216 28636 24268 28645
rect 26516 28636 26568 28688
rect 23848 28543 23900 28552
rect 23848 28509 23857 28543
rect 23857 28509 23891 28543
rect 23891 28509 23900 28543
rect 23848 28500 23900 28509
rect 24216 28500 24268 28552
rect 24492 28500 24544 28552
rect 23204 28364 23256 28416
rect 25504 28500 25556 28552
rect 27068 28568 27120 28620
rect 25872 28500 25924 28552
rect 26240 28543 26292 28552
rect 26240 28509 26249 28543
rect 26249 28509 26283 28543
rect 26283 28509 26292 28543
rect 26240 28500 26292 28509
rect 26332 28543 26384 28552
rect 26332 28509 26341 28543
rect 26341 28509 26375 28543
rect 26375 28509 26384 28543
rect 26332 28500 26384 28509
rect 25688 28475 25740 28484
rect 25688 28441 25697 28475
rect 25697 28441 25731 28475
rect 25731 28441 25740 28475
rect 25688 28432 25740 28441
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 25780 28364 25832 28416
rect 27068 28475 27120 28484
rect 27068 28441 27077 28475
rect 27077 28441 27111 28475
rect 27111 28441 27120 28475
rect 27068 28432 27120 28441
rect 26056 28407 26108 28416
rect 26056 28373 26065 28407
rect 26065 28373 26099 28407
rect 26099 28373 26108 28407
rect 26056 28364 26108 28373
rect 27896 28364 27948 28416
rect 28954 28636 29006 28688
rect 29092 28500 29144 28552
rect 29184 28525 29193 28552
rect 29193 28525 29227 28552
rect 29227 28525 29236 28552
rect 29184 28500 29236 28525
rect 33140 28568 33192 28620
rect 34796 28568 34848 28620
rect 31484 28543 31536 28552
rect 31484 28509 31493 28543
rect 31493 28509 31527 28543
rect 31527 28509 31536 28543
rect 31484 28500 31536 28509
rect 33048 28500 33100 28552
rect 28540 28407 28592 28416
rect 28540 28373 28549 28407
rect 28549 28373 28583 28407
rect 28583 28373 28592 28407
rect 28540 28364 28592 28373
rect 31392 28432 31444 28484
rect 31760 28475 31812 28484
rect 31760 28441 31769 28475
rect 31769 28441 31803 28475
rect 31803 28441 31812 28475
rect 31760 28432 31812 28441
rect 29736 28364 29788 28416
rect 33508 28432 33560 28484
rect 33140 28364 33192 28416
rect 33232 28407 33284 28416
rect 33232 28373 33241 28407
rect 33241 28373 33275 28407
rect 33275 28373 33284 28407
rect 33232 28364 33284 28373
rect 34244 28407 34296 28416
rect 34244 28373 34253 28407
rect 34253 28373 34287 28407
rect 34287 28373 34296 28407
rect 34244 28364 34296 28373
rect 34520 28364 34572 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4344 28160 4396 28212
rect 6920 28160 6972 28212
rect 9128 28160 9180 28212
rect 4712 28092 4764 28144
rect 6276 28092 6328 28144
rect 8116 28024 8168 28076
rect 11336 28067 11388 28076
rect 11336 28033 11345 28067
rect 11345 28033 11379 28067
rect 11379 28033 11388 28067
rect 11336 28024 11388 28033
rect 11704 28092 11756 28144
rect 12256 28092 12308 28144
rect 14556 28135 14608 28144
rect 14556 28101 14565 28135
rect 14565 28101 14599 28135
rect 14599 28101 14608 28135
rect 14556 28092 14608 28101
rect 14648 28092 14700 28144
rect 14372 28067 14424 28076
rect 14372 28033 14381 28067
rect 14381 28033 14415 28067
rect 14415 28033 14424 28067
rect 14372 28024 14424 28033
rect 14740 28024 14792 28076
rect 15200 28024 15252 28076
rect 7012 27999 7064 28008
rect 7012 27965 7021 27999
rect 7021 27965 7055 27999
rect 7055 27965 7064 27999
rect 7012 27956 7064 27965
rect 5908 27863 5960 27872
rect 5908 27829 5917 27863
rect 5917 27829 5951 27863
rect 5951 27829 5960 27863
rect 11060 27888 11112 27940
rect 13268 27999 13320 28008
rect 13268 27965 13277 27999
rect 13277 27965 13311 27999
rect 13311 27965 13320 27999
rect 16488 28092 16540 28144
rect 13268 27956 13320 27965
rect 16120 28024 16172 28076
rect 17408 28067 17460 28076
rect 17408 28033 17417 28067
rect 17417 28033 17451 28067
rect 17451 28033 17460 28067
rect 17408 28024 17460 28033
rect 17500 28067 17552 28076
rect 17500 28033 17509 28067
rect 17509 28033 17543 28067
rect 17543 28033 17552 28067
rect 17500 28024 17552 28033
rect 17960 28160 18012 28212
rect 18788 28160 18840 28212
rect 17776 28092 17828 28144
rect 18144 28024 18196 28076
rect 20536 28160 20588 28212
rect 20076 28024 20128 28076
rect 20168 28067 20220 28076
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 20352 28092 20404 28144
rect 20720 28092 20772 28144
rect 21088 28160 21140 28212
rect 22008 28203 22060 28212
rect 22008 28169 22017 28203
rect 22017 28169 22051 28203
rect 22051 28169 22060 28203
rect 22008 28160 22060 28169
rect 22100 28203 22152 28212
rect 22100 28169 22109 28203
rect 22109 28169 22143 28203
rect 22143 28169 22152 28203
rect 22100 28160 22152 28169
rect 22744 28160 22796 28212
rect 22928 28160 22980 28212
rect 21824 28135 21876 28144
rect 21824 28101 21833 28135
rect 21833 28101 21867 28135
rect 21867 28101 21876 28135
rect 21824 28092 21876 28101
rect 22560 28092 22612 28144
rect 21272 28067 21324 28076
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 21272 28024 21324 28033
rect 22284 28024 22336 28076
rect 22928 28067 22980 28076
rect 22928 28033 22937 28067
rect 22937 28033 22971 28067
rect 22971 28033 22980 28067
rect 22928 28024 22980 28033
rect 14188 27931 14240 27940
rect 14188 27897 14197 27931
rect 14197 27897 14231 27931
rect 14231 27897 14240 27931
rect 14188 27888 14240 27897
rect 14556 27888 14608 27940
rect 15384 27888 15436 27940
rect 16304 27888 16356 27940
rect 19432 27888 19484 27940
rect 19800 27931 19852 27940
rect 19800 27897 19809 27931
rect 19809 27897 19843 27931
rect 19843 27897 19852 27931
rect 19800 27888 19852 27897
rect 19984 27888 20036 27940
rect 21456 27956 21508 28008
rect 21732 27956 21784 28008
rect 23112 28067 23164 28076
rect 23112 28033 23126 28067
rect 23126 28033 23160 28067
rect 23160 28033 23164 28067
rect 23112 28024 23164 28033
rect 23296 28024 23348 28076
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 23572 28092 23624 28144
rect 23940 28092 23992 28144
rect 22376 27888 22428 27940
rect 22652 27888 22704 27940
rect 22928 27888 22980 27940
rect 5908 27820 5960 27829
rect 8392 27820 8444 27872
rect 11520 27820 11572 27872
rect 16764 27820 16816 27872
rect 17224 27820 17276 27872
rect 19340 27820 19392 27872
rect 19524 27863 19576 27872
rect 19524 27829 19533 27863
rect 19533 27829 19567 27863
rect 19567 27829 19576 27863
rect 19524 27820 19576 27829
rect 20996 27863 21048 27872
rect 20996 27829 21005 27863
rect 21005 27829 21039 27863
rect 21039 27829 21048 27863
rect 20996 27820 21048 27829
rect 21456 27863 21508 27872
rect 21456 27829 21465 27863
rect 21465 27829 21499 27863
rect 21499 27829 21508 27863
rect 21456 27820 21508 27829
rect 21640 27820 21692 27872
rect 25412 28160 25464 28212
rect 26056 28160 26108 28212
rect 24124 28024 24176 28076
rect 26148 28067 26200 28076
rect 26148 28033 26157 28067
rect 26157 28033 26191 28067
rect 26191 28033 26200 28067
rect 26148 28024 26200 28033
rect 27068 28203 27120 28212
rect 27068 28169 27077 28203
rect 27077 28169 27111 28203
rect 27111 28169 27120 28203
rect 27068 28160 27120 28169
rect 29184 28160 29236 28212
rect 26976 28092 27028 28144
rect 26700 28024 26752 28076
rect 26792 28024 26844 28076
rect 27252 28067 27304 28076
rect 27252 28033 27261 28067
rect 27261 28033 27295 28067
rect 27295 28033 27304 28067
rect 27252 28024 27304 28033
rect 29000 28048 29052 28100
rect 29092 28067 29144 28076
rect 29092 28033 29101 28067
rect 29101 28033 29135 28067
rect 29135 28033 29144 28067
rect 29092 28024 29144 28033
rect 29920 28135 29972 28144
rect 29920 28101 29929 28135
rect 29929 28101 29963 28135
rect 29963 28101 29972 28135
rect 29920 28092 29972 28101
rect 30012 28135 30064 28144
rect 30012 28101 30021 28135
rect 30021 28101 30055 28135
rect 30055 28101 30064 28135
rect 30012 28092 30064 28101
rect 28816 27956 28868 28008
rect 26332 27888 26384 27940
rect 29460 28024 29512 28076
rect 29736 28067 29788 28076
rect 29736 28033 29746 28067
rect 29746 28033 29780 28067
rect 29780 28033 29788 28067
rect 29736 28024 29788 28033
rect 30104 28067 30156 28076
rect 30104 28033 30118 28067
rect 30118 28033 30152 28067
rect 30152 28033 30156 28067
rect 31760 28203 31812 28212
rect 31760 28169 31769 28203
rect 31769 28169 31803 28203
rect 31803 28169 31812 28203
rect 31760 28160 31812 28169
rect 30380 28092 30432 28144
rect 30104 28024 30156 28033
rect 30840 28067 30892 28076
rect 30840 28033 30849 28067
rect 30849 28033 30883 28067
rect 30883 28033 30892 28067
rect 30840 28024 30892 28033
rect 34244 28160 34296 28212
rect 33968 28092 34020 28144
rect 34520 28160 34572 28212
rect 32496 28067 32548 28076
rect 32496 28033 32505 28067
rect 32505 28033 32539 28067
rect 32539 28033 32548 28067
rect 32496 28024 32548 28033
rect 33232 28024 33284 28076
rect 33508 28024 33560 28076
rect 34796 28092 34848 28144
rect 32772 27999 32824 28008
rect 32772 27965 32781 27999
rect 32781 27965 32815 27999
rect 32815 27965 32824 27999
rect 32772 27956 32824 27965
rect 23296 27863 23348 27872
rect 23296 27829 23305 27863
rect 23305 27829 23339 27863
rect 23339 27829 23348 27863
rect 23296 27820 23348 27829
rect 23756 27820 23808 27872
rect 25688 27820 25740 27872
rect 30288 27820 30340 27872
rect 30380 27863 30432 27872
rect 30380 27829 30389 27863
rect 30389 27829 30423 27863
rect 30423 27829 30432 27863
rect 30380 27820 30432 27829
rect 33784 27999 33836 28008
rect 33784 27965 33793 27999
rect 33793 27965 33827 27999
rect 33827 27965 33836 27999
rect 33784 27956 33836 27965
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4712 27659 4764 27668
rect 4712 27625 4721 27659
rect 4721 27625 4755 27659
rect 4755 27625 4764 27659
rect 4712 27616 4764 27625
rect 7012 27616 7064 27668
rect 8116 27616 8168 27668
rect 8668 27616 8720 27668
rect 11336 27616 11388 27668
rect 11796 27616 11848 27668
rect 6828 27480 6880 27532
rect 5908 27412 5960 27464
rect 10600 27548 10652 27600
rect 11704 27548 11756 27600
rect 12072 27548 12124 27600
rect 6736 27344 6788 27396
rect 8392 27412 8444 27464
rect 8484 27455 8536 27464
rect 8484 27421 8493 27455
rect 8493 27421 8527 27455
rect 8527 27421 8536 27455
rect 8484 27412 8536 27421
rect 8852 27480 8904 27532
rect 10692 27480 10744 27532
rect 12348 27480 12400 27532
rect 13268 27548 13320 27600
rect 14556 27591 14608 27600
rect 14556 27557 14565 27591
rect 14565 27557 14599 27591
rect 14599 27557 14608 27591
rect 14556 27548 14608 27557
rect 14648 27548 14700 27600
rect 13820 27480 13872 27532
rect 14188 27480 14240 27532
rect 15660 27480 15712 27532
rect 13636 27412 13688 27464
rect 14464 27412 14516 27464
rect 15476 27412 15528 27464
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 16028 27455 16080 27464
rect 12624 27344 12676 27396
rect 15384 27344 15436 27396
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 16488 27412 16540 27464
rect 16672 27455 16724 27464
rect 16672 27421 16681 27455
rect 16681 27421 16715 27455
rect 16715 27421 16724 27455
rect 16672 27412 16724 27421
rect 17040 27480 17092 27532
rect 17868 27480 17920 27532
rect 15936 27387 15988 27396
rect 15936 27353 15945 27387
rect 15945 27353 15979 27387
rect 15979 27353 15988 27387
rect 15936 27344 15988 27353
rect 8300 27276 8352 27328
rect 9404 27276 9456 27328
rect 10968 27276 11020 27328
rect 11520 27276 11572 27328
rect 11796 27276 11848 27328
rect 13636 27319 13688 27328
rect 13636 27285 13645 27319
rect 13645 27285 13679 27319
rect 13679 27285 13688 27319
rect 13636 27276 13688 27285
rect 14372 27276 14424 27328
rect 14832 27319 14884 27328
rect 14832 27285 14841 27319
rect 14841 27285 14875 27319
rect 14875 27285 14884 27319
rect 14832 27276 14884 27285
rect 15660 27276 15712 27328
rect 17408 27412 17460 27464
rect 19800 27616 19852 27668
rect 20076 27616 20128 27668
rect 20628 27616 20680 27668
rect 21272 27616 21324 27668
rect 24492 27616 24544 27668
rect 25044 27616 25096 27668
rect 26148 27616 26200 27668
rect 26516 27616 26568 27668
rect 27252 27616 27304 27668
rect 29184 27616 29236 27668
rect 32496 27616 32548 27668
rect 33692 27659 33744 27668
rect 33692 27625 33701 27659
rect 33701 27625 33735 27659
rect 33735 27625 33744 27659
rect 33692 27616 33744 27625
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 19524 27412 19576 27464
rect 20076 27412 20128 27464
rect 20444 27412 20496 27464
rect 20812 27455 20864 27464
rect 20812 27421 20821 27455
rect 20821 27421 20855 27455
rect 20855 27421 20864 27455
rect 20812 27412 20864 27421
rect 21088 27412 21140 27464
rect 21456 27480 21508 27532
rect 23296 27523 23348 27532
rect 23296 27489 23305 27523
rect 23305 27489 23339 27523
rect 23339 27489 23348 27523
rect 23296 27480 23348 27489
rect 23756 27480 23808 27532
rect 21824 27412 21876 27464
rect 22192 27412 22244 27464
rect 19984 27344 20036 27396
rect 17132 27276 17184 27328
rect 18052 27276 18104 27328
rect 20996 27344 21048 27396
rect 22560 27455 22612 27464
rect 22560 27421 22569 27455
rect 22569 27421 22603 27455
rect 22603 27421 22612 27455
rect 22560 27412 22612 27421
rect 23204 27455 23256 27464
rect 23204 27421 23213 27455
rect 23213 27421 23247 27455
rect 23247 27421 23256 27455
rect 23204 27412 23256 27421
rect 23388 27344 23440 27396
rect 23664 27455 23716 27464
rect 23664 27421 23673 27455
rect 23673 27421 23707 27455
rect 23707 27421 23716 27455
rect 23664 27412 23716 27421
rect 24124 27412 24176 27464
rect 28908 27548 28960 27600
rect 29920 27548 29972 27600
rect 30380 27548 30432 27600
rect 30656 27548 30708 27600
rect 30840 27548 30892 27600
rect 34704 27548 34756 27600
rect 24584 27480 24636 27532
rect 27528 27412 27580 27464
rect 29092 27412 29144 27464
rect 29368 27412 29420 27464
rect 30748 27455 30800 27464
rect 30748 27421 30757 27455
rect 30757 27421 30791 27455
rect 30791 27421 30800 27455
rect 30748 27412 30800 27421
rect 23020 27276 23072 27328
rect 23572 27276 23624 27328
rect 24400 27276 24452 27328
rect 25596 27276 25648 27328
rect 27804 27344 27856 27396
rect 30840 27344 30892 27396
rect 28632 27276 28684 27328
rect 29460 27276 29512 27328
rect 31024 27455 31076 27464
rect 31024 27421 31033 27455
rect 31033 27421 31067 27455
rect 31067 27421 31076 27455
rect 31024 27412 31076 27421
rect 31208 27412 31260 27464
rect 31300 27344 31352 27396
rect 32404 27412 32456 27464
rect 33784 27276 33836 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 6828 27072 6880 27124
rect 5908 26979 5960 26988
rect 5908 26945 5917 26979
rect 5917 26945 5951 26979
rect 5951 26945 5960 26979
rect 5908 26936 5960 26945
rect 8300 27004 8352 27056
rect 8668 27004 8720 27056
rect 8392 26911 8444 26920
rect 8392 26877 8401 26911
rect 8401 26877 8435 26911
rect 8435 26877 8444 26911
rect 8392 26868 8444 26877
rect 10600 27004 10652 27056
rect 10140 26936 10192 26988
rect 5448 26732 5500 26784
rect 7380 26732 7432 26784
rect 7748 26732 7800 26784
rect 9496 26800 9548 26852
rect 10600 26911 10652 26920
rect 10600 26877 10609 26911
rect 10609 26877 10643 26911
rect 10643 26877 10652 26911
rect 10600 26868 10652 26877
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 11520 27115 11572 27124
rect 11520 27081 11529 27115
rect 11529 27081 11563 27115
rect 11563 27081 11572 27115
rect 11520 27072 11572 27081
rect 15200 27072 15252 27124
rect 16672 27115 16724 27124
rect 16672 27081 16681 27115
rect 16681 27081 16715 27115
rect 16715 27081 16724 27115
rect 16672 27072 16724 27081
rect 16856 27072 16908 27124
rect 16948 27072 17000 27124
rect 11980 27004 12032 27056
rect 12808 27004 12860 27056
rect 11796 26868 11848 26920
rect 12900 26979 12952 26988
rect 12900 26945 12909 26979
rect 12909 26945 12943 26979
rect 12943 26945 12952 26979
rect 12900 26936 12952 26945
rect 13084 27004 13136 27056
rect 13912 27004 13964 27056
rect 13268 26979 13320 26988
rect 13268 26945 13277 26979
rect 13277 26945 13311 26979
rect 13311 26945 13320 26979
rect 13268 26936 13320 26945
rect 13360 26979 13412 26988
rect 13360 26945 13374 26979
rect 13374 26945 13408 26979
rect 13408 26945 13412 26979
rect 13360 26936 13412 26945
rect 13544 26936 13596 26988
rect 13636 26936 13688 26988
rect 14188 26868 14240 26920
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 16120 27004 16172 27056
rect 15844 26936 15896 26988
rect 16028 26936 16080 26988
rect 16764 26936 16816 26988
rect 18144 27072 18196 27124
rect 18328 26979 18380 26988
rect 18328 26945 18337 26979
rect 18337 26945 18371 26979
rect 18371 26945 18380 26979
rect 18328 26936 18380 26945
rect 18420 26979 18472 26988
rect 18420 26945 18429 26979
rect 18429 26945 18463 26979
rect 18463 26945 18472 26979
rect 18420 26936 18472 26945
rect 18696 26936 18748 26988
rect 18788 26979 18840 26988
rect 18788 26945 18797 26979
rect 18797 26945 18831 26979
rect 18831 26945 18840 26979
rect 18788 26936 18840 26945
rect 19064 27047 19116 27056
rect 19064 27013 19073 27047
rect 19073 27013 19107 27047
rect 19107 27013 19116 27047
rect 19064 27004 19116 27013
rect 20720 27072 20772 27124
rect 23756 27072 23808 27124
rect 25872 27072 25924 27124
rect 29552 27072 29604 27124
rect 34704 27072 34756 27124
rect 34796 27072 34848 27124
rect 35348 27072 35400 27124
rect 20996 27004 21048 27056
rect 24400 27004 24452 27056
rect 24860 27004 24912 27056
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 25780 26979 25832 26988
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 27804 27004 27856 27056
rect 28540 27004 28592 27056
rect 10600 26732 10652 26784
rect 10968 26732 11020 26784
rect 12256 26732 12308 26784
rect 26056 26936 26108 26988
rect 27620 26979 27672 26988
rect 27620 26945 27629 26979
rect 27629 26945 27663 26979
rect 27663 26945 27672 26979
rect 27620 26936 27672 26945
rect 28632 26979 28684 26988
rect 28632 26945 28641 26979
rect 28641 26945 28675 26979
rect 28675 26945 28684 26979
rect 28632 26936 28684 26945
rect 28724 26979 28776 26988
rect 28724 26945 28734 26979
rect 28734 26945 28768 26979
rect 28768 26945 28776 26979
rect 28724 26936 28776 26945
rect 28908 26979 28960 26988
rect 28908 26945 28917 26979
rect 28917 26945 28951 26979
rect 28951 26945 28960 26979
rect 28908 26936 28960 26945
rect 30104 26936 30156 26988
rect 30748 26936 30800 26988
rect 31024 26936 31076 26988
rect 34336 26979 34388 26988
rect 34336 26945 34345 26979
rect 34345 26945 34379 26979
rect 34379 26945 34388 26979
rect 34336 26936 34388 26945
rect 13820 26732 13872 26784
rect 14556 26732 14608 26784
rect 18880 26800 18932 26852
rect 18972 26800 19024 26852
rect 19064 26800 19116 26852
rect 30288 26868 30340 26920
rect 16488 26732 16540 26784
rect 24124 26800 24176 26852
rect 31300 26800 31352 26852
rect 19340 26775 19392 26784
rect 19340 26741 19349 26775
rect 19349 26741 19383 26775
rect 19383 26741 19392 26775
rect 19340 26732 19392 26741
rect 21824 26732 21876 26784
rect 22284 26732 22336 26784
rect 25596 26732 25648 26784
rect 26148 26775 26200 26784
rect 26148 26741 26157 26775
rect 26157 26741 26191 26775
rect 26191 26741 26200 26775
rect 26148 26732 26200 26741
rect 27436 26775 27488 26784
rect 27436 26741 27445 26775
rect 27445 26741 27479 26775
rect 27479 26741 27488 26775
rect 27436 26732 27488 26741
rect 29276 26775 29328 26784
rect 29276 26741 29285 26775
rect 29285 26741 29319 26775
rect 29319 26741 29328 26775
rect 29276 26732 29328 26741
rect 32588 26732 32640 26784
rect 34612 26732 34664 26784
rect 34796 26732 34848 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5356 26528 5408 26580
rect 8392 26460 8444 26512
rect 9496 26460 9548 26512
rect 4068 26392 4120 26444
rect 7104 26392 7156 26444
rect 8668 26392 8720 26444
rect 6644 26324 6696 26376
rect 5264 26256 5316 26308
rect 5448 26256 5500 26308
rect 7196 26256 7248 26308
rect 10600 26528 10652 26580
rect 11980 26571 12032 26580
rect 11980 26537 11989 26571
rect 11989 26537 12023 26571
rect 12023 26537 12032 26571
rect 11980 26528 12032 26537
rect 12164 26528 12216 26580
rect 12900 26528 12952 26580
rect 19340 26528 19392 26580
rect 14188 26503 14240 26512
rect 14188 26469 14197 26503
rect 14197 26469 14231 26503
rect 14231 26469 14240 26503
rect 14188 26460 14240 26469
rect 15660 26460 15712 26512
rect 13268 26392 13320 26444
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 14648 26367 14700 26376
rect 14648 26333 14657 26367
rect 14657 26333 14691 26367
rect 14691 26333 14700 26367
rect 14648 26324 14700 26333
rect 14924 26367 14976 26376
rect 14924 26333 14933 26367
rect 14933 26333 14967 26367
rect 14967 26333 14976 26367
rect 14924 26324 14976 26333
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 16580 26367 16632 26376
rect 16580 26333 16589 26367
rect 16589 26333 16623 26367
rect 16623 26333 16632 26367
rect 16580 26324 16632 26333
rect 17132 26367 17184 26376
rect 17132 26333 17142 26367
rect 17142 26333 17176 26367
rect 17176 26333 17184 26367
rect 17132 26324 17184 26333
rect 17316 26367 17368 26376
rect 17316 26333 17325 26367
rect 17325 26333 17359 26367
rect 17359 26333 17368 26367
rect 17316 26324 17368 26333
rect 10968 26256 11020 26308
rect 8944 26188 8996 26240
rect 13084 26188 13136 26240
rect 13360 26188 13412 26240
rect 15752 26256 15804 26308
rect 18788 26392 18840 26444
rect 17684 26324 17736 26376
rect 17776 26367 17828 26376
rect 17776 26333 17785 26367
rect 17785 26333 17819 26367
rect 17819 26333 17828 26367
rect 17776 26324 17828 26333
rect 16304 26188 16356 26240
rect 18420 26324 18472 26376
rect 20904 26324 20956 26376
rect 22192 26528 22244 26580
rect 22468 26460 22520 26512
rect 22744 26460 22796 26512
rect 21456 26392 21508 26444
rect 21180 26367 21232 26376
rect 21180 26333 21189 26367
rect 21189 26333 21223 26367
rect 21223 26333 21232 26367
rect 21180 26324 21232 26333
rect 18144 26231 18196 26240
rect 18144 26197 18153 26231
rect 18153 26197 18187 26231
rect 18187 26197 18196 26231
rect 18144 26188 18196 26197
rect 18880 26256 18932 26308
rect 20076 26256 20128 26308
rect 20536 26256 20588 26308
rect 21548 26256 21600 26308
rect 25872 26392 25924 26444
rect 23296 26324 23348 26376
rect 23848 26324 23900 26376
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 24676 26299 24728 26308
rect 24676 26265 24685 26299
rect 24685 26265 24719 26299
rect 24719 26265 24728 26299
rect 24676 26256 24728 26265
rect 25412 26256 25464 26308
rect 20812 26188 20864 26240
rect 22560 26188 22612 26240
rect 25504 26188 25556 26240
rect 26516 26460 26568 26512
rect 26700 26460 26752 26512
rect 27436 26392 27488 26444
rect 30656 26460 30708 26512
rect 26332 26299 26384 26308
rect 26332 26265 26341 26299
rect 26341 26265 26375 26299
rect 26375 26265 26384 26299
rect 26332 26256 26384 26265
rect 27068 26367 27120 26376
rect 27068 26333 27077 26367
rect 27077 26333 27111 26367
rect 27111 26333 27120 26367
rect 27068 26324 27120 26333
rect 29092 26324 29144 26376
rect 29276 26324 29328 26376
rect 30288 26367 30340 26376
rect 30288 26333 30297 26367
rect 30297 26333 30331 26367
rect 30331 26333 30340 26367
rect 30288 26324 30340 26333
rect 30472 26324 30524 26376
rect 30748 26324 30800 26376
rect 27804 26256 27856 26308
rect 31024 26367 31076 26376
rect 31024 26333 31033 26367
rect 31033 26333 31067 26367
rect 31067 26333 31076 26367
rect 31024 26324 31076 26333
rect 34336 26528 34388 26580
rect 34704 26528 34756 26580
rect 34796 26528 34848 26580
rect 32680 26460 32732 26512
rect 33784 26392 33836 26444
rect 34244 26392 34296 26444
rect 31392 26367 31444 26376
rect 31392 26333 31401 26367
rect 31401 26333 31435 26367
rect 31435 26333 31444 26367
rect 31392 26324 31444 26333
rect 34612 26392 34664 26444
rect 28356 26188 28408 26240
rect 28724 26188 28776 26240
rect 29092 26188 29144 26240
rect 30564 26188 30616 26240
rect 31300 26256 31352 26308
rect 31760 26256 31812 26308
rect 31208 26188 31260 26240
rect 33692 26299 33744 26308
rect 33692 26265 33701 26299
rect 33701 26265 33735 26299
rect 33735 26265 33744 26299
rect 33692 26256 33744 26265
rect 32496 26188 32548 26240
rect 34336 26188 34388 26240
rect 35440 26256 35492 26308
rect 36544 26256 36596 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5908 25984 5960 26036
rect 11060 25984 11112 26036
rect 12164 25984 12216 26036
rect 7196 25916 7248 25968
rect 15384 25984 15436 26036
rect 13728 25916 13780 25968
rect 23204 25984 23256 26036
rect 23480 25984 23532 26036
rect 24676 25984 24728 26036
rect 24952 25984 25004 26036
rect 25136 25984 25188 26036
rect 25872 25984 25924 26036
rect 6000 25891 6052 25900
rect 6000 25857 6009 25891
rect 6009 25857 6043 25891
rect 6043 25857 6052 25891
rect 6000 25848 6052 25857
rect 6828 25780 6880 25832
rect 10416 25891 10468 25900
rect 10416 25857 10425 25891
rect 10425 25857 10459 25891
rect 10459 25857 10468 25891
rect 10416 25848 10468 25857
rect 11888 25891 11940 25900
rect 11888 25857 11897 25891
rect 11897 25857 11931 25891
rect 11931 25857 11940 25891
rect 11888 25848 11940 25857
rect 14648 25848 14700 25900
rect 15108 25848 15160 25900
rect 16120 25848 16172 25900
rect 18236 25891 18288 25900
rect 18236 25857 18245 25891
rect 18245 25857 18279 25891
rect 18279 25857 18288 25891
rect 18236 25848 18288 25857
rect 5632 25644 5684 25696
rect 9404 25712 9456 25764
rect 7932 25644 7984 25696
rect 10048 25644 10100 25696
rect 12072 25687 12124 25696
rect 12072 25653 12081 25687
rect 12081 25653 12115 25687
rect 12115 25653 12124 25687
rect 12072 25644 12124 25653
rect 12624 25712 12676 25764
rect 16028 25712 16080 25764
rect 17960 25780 18012 25832
rect 20352 25916 20404 25968
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 22744 25916 22796 25968
rect 21180 25848 21232 25900
rect 21456 25848 21508 25900
rect 22192 25848 22244 25900
rect 19708 25712 19760 25764
rect 19984 25712 20036 25764
rect 20628 25712 20680 25764
rect 16580 25644 16632 25696
rect 18512 25644 18564 25696
rect 18604 25687 18656 25696
rect 18604 25653 18613 25687
rect 18613 25653 18647 25687
rect 18647 25653 18656 25687
rect 18604 25644 18656 25653
rect 20444 25687 20496 25696
rect 20444 25653 20453 25687
rect 20453 25653 20487 25687
rect 20487 25653 20496 25687
rect 20444 25644 20496 25653
rect 20812 25687 20864 25696
rect 20812 25653 20821 25687
rect 20821 25653 20855 25687
rect 20855 25653 20864 25687
rect 20812 25644 20864 25653
rect 22192 25687 22244 25696
rect 22192 25653 22201 25687
rect 22201 25653 22235 25687
rect 22235 25653 22244 25687
rect 22192 25644 22244 25653
rect 22560 25891 22612 25900
rect 22560 25857 22569 25891
rect 22569 25857 22603 25891
rect 22603 25857 22612 25891
rect 22560 25848 22612 25857
rect 22468 25755 22520 25764
rect 22468 25721 22477 25755
rect 22477 25721 22511 25755
rect 22511 25721 22520 25755
rect 22468 25712 22520 25721
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 23296 25848 23348 25900
rect 23664 25891 23716 25900
rect 23664 25857 23673 25891
rect 23673 25857 23707 25891
rect 23707 25857 23716 25891
rect 23664 25848 23716 25857
rect 25688 25916 25740 25968
rect 23848 25780 23900 25832
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 24768 25848 24820 25900
rect 24952 25848 25004 25900
rect 26240 25984 26292 26036
rect 26608 25984 26660 26036
rect 27068 25984 27120 26036
rect 27620 25984 27672 26036
rect 24124 25823 24176 25832
rect 24124 25789 24133 25823
rect 24133 25789 24167 25823
rect 24167 25789 24176 25823
rect 24124 25780 24176 25789
rect 26148 25848 26200 25900
rect 28264 25916 28316 25968
rect 28908 25916 28960 25968
rect 29644 25916 29696 25968
rect 31300 25984 31352 26036
rect 31392 25984 31444 26036
rect 31760 26027 31812 26036
rect 31760 25993 31769 26027
rect 31769 25993 31803 26027
rect 31803 25993 31812 26027
rect 31760 25984 31812 25993
rect 27436 25848 27488 25900
rect 28356 25848 28408 25900
rect 29000 25891 29052 25900
rect 29000 25857 29009 25891
rect 29009 25857 29043 25891
rect 29043 25857 29052 25891
rect 29000 25848 29052 25857
rect 32404 25984 32456 26036
rect 32588 26027 32640 26036
rect 32588 25993 32597 26027
rect 32597 25993 32631 26027
rect 32631 25993 32640 26027
rect 32588 25984 32640 25993
rect 33968 26027 34020 26036
rect 33968 25993 33977 26027
rect 33977 25993 34011 26027
rect 34011 25993 34020 26027
rect 33968 25984 34020 25993
rect 32496 25959 32548 25968
rect 32496 25925 32505 25959
rect 32505 25925 32539 25959
rect 32539 25925 32548 25959
rect 32496 25916 32548 25925
rect 35348 25916 35400 25968
rect 28816 25780 28868 25832
rect 29092 25823 29144 25832
rect 29092 25789 29101 25823
rect 29101 25789 29135 25823
rect 29135 25789 29144 25823
rect 29092 25780 29144 25789
rect 30380 25780 30432 25832
rect 22744 25712 22796 25764
rect 23296 25712 23348 25764
rect 24768 25712 24820 25764
rect 23480 25687 23532 25696
rect 23480 25653 23489 25687
rect 23489 25653 23523 25687
rect 23523 25653 23532 25687
rect 23480 25644 23532 25653
rect 24032 25687 24084 25696
rect 24032 25653 24041 25687
rect 24041 25653 24075 25687
rect 24075 25653 24084 25687
rect 24032 25644 24084 25653
rect 25688 25644 25740 25696
rect 26516 25644 26568 25696
rect 32772 25823 32824 25832
rect 32772 25789 32781 25823
rect 32781 25789 32815 25823
rect 32815 25789 32824 25823
rect 32772 25780 32824 25789
rect 32956 25780 33008 25832
rect 33784 25780 33836 25832
rect 34336 25823 34388 25832
rect 34336 25789 34345 25823
rect 34345 25789 34379 25823
rect 34379 25789 34388 25823
rect 34336 25780 34388 25789
rect 34612 25823 34664 25832
rect 34612 25789 34621 25823
rect 34621 25789 34655 25823
rect 34655 25789 34664 25823
rect 34612 25780 34664 25789
rect 31760 25644 31812 25696
rect 32496 25644 32548 25696
rect 33508 25687 33560 25696
rect 33508 25653 33517 25687
rect 33517 25653 33551 25687
rect 33551 25653 33560 25687
rect 33508 25644 33560 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5632 25440 5684 25492
rect 6000 25440 6052 25492
rect 7932 25440 7984 25492
rect 9772 25440 9824 25492
rect 10416 25440 10468 25492
rect 7656 25372 7708 25424
rect 7748 25347 7800 25356
rect 7748 25313 7757 25347
rect 7757 25313 7791 25347
rect 7791 25313 7800 25347
rect 7748 25304 7800 25313
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 1952 25211 2004 25220
rect 1952 25177 1961 25211
rect 1961 25177 1995 25211
rect 1995 25177 2004 25211
rect 1952 25168 2004 25177
rect 4068 25168 4120 25220
rect 2780 25100 2832 25152
rect 6644 25236 6696 25288
rect 8024 25372 8076 25424
rect 9680 25372 9732 25424
rect 13268 25440 13320 25492
rect 15384 25440 15436 25492
rect 10048 25304 10100 25356
rect 9404 25279 9456 25288
rect 9404 25245 9413 25279
rect 9413 25245 9447 25279
rect 9447 25245 9456 25279
rect 9404 25236 9456 25245
rect 11060 25236 11112 25288
rect 11336 25236 11388 25288
rect 15108 25372 15160 25424
rect 17040 25372 17092 25424
rect 12164 25347 12216 25356
rect 12164 25313 12173 25347
rect 12173 25313 12207 25347
rect 12207 25313 12216 25347
rect 12164 25304 12216 25313
rect 12900 25304 12952 25356
rect 13360 25304 13412 25356
rect 13728 25347 13780 25356
rect 13728 25313 13737 25347
rect 13737 25313 13771 25347
rect 13771 25313 13780 25347
rect 13728 25304 13780 25313
rect 18604 25304 18656 25356
rect 14096 25236 14148 25288
rect 14188 25279 14240 25288
rect 14188 25245 14197 25279
rect 14197 25245 14231 25279
rect 14231 25245 14240 25279
rect 14188 25236 14240 25245
rect 14648 25279 14700 25288
rect 14648 25245 14657 25279
rect 14657 25245 14691 25279
rect 14691 25245 14700 25279
rect 14648 25236 14700 25245
rect 16672 25236 16724 25288
rect 18144 25236 18196 25288
rect 18696 25236 18748 25288
rect 16764 25168 16816 25220
rect 19708 25236 19760 25288
rect 7656 25143 7708 25152
rect 7656 25109 7665 25143
rect 7665 25109 7699 25143
rect 7699 25109 7708 25143
rect 7656 25100 7708 25109
rect 7840 25100 7892 25152
rect 8392 25143 8444 25152
rect 8392 25109 8401 25143
rect 8401 25109 8435 25143
rect 8435 25109 8444 25143
rect 8392 25100 8444 25109
rect 12072 25143 12124 25152
rect 12072 25109 12081 25143
rect 12081 25109 12115 25143
rect 12115 25109 12124 25143
rect 12072 25100 12124 25109
rect 12716 25100 12768 25152
rect 13084 25100 13136 25152
rect 17224 25100 17276 25152
rect 18236 25143 18288 25152
rect 18236 25109 18245 25143
rect 18245 25109 18279 25143
rect 18279 25109 18288 25143
rect 18236 25100 18288 25109
rect 19156 25168 19208 25220
rect 20168 25440 20220 25492
rect 20352 25483 20404 25492
rect 20352 25449 20361 25483
rect 20361 25449 20395 25483
rect 20395 25449 20404 25483
rect 20352 25440 20404 25449
rect 20720 25440 20772 25492
rect 21732 25440 21784 25492
rect 22284 25372 22336 25424
rect 22560 25372 22612 25424
rect 22744 25440 22796 25492
rect 24032 25440 24084 25492
rect 24676 25440 24728 25492
rect 25320 25483 25372 25492
rect 25320 25449 25329 25483
rect 25329 25449 25363 25483
rect 25363 25449 25372 25483
rect 25320 25440 25372 25449
rect 26148 25440 26200 25492
rect 26884 25440 26936 25492
rect 29000 25440 29052 25492
rect 33508 25440 33560 25492
rect 34612 25440 34664 25492
rect 20444 25304 20496 25356
rect 19984 25100 20036 25152
rect 20720 25236 20772 25288
rect 22928 25304 22980 25356
rect 23112 25304 23164 25356
rect 22192 25236 22244 25288
rect 22376 25236 22428 25288
rect 23848 25304 23900 25356
rect 23296 25236 23348 25288
rect 24584 25304 24636 25356
rect 24676 25304 24728 25356
rect 21548 25211 21600 25220
rect 21548 25177 21557 25211
rect 21557 25177 21591 25211
rect 21591 25177 21600 25211
rect 21548 25168 21600 25177
rect 20628 25100 20680 25152
rect 24952 25168 25004 25220
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 26884 25304 26936 25356
rect 32956 25372 33008 25424
rect 25412 25168 25464 25220
rect 22928 25100 22980 25152
rect 25504 25100 25556 25152
rect 26516 25279 26568 25288
rect 26516 25245 26525 25279
rect 26525 25245 26559 25279
rect 26559 25245 26568 25279
rect 26516 25236 26568 25245
rect 26608 25279 26660 25288
rect 26608 25245 26617 25279
rect 26617 25245 26651 25279
rect 26651 25245 26660 25279
rect 26608 25236 26660 25245
rect 26700 25236 26752 25288
rect 30196 25236 30248 25288
rect 30380 25236 30432 25288
rect 32036 25236 32088 25288
rect 32496 25236 32548 25288
rect 28540 25100 28592 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 1952 24896 2004 24948
rect 7656 24896 7708 24948
rect 1676 24828 1728 24880
rect 1492 24803 1544 24812
rect 1492 24769 1501 24803
rect 1501 24769 1535 24803
rect 1535 24769 1544 24803
rect 1492 24760 1544 24769
rect 2780 24871 2832 24880
rect 2780 24837 2789 24871
rect 2789 24837 2823 24871
rect 2823 24837 2832 24871
rect 2780 24828 2832 24837
rect 6644 24828 6696 24880
rect 8392 24828 8444 24880
rect 8668 24828 8720 24880
rect 9680 24896 9732 24948
rect 10048 24896 10100 24948
rect 12256 24896 12308 24948
rect 15936 24896 15988 24948
rect 18420 24896 18472 24948
rect 20812 24896 20864 24948
rect 22468 24896 22520 24948
rect 2872 24735 2924 24744
rect 2872 24701 2881 24735
rect 2881 24701 2915 24735
rect 2915 24701 2924 24735
rect 2872 24692 2924 24701
rect 3148 24692 3200 24744
rect 3700 24735 3752 24744
rect 3700 24701 3709 24735
rect 3709 24701 3743 24735
rect 3743 24701 3752 24735
rect 3700 24692 3752 24701
rect 4068 24692 4120 24744
rect 6184 24760 6236 24812
rect 11704 24760 11756 24812
rect 12532 24760 12584 24812
rect 5448 24692 5500 24744
rect 7840 24735 7892 24744
rect 7840 24701 7849 24735
rect 7849 24701 7883 24735
rect 7883 24701 7892 24735
rect 7840 24692 7892 24701
rect 9772 24692 9824 24744
rect 10232 24735 10284 24744
rect 10232 24701 10241 24735
rect 10241 24701 10275 24735
rect 10275 24701 10284 24735
rect 10232 24692 10284 24701
rect 4804 24556 4856 24608
rect 5264 24556 5316 24608
rect 10048 24556 10100 24608
rect 13544 24760 13596 24812
rect 13820 24760 13872 24812
rect 14740 24760 14792 24812
rect 16120 24803 16172 24812
rect 16120 24769 16129 24803
rect 16129 24769 16163 24803
rect 16163 24769 16172 24803
rect 16120 24760 16172 24769
rect 16304 24803 16356 24812
rect 16304 24769 16313 24803
rect 16313 24769 16347 24803
rect 16347 24769 16356 24803
rect 16304 24760 16356 24769
rect 16672 24760 16724 24812
rect 19432 24828 19484 24880
rect 20628 24871 20680 24880
rect 20628 24837 20637 24871
rect 20637 24837 20671 24871
rect 20671 24837 20680 24871
rect 20628 24828 20680 24837
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18052 24803 18104 24812
rect 18052 24769 18061 24803
rect 18061 24769 18095 24803
rect 18095 24769 18104 24803
rect 18052 24760 18104 24769
rect 18144 24760 18196 24812
rect 18420 24760 18472 24812
rect 12348 24556 12400 24608
rect 13360 24624 13412 24676
rect 14096 24692 14148 24744
rect 14188 24735 14240 24744
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 17132 24692 17184 24744
rect 13268 24556 13320 24608
rect 13636 24556 13688 24608
rect 16028 24624 16080 24676
rect 18696 24692 18748 24744
rect 16488 24599 16540 24608
rect 16488 24565 16497 24599
rect 16497 24565 16531 24599
rect 16531 24565 16540 24599
rect 16488 24556 16540 24565
rect 18328 24624 18380 24676
rect 20168 24760 20220 24812
rect 20536 24803 20588 24812
rect 20536 24769 20543 24803
rect 20543 24769 20588 24803
rect 20536 24760 20588 24769
rect 20904 24760 20956 24812
rect 21272 24760 21324 24812
rect 22100 24803 22152 24812
rect 22100 24769 22109 24803
rect 22109 24769 22143 24803
rect 22143 24769 22152 24803
rect 22100 24760 22152 24769
rect 24584 24828 24636 24880
rect 25780 24896 25832 24948
rect 27988 24896 28040 24948
rect 28356 24896 28408 24948
rect 30656 24896 30708 24948
rect 33876 24896 33928 24948
rect 26700 24828 26752 24880
rect 27436 24828 27488 24880
rect 31760 24828 31812 24880
rect 32496 24828 32548 24880
rect 22284 24760 22336 24812
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 20996 24692 21048 24744
rect 19064 24624 19116 24676
rect 24216 24760 24268 24812
rect 24952 24760 25004 24812
rect 25504 24803 25556 24812
rect 25504 24769 25513 24803
rect 25513 24769 25547 24803
rect 25547 24769 25556 24803
rect 25504 24760 25556 24769
rect 26056 24760 26108 24812
rect 27528 24760 27580 24812
rect 28264 24760 28316 24812
rect 28632 24803 28684 24812
rect 28632 24769 28641 24803
rect 28641 24769 28675 24803
rect 28675 24769 28684 24803
rect 28632 24760 28684 24769
rect 26516 24692 26568 24744
rect 26700 24692 26752 24744
rect 28908 24692 28960 24744
rect 29920 24760 29972 24812
rect 32128 24803 32180 24812
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 32312 24803 32364 24812
rect 32312 24769 32321 24803
rect 32321 24769 32355 24803
rect 32355 24769 32364 24803
rect 32312 24760 32364 24769
rect 32404 24803 32456 24812
rect 32404 24769 32413 24803
rect 32413 24769 32447 24803
rect 32447 24769 32456 24803
rect 32404 24760 32456 24769
rect 26608 24624 26660 24676
rect 30472 24624 30524 24676
rect 32036 24624 32088 24676
rect 21088 24556 21140 24608
rect 22192 24556 22244 24608
rect 30656 24556 30708 24608
rect 32220 24599 32272 24608
rect 32220 24565 32229 24599
rect 32229 24565 32263 24599
rect 32263 24565 32272 24599
rect 32220 24556 32272 24565
rect 32588 24624 32640 24676
rect 32864 24803 32916 24812
rect 32864 24769 32873 24803
rect 32873 24769 32907 24803
rect 32907 24769 32916 24803
rect 32864 24760 32916 24769
rect 32956 24760 33008 24812
rect 35348 24556 35400 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3700 24352 3752 24404
rect 8668 24352 8720 24404
rect 12072 24352 12124 24404
rect 12532 24352 12584 24404
rect 3148 24080 3200 24132
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 5448 24216 5500 24268
rect 8300 24216 8352 24268
rect 12716 24284 12768 24336
rect 13636 24327 13688 24336
rect 13636 24293 13645 24327
rect 13645 24293 13679 24327
rect 13679 24293 13688 24327
rect 13636 24284 13688 24293
rect 14648 24352 14700 24404
rect 16304 24352 16356 24404
rect 14740 24284 14792 24336
rect 15476 24284 15528 24336
rect 17868 24395 17920 24404
rect 17868 24361 17877 24395
rect 17877 24361 17911 24395
rect 17911 24361 17920 24395
rect 17868 24352 17920 24361
rect 18328 24352 18380 24404
rect 11428 24216 11480 24268
rect 4896 24055 4948 24064
rect 4896 24021 4905 24055
rect 4905 24021 4939 24055
rect 4939 24021 4948 24055
rect 4896 24012 4948 24021
rect 6736 24123 6788 24132
rect 6736 24089 6745 24123
rect 6745 24089 6779 24123
rect 6779 24089 6788 24123
rect 6736 24080 6788 24089
rect 12716 24191 12768 24200
rect 12716 24157 12725 24191
rect 12725 24157 12759 24191
rect 12759 24157 12768 24191
rect 12716 24148 12768 24157
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 14096 24259 14148 24268
rect 14096 24225 14105 24259
rect 14105 24225 14139 24259
rect 14139 24225 14148 24259
rect 14096 24216 14148 24225
rect 15108 24216 15160 24268
rect 13820 24148 13872 24200
rect 14188 24148 14240 24200
rect 13728 24080 13780 24132
rect 14004 24080 14056 24132
rect 15292 24191 15344 24200
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 15384 24148 15436 24200
rect 15752 24191 15804 24200
rect 15752 24157 15761 24191
rect 15761 24157 15795 24191
rect 15795 24157 15804 24191
rect 15752 24148 15804 24157
rect 16028 24191 16080 24200
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 16304 24216 16356 24268
rect 16948 24216 17000 24268
rect 16396 24148 16448 24200
rect 18052 24148 18104 24200
rect 18604 24284 18656 24336
rect 19984 24352 20036 24404
rect 20260 24284 20312 24336
rect 19064 24216 19116 24268
rect 20536 24216 20588 24268
rect 20996 24352 21048 24404
rect 21272 24352 21324 24404
rect 22100 24352 22152 24404
rect 22652 24352 22704 24404
rect 24400 24352 24452 24404
rect 22008 24216 22060 24268
rect 17316 24080 17368 24132
rect 19432 24148 19484 24200
rect 19984 24191 20036 24200
rect 19984 24157 19993 24191
rect 19993 24157 20027 24191
rect 20027 24157 20036 24191
rect 19984 24148 20036 24157
rect 20444 24191 20496 24200
rect 20444 24157 20451 24191
rect 20451 24157 20496 24191
rect 20444 24148 20496 24157
rect 6920 24012 6972 24064
rect 7564 24012 7616 24064
rect 10140 24012 10192 24064
rect 11244 24012 11296 24064
rect 12072 24012 12124 24064
rect 12256 24012 12308 24064
rect 15844 24012 15896 24064
rect 16856 24012 16908 24064
rect 19340 24080 19392 24132
rect 18420 24012 18472 24064
rect 19248 24012 19300 24064
rect 22100 24148 22152 24200
rect 22560 24148 22612 24200
rect 22744 24191 22796 24200
rect 22744 24157 22753 24191
rect 22753 24157 22787 24191
rect 22787 24157 22796 24191
rect 22744 24148 22796 24157
rect 23388 24284 23440 24336
rect 24860 24284 24912 24336
rect 25504 24352 25556 24404
rect 26700 24352 26752 24404
rect 28632 24352 28684 24404
rect 28724 24352 28776 24404
rect 30564 24352 30616 24404
rect 25596 24216 25648 24268
rect 23112 24148 23164 24200
rect 24768 24148 24820 24200
rect 25688 24148 25740 24200
rect 26884 24216 26936 24268
rect 28908 24284 28960 24336
rect 29184 24284 29236 24336
rect 26608 24148 26660 24200
rect 26792 24148 26844 24200
rect 27344 24148 27396 24200
rect 27804 24148 27856 24200
rect 28816 24259 28868 24268
rect 28816 24225 28825 24259
rect 28825 24225 28859 24259
rect 28859 24225 28868 24259
rect 28816 24216 28868 24225
rect 30196 24148 30248 24200
rect 30380 24191 30432 24200
rect 30380 24157 30389 24191
rect 30389 24157 30423 24191
rect 30423 24157 30432 24191
rect 30380 24148 30432 24157
rect 31024 24284 31076 24336
rect 32864 24352 32916 24404
rect 32128 24284 32180 24336
rect 32496 24327 32548 24336
rect 32496 24293 32505 24327
rect 32505 24293 32539 24327
rect 32539 24293 32548 24327
rect 32496 24284 32548 24293
rect 30656 24191 30708 24200
rect 30656 24157 30665 24191
rect 30665 24157 30699 24191
rect 30699 24157 30708 24191
rect 30656 24148 30708 24157
rect 20168 24012 20220 24064
rect 21640 24080 21692 24132
rect 22008 24080 22060 24132
rect 23756 24080 23808 24132
rect 20628 24012 20680 24064
rect 20904 24055 20956 24064
rect 20904 24021 20913 24055
rect 20913 24021 20947 24055
rect 20947 24021 20956 24055
rect 20904 24012 20956 24021
rect 21272 24055 21324 24064
rect 21272 24021 21281 24055
rect 21281 24021 21315 24055
rect 21315 24021 21324 24055
rect 21272 24012 21324 24021
rect 21364 24055 21416 24064
rect 21364 24021 21373 24055
rect 21373 24021 21407 24055
rect 21407 24021 21416 24055
rect 21364 24012 21416 24021
rect 22192 24012 22244 24064
rect 22744 24012 22796 24064
rect 23388 24012 23440 24064
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 24768 24012 24820 24064
rect 24952 24055 25004 24064
rect 24952 24021 24961 24055
rect 24961 24021 24995 24055
rect 24995 24021 25004 24055
rect 26516 24080 26568 24132
rect 26976 24123 27028 24132
rect 26976 24089 26985 24123
rect 26985 24089 27019 24123
rect 27019 24089 27028 24123
rect 26976 24080 27028 24089
rect 30840 24148 30892 24200
rect 31484 24216 31536 24268
rect 32036 24191 32088 24200
rect 32036 24157 32045 24191
rect 32045 24157 32079 24191
rect 32079 24157 32088 24191
rect 32036 24148 32088 24157
rect 32128 24191 32180 24200
rect 32128 24157 32137 24191
rect 32137 24157 32171 24191
rect 32171 24157 32180 24191
rect 32128 24148 32180 24157
rect 32404 24191 32456 24200
rect 32404 24157 32413 24191
rect 32413 24157 32447 24191
rect 32447 24157 32456 24191
rect 32404 24148 32456 24157
rect 32588 24148 32640 24200
rect 32956 24148 33008 24200
rect 33876 24148 33928 24200
rect 33968 24191 34020 24200
rect 33968 24157 33977 24191
rect 33977 24157 34011 24191
rect 34011 24157 34020 24191
rect 33968 24148 34020 24157
rect 34244 24216 34296 24268
rect 24952 24012 25004 24021
rect 26240 24012 26292 24064
rect 27620 24012 27672 24064
rect 28540 24012 28592 24064
rect 30748 24012 30800 24064
rect 30840 24055 30892 24064
rect 30840 24021 30849 24055
rect 30849 24021 30883 24055
rect 30883 24021 30892 24055
rect 30840 24012 30892 24021
rect 31208 24055 31260 24064
rect 31208 24021 31217 24055
rect 31217 24021 31251 24055
rect 31251 24021 31260 24055
rect 31208 24012 31260 24021
rect 31852 24055 31904 24064
rect 31852 24021 31861 24055
rect 31861 24021 31895 24055
rect 31895 24021 31904 24055
rect 31852 24012 31904 24021
rect 32220 24012 32272 24064
rect 35072 24080 35124 24132
rect 32956 24055 33008 24064
rect 32956 24021 32965 24055
rect 32965 24021 32999 24055
rect 32999 24021 33008 24055
rect 32956 24012 33008 24021
rect 34520 24055 34572 24064
rect 34520 24021 34529 24055
rect 34529 24021 34563 24055
rect 34563 24021 34572 24055
rect 34520 24012 34572 24021
rect 34704 24012 34756 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 6736 23808 6788 23860
rect 1676 23740 1728 23792
rect 4068 23740 4120 23792
rect 10324 23808 10376 23860
rect 12716 23808 12768 23860
rect 1768 23604 1820 23656
rect 6920 23604 6972 23656
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 7656 23604 7708 23613
rect 11612 23740 11664 23792
rect 10784 23672 10836 23724
rect 11428 23672 11480 23724
rect 11520 23604 11572 23656
rect 13360 23808 13412 23860
rect 13912 23808 13964 23860
rect 14464 23808 14516 23860
rect 13268 23783 13320 23792
rect 13268 23749 13277 23783
rect 13277 23749 13311 23783
rect 13311 23749 13320 23783
rect 13268 23740 13320 23749
rect 13544 23740 13596 23792
rect 13360 23672 13412 23724
rect 13728 23715 13780 23724
rect 13728 23681 13737 23715
rect 13737 23681 13771 23715
rect 13771 23681 13780 23715
rect 13728 23672 13780 23681
rect 15292 23740 15344 23792
rect 15936 23740 15988 23792
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 14280 23672 14332 23724
rect 15200 23672 15252 23724
rect 15844 23715 15896 23724
rect 15844 23681 15853 23715
rect 15853 23681 15887 23715
rect 15887 23681 15896 23715
rect 15844 23672 15896 23681
rect 18328 23808 18380 23860
rect 18512 23808 18564 23860
rect 22100 23808 22152 23860
rect 22192 23808 22244 23860
rect 15568 23604 15620 23656
rect 7104 23536 7156 23588
rect 13912 23536 13964 23588
rect 16120 23536 16172 23588
rect 16212 23536 16264 23588
rect 17040 23604 17092 23656
rect 17408 23672 17460 23724
rect 18420 23715 18472 23724
rect 18420 23681 18429 23715
rect 18429 23681 18463 23715
rect 18463 23681 18472 23715
rect 18420 23672 18472 23681
rect 18512 23672 18564 23724
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 19432 23740 19484 23792
rect 20352 23740 20404 23792
rect 21364 23740 21416 23792
rect 20536 23672 20588 23724
rect 20812 23672 20864 23724
rect 21456 23672 21508 23724
rect 21732 23672 21784 23724
rect 22744 23740 22796 23792
rect 23112 23740 23164 23792
rect 21824 23604 21876 23656
rect 22652 23715 22704 23724
rect 22652 23681 22662 23715
rect 22662 23681 22696 23715
rect 22696 23681 22704 23715
rect 22652 23672 22704 23681
rect 23388 23808 23440 23860
rect 17224 23536 17276 23588
rect 21272 23536 21324 23588
rect 3332 23468 3384 23520
rect 10232 23468 10284 23520
rect 13360 23468 13412 23520
rect 13636 23468 13688 23520
rect 14188 23468 14240 23520
rect 18144 23468 18196 23520
rect 18972 23468 19024 23520
rect 19248 23468 19300 23520
rect 21916 23536 21968 23588
rect 23020 23536 23072 23588
rect 23112 23536 23164 23588
rect 23572 23672 23624 23724
rect 25320 23740 25372 23792
rect 26240 23808 26292 23860
rect 28724 23808 28776 23860
rect 29184 23808 29236 23860
rect 30840 23808 30892 23860
rect 32128 23808 32180 23860
rect 32312 23808 32364 23860
rect 32404 23851 32456 23860
rect 32404 23817 32413 23851
rect 32413 23817 32447 23851
rect 32447 23817 32456 23851
rect 32404 23808 32456 23817
rect 34520 23808 34572 23860
rect 35348 23808 35400 23860
rect 26516 23740 26568 23792
rect 27988 23740 28040 23792
rect 28264 23740 28316 23792
rect 29644 23740 29696 23792
rect 24124 23672 24176 23724
rect 27068 23672 27120 23724
rect 27252 23715 27304 23724
rect 27252 23681 27261 23715
rect 27261 23681 27295 23715
rect 27295 23681 27304 23715
rect 27252 23672 27304 23681
rect 27344 23715 27396 23724
rect 27344 23681 27353 23715
rect 27353 23681 27387 23715
rect 27387 23681 27396 23715
rect 27344 23672 27396 23681
rect 23940 23604 23992 23656
rect 24584 23647 24636 23656
rect 24584 23613 24593 23647
rect 24593 23613 24627 23647
rect 24627 23613 24636 23647
rect 24584 23604 24636 23613
rect 24676 23604 24728 23656
rect 27620 23672 27672 23724
rect 31024 23740 31076 23792
rect 21640 23468 21692 23520
rect 22376 23468 22428 23520
rect 22652 23468 22704 23520
rect 31484 23604 31536 23656
rect 33968 23604 34020 23656
rect 31116 23536 31168 23588
rect 33232 23536 33284 23588
rect 35072 23647 35124 23656
rect 35072 23613 35081 23647
rect 35081 23613 35115 23647
rect 35115 23613 35124 23647
rect 35072 23604 35124 23613
rect 34796 23536 34848 23588
rect 25596 23468 25648 23520
rect 32772 23468 32824 23520
rect 34244 23468 34296 23520
rect 34612 23511 34664 23520
rect 34612 23477 34621 23511
rect 34621 23477 34655 23511
rect 34655 23477 34664 23511
rect 34612 23468 34664 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1768 23307 1820 23316
rect 1768 23273 1777 23307
rect 1777 23273 1811 23307
rect 1811 23273 1820 23307
rect 1768 23264 1820 23273
rect 2872 23264 2924 23316
rect 3148 23128 3200 23180
rect 3332 23060 3384 23112
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 7656 23264 7708 23316
rect 8116 23264 8168 23316
rect 4804 23171 4856 23180
rect 4804 23137 4813 23171
rect 4813 23137 4847 23171
rect 4847 23137 4856 23171
rect 4804 23128 4856 23137
rect 5448 23128 5500 23180
rect 5632 23128 5684 23180
rect 6368 23196 6420 23248
rect 7288 23196 7340 23248
rect 6920 23128 6972 23180
rect 4160 23060 4212 23069
rect 4620 23060 4672 23112
rect 6184 23060 6236 23112
rect 9404 23196 9456 23248
rect 11336 23196 11388 23248
rect 13728 23196 13780 23248
rect 13820 23239 13872 23248
rect 13820 23205 13829 23239
rect 13829 23205 13863 23239
rect 13863 23205 13872 23239
rect 13820 23196 13872 23205
rect 14188 23264 14240 23316
rect 16948 23264 17000 23316
rect 3608 22992 3660 23044
rect 4344 22992 4396 23044
rect 4988 22992 5040 23044
rect 5080 23035 5132 23044
rect 5080 23001 5089 23035
rect 5089 23001 5123 23035
rect 5123 23001 5132 23035
rect 5080 22992 5132 23001
rect 7012 23035 7064 23044
rect 2780 22967 2832 22976
rect 2780 22933 2789 22967
rect 2789 22933 2823 22967
rect 2823 22933 2832 22967
rect 2780 22924 2832 22933
rect 7012 23001 7021 23035
rect 7021 23001 7055 23035
rect 7055 23001 7064 23035
rect 7012 22992 7064 23001
rect 6644 22967 6696 22976
rect 6644 22933 6653 22967
rect 6653 22933 6687 22967
rect 6687 22933 6696 22967
rect 6644 22924 6696 22933
rect 6736 22924 6788 22976
rect 8484 23103 8536 23112
rect 8484 23069 8519 23103
rect 8519 23069 8536 23103
rect 8484 23060 8536 23069
rect 8668 23103 8720 23112
rect 8668 23069 8677 23103
rect 8677 23069 8711 23103
rect 8711 23069 8720 23103
rect 8668 23060 8720 23069
rect 10232 23128 10284 23180
rect 13452 23128 13504 23180
rect 12900 23060 12952 23112
rect 15108 23128 15160 23180
rect 16028 23196 16080 23248
rect 16304 23239 16356 23248
rect 16304 23205 16313 23239
rect 16313 23205 16347 23239
rect 16347 23205 16356 23239
rect 16304 23196 16356 23205
rect 17592 23196 17644 23248
rect 16672 23128 16724 23180
rect 17040 23171 17092 23180
rect 17040 23137 17049 23171
rect 17049 23137 17083 23171
rect 17083 23137 17092 23171
rect 17040 23128 17092 23137
rect 18604 23264 18656 23316
rect 20628 23264 20680 23316
rect 21640 23264 21692 23316
rect 17776 23196 17828 23248
rect 21364 23196 21416 23248
rect 18880 23128 18932 23180
rect 21180 23128 21232 23180
rect 21640 23128 21692 23180
rect 8300 23035 8352 23044
rect 8300 23001 8309 23035
rect 8309 23001 8343 23035
rect 8343 23001 8352 23035
rect 8300 22992 8352 23001
rect 8944 23035 8996 23044
rect 8944 23001 8953 23035
rect 8953 23001 8987 23035
rect 8987 23001 8996 23035
rect 8944 22992 8996 23001
rect 9128 23035 9180 23044
rect 9128 23001 9137 23035
rect 9137 23001 9171 23035
rect 9171 23001 9180 23035
rect 9128 22992 9180 23001
rect 11888 23035 11940 23044
rect 11888 23001 11897 23035
rect 11897 23001 11931 23035
rect 11931 23001 11940 23035
rect 13728 23060 13780 23112
rect 14188 23060 14240 23112
rect 15292 23060 15344 23112
rect 16212 23103 16264 23112
rect 16212 23069 16221 23103
rect 16221 23069 16255 23103
rect 16255 23069 16264 23103
rect 16212 23060 16264 23069
rect 16396 23060 16448 23112
rect 17408 23060 17460 23112
rect 18512 23060 18564 23112
rect 18604 23103 18656 23112
rect 18604 23069 18613 23103
rect 18613 23069 18647 23103
rect 18647 23069 18656 23103
rect 18604 23060 18656 23069
rect 11888 22992 11940 23001
rect 16948 22992 17000 23044
rect 17500 23035 17552 23044
rect 17500 23001 17509 23035
rect 17509 23001 17543 23035
rect 17543 23001 17552 23035
rect 17500 22992 17552 23001
rect 19064 23060 19116 23112
rect 20720 23060 20772 23112
rect 18972 22992 19024 23044
rect 15016 22924 15068 22976
rect 15108 22924 15160 22976
rect 18604 22924 18656 22976
rect 18880 22924 18932 22976
rect 19892 22992 19944 23044
rect 20076 22992 20128 23044
rect 20260 22992 20312 23044
rect 20536 22992 20588 23044
rect 22928 23264 22980 23316
rect 24584 23264 24636 23316
rect 28816 23264 28868 23316
rect 33876 23264 33928 23316
rect 35624 23264 35676 23316
rect 22192 23171 22244 23180
rect 22192 23137 22201 23171
rect 22201 23137 22235 23171
rect 22235 23137 22244 23171
rect 22192 23128 22244 23137
rect 21916 23060 21968 23112
rect 22100 23103 22152 23112
rect 22100 23069 22109 23103
rect 22109 23069 22143 23103
rect 22143 23069 22152 23103
rect 22100 23060 22152 23069
rect 22376 23128 22428 23180
rect 22652 23128 22704 23180
rect 34244 23196 34296 23248
rect 24492 23128 24544 23180
rect 25320 23128 25372 23180
rect 22560 23060 22612 23112
rect 22744 23060 22796 23112
rect 23112 23060 23164 23112
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 25228 23103 25280 23112
rect 25228 23069 25237 23103
rect 25237 23069 25271 23103
rect 25271 23069 25280 23103
rect 25228 23060 25280 23069
rect 26516 23128 26568 23180
rect 27252 23128 27304 23180
rect 25596 23103 25648 23112
rect 25596 23069 25610 23103
rect 25610 23069 25644 23103
rect 25644 23069 25648 23103
rect 25596 23060 25648 23069
rect 26608 23060 26660 23112
rect 25504 23035 25556 23044
rect 25504 23001 25513 23035
rect 25513 23001 25547 23035
rect 25547 23001 25556 23035
rect 25504 22992 25556 23001
rect 27068 23035 27120 23044
rect 27068 23001 27077 23035
rect 27077 23001 27111 23035
rect 27111 23001 27120 23035
rect 27068 22992 27120 23001
rect 31208 23060 31260 23112
rect 32128 23060 32180 23112
rect 33968 23060 34020 23112
rect 35624 23060 35676 23112
rect 37280 23060 37332 23112
rect 35808 22992 35860 23044
rect 20996 22924 21048 22976
rect 22100 22924 22152 22976
rect 22376 22924 22428 22976
rect 22560 22924 22612 22976
rect 23664 22924 23716 22976
rect 24400 22924 24452 22976
rect 30932 22924 30984 22976
rect 32312 22924 32364 22976
rect 33600 22924 33652 22976
rect 35348 22967 35400 22976
rect 35348 22933 35357 22967
rect 35357 22933 35391 22967
rect 35391 22933 35400 22967
rect 35348 22924 35400 22933
rect 35900 22967 35952 22976
rect 35900 22933 35909 22967
rect 35909 22933 35943 22967
rect 35943 22933 35952 22967
rect 35900 22924 35952 22933
rect 37372 22967 37424 22976
rect 37372 22933 37381 22967
rect 37381 22933 37415 22967
rect 37415 22933 37424 22967
rect 37372 22924 37424 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1492 22720 1544 22772
rect 2688 22720 2740 22772
rect 2780 22720 2832 22772
rect 3608 22720 3660 22772
rect 3976 22720 4028 22772
rect 5080 22720 5132 22772
rect 2504 22627 2556 22636
rect 2504 22593 2513 22627
rect 2513 22593 2547 22627
rect 2547 22593 2556 22627
rect 2504 22584 2556 22593
rect 2596 22627 2648 22636
rect 2596 22593 2605 22627
rect 2605 22593 2639 22627
rect 2639 22593 2648 22627
rect 2596 22584 2648 22593
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2780 22584 2832 22593
rect 3700 22695 3752 22704
rect 3700 22661 3709 22695
rect 3709 22661 3743 22695
rect 3743 22661 3752 22695
rect 3700 22652 3752 22661
rect 4160 22652 4212 22704
rect 4252 22695 4304 22704
rect 4252 22661 4261 22695
rect 4261 22661 4295 22695
rect 4295 22661 4304 22695
rect 4252 22652 4304 22661
rect 3056 22627 3108 22636
rect 3056 22593 3065 22627
rect 3065 22593 3099 22627
rect 3099 22593 3108 22627
rect 3056 22584 3108 22593
rect 3516 22627 3568 22636
rect 3516 22593 3525 22627
rect 3525 22593 3559 22627
rect 3559 22593 3568 22627
rect 3516 22584 3568 22593
rect 3976 22627 4028 22636
rect 3976 22593 3985 22627
rect 3985 22593 4019 22627
rect 4019 22593 4028 22627
rect 3976 22584 4028 22593
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 4620 22584 4672 22636
rect 6644 22720 6696 22772
rect 7196 22720 7248 22772
rect 4344 22516 4396 22568
rect 3240 22380 3292 22432
rect 4252 22380 4304 22432
rect 4804 22380 4856 22432
rect 6736 22584 6788 22636
rect 6920 22627 6972 22636
rect 6920 22593 6929 22627
rect 6929 22593 6963 22627
rect 6963 22593 6972 22627
rect 6920 22584 6972 22593
rect 7104 22627 7156 22636
rect 7104 22593 7139 22627
rect 7139 22593 7156 22627
rect 7104 22584 7156 22593
rect 7656 22720 7708 22772
rect 8300 22763 8352 22772
rect 8300 22729 8309 22763
rect 8309 22729 8343 22763
rect 8343 22729 8352 22763
rect 8300 22720 8352 22729
rect 9864 22720 9916 22772
rect 11520 22763 11572 22772
rect 11520 22729 11529 22763
rect 11529 22729 11563 22763
rect 11563 22729 11572 22763
rect 11520 22720 11572 22729
rect 11888 22763 11940 22772
rect 11888 22729 11897 22763
rect 11897 22729 11931 22763
rect 11931 22729 11940 22763
rect 11888 22720 11940 22729
rect 11980 22720 12032 22772
rect 7380 22652 7432 22704
rect 7472 22584 7524 22636
rect 8116 22652 8168 22704
rect 8944 22652 8996 22704
rect 10968 22652 11020 22704
rect 7196 22380 7248 22432
rect 7288 22380 7340 22432
rect 7564 22380 7616 22432
rect 15016 22720 15068 22772
rect 21088 22720 21140 22772
rect 21456 22720 21508 22772
rect 21916 22720 21968 22772
rect 12440 22584 12492 22636
rect 14280 22627 14332 22636
rect 14280 22593 14289 22627
rect 14289 22593 14323 22627
rect 14323 22593 14332 22627
rect 14280 22584 14332 22593
rect 14740 22584 14792 22636
rect 10784 22516 10836 22568
rect 11980 22559 12032 22568
rect 11980 22525 11989 22559
rect 11989 22525 12023 22559
rect 12023 22525 12032 22559
rect 11980 22516 12032 22525
rect 12164 22559 12216 22568
rect 12164 22525 12173 22559
rect 12173 22525 12207 22559
rect 12207 22525 12216 22559
rect 12164 22516 12216 22525
rect 15752 22652 15804 22704
rect 15016 22627 15068 22636
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 15384 22584 15436 22636
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 15844 22584 15896 22636
rect 18144 22652 18196 22704
rect 17316 22627 17368 22636
rect 17316 22593 17325 22627
rect 17325 22593 17359 22627
rect 17359 22593 17368 22627
rect 17316 22584 17368 22593
rect 17684 22627 17736 22636
rect 17684 22593 17693 22627
rect 17693 22593 17727 22627
rect 17727 22593 17736 22627
rect 17684 22584 17736 22593
rect 11428 22448 11480 22500
rect 13176 22448 13228 22500
rect 13728 22448 13780 22500
rect 8392 22380 8444 22432
rect 8484 22380 8536 22432
rect 8668 22380 8720 22432
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 15200 22491 15252 22500
rect 15200 22457 15209 22491
rect 15209 22457 15243 22491
rect 15243 22457 15252 22491
rect 15200 22448 15252 22457
rect 16856 22559 16908 22568
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 17132 22559 17184 22568
rect 17132 22525 17141 22559
rect 17141 22525 17175 22559
rect 17175 22525 17184 22559
rect 17132 22516 17184 22525
rect 17592 22559 17644 22568
rect 16488 22448 16540 22500
rect 17592 22525 17601 22559
rect 17601 22525 17635 22559
rect 17635 22525 17644 22559
rect 17592 22516 17644 22525
rect 21824 22652 21876 22704
rect 22744 22720 22796 22772
rect 27252 22720 27304 22772
rect 31208 22720 31260 22772
rect 18328 22584 18380 22636
rect 18972 22627 19024 22636
rect 18972 22593 18981 22627
rect 18981 22593 19015 22627
rect 19015 22593 19024 22627
rect 18972 22584 19024 22593
rect 19064 22627 19116 22636
rect 19064 22593 19073 22627
rect 19073 22593 19107 22627
rect 19107 22593 19116 22627
rect 19064 22584 19116 22593
rect 19248 22584 19300 22636
rect 20444 22627 20496 22636
rect 20444 22593 20453 22627
rect 20453 22593 20487 22627
rect 20487 22593 20496 22627
rect 20444 22584 20496 22593
rect 20628 22584 20680 22636
rect 18880 22516 18932 22568
rect 20536 22448 20588 22500
rect 20904 22584 20956 22636
rect 21180 22627 21232 22636
rect 21180 22593 21189 22627
rect 21189 22593 21223 22627
rect 21223 22593 21232 22627
rect 21180 22584 21232 22593
rect 22468 22584 22520 22636
rect 25596 22584 25648 22636
rect 26332 22584 26384 22636
rect 26976 22627 27028 22636
rect 26976 22593 26985 22627
rect 26985 22593 27019 22627
rect 27019 22593 27028 22627
rect 26976 22584 27028 22593
rect 27252 22627 27304 22636
rect 27252 22593 27261 22627
rect 27261 22593 27295 22627
rect 27295 22593 27304 22627
rect 27252 22584 27304 22593
rect 27344 22627 27396 22636
rect 27344 22593 27353 22627
rect 27353 22593 27387 22627
rect 27387 22593 27396 22627
rect 27344 22584 27396 22593
rect 27620 22584 27672 22636
rect 27712 22584 27764 22636
rect 28724 22627 28776 22636
rect 28724 22593 28733 22627
rect 28733 22593 28767 22627
rect 28767 22593 28776 22627
rect 28724 22584 28776 22593
rect 21180 22448 21232 22500
rect 21456 22516 21508 22568
rect 22376 22516 22428 22568
rect 23112 22516 23164 22568
rect 28816 22516 28868 22568
rect 29460 22627 29512 22636
rect 29460 22593 29469 22627
rect 29469 22593 29503 22627
rect 29503 22593 29512 22627
rect 29460 22584 29512 22593
rect 32128 22652 32180 22704
rect 30012 22516 30064 22568
rect 22744 22448 22796 22500
rect 19340 22380 19392 22432
rect 20352 22423 20404 22432
rect 20352 22389 20361 22423
rect 20361 22389 20395 22423
rect 20395 22389 20404 22423
rect 20352 22380 20404 22389
rect 20812 22423 20864 22432
rect 20812 22389 20821 22423
rect 20821 22389 20855 22423
rect 20855 22389 20864 22423
rect 20812 22380 20864 22389
rect 21364 22380 21416 22432
rect 21732 22380 21784 22432
rect 21824 22423 21876 22432
rect 21824 22389 21833 22423
rect 21833 22389 21867 22423
rect 21867 22389 21876 22423
rect 21824 22380 21876 22389
rect 22284 22380 22336 22432
rect 31024 22448 31076 22500
rect 31760 22516 31812 22568
rect 32312 22720 32364 22772
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 32956 22584 33008 22636
rect 34152 22627 34204 22636
rect 34152 22593 34161 22627
rect 34161 22593 34195 22627
rect 34195 22593 34204 22627
rect 34152 22584 34204 22593
rect 34704 22720 34756 22772
rect 35900 22720 35952 22772
rect 37372 22720 37424 22772
rect 34796 22652 34848 22704
rect 34704 22627 34756 22636
rect 34704 22593 34713 22627
rect 34713 22593 34747 22627
rect 34747 22593 34756 22627
rect 34704 22584 34756 22593
rect 35808 22652 35860 22704
rect 33508 22448 33560 22500
rect 29092 22423 29144 22432
rect 29092 22389 29101 22423
rect 29101 22389 29135 22423
rect 29135 22389 29144 22423
rect 29092 22380 29144 22389
rect 29736 22380 29788 22432
rect 31484 22423 31536 22432
rect 31484 22389 31493 22423
rect 31493 22389 31527 22423
rect 31527 22389 31536 22423
rect 31484 22380 31536 22389
rect 32128 22423 32180 22432
rect 32128 22389 32137 22423
rect 32137 22389 32171 22423
rect 32171 22389 32180 22423
rect 32128 22380 32180 22389
rect 34244 22423 34296 22432
rect 34244 22389 34253 22423
rect 34253 22389 34287 22423
rect 34287 22389 34296 22423
rect 34244 22380 34296 22389
rect 37832 22491 37884 22500
rect 37832 22457 37841 22491
rect 37841 22457 37875 22491
rect 37875 22457 37884 22491
rect 37832 22448 37884 22457
rect 35900 22423 35952 22432
rect 35900 22389 35909 22423
rect 35909 22389 35943 22423
rect 35943 22389 35952 22423
rect 35900 22380 35952 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3516 22176 3568 22228
rect 6920 22176 6972 22228
rect 7012 22176 7064 22228
rect 7472 22176 7524 22228
rect 3332 22108 3384 22160
rect 3240 22040 3292 22092
rect 4988 22108 5040 22160
rect 4896 22040 4948 22092
rect 4804 22015 4856 22024
rect 3884 21904 3936 21956
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 4160 21836 4212 21888
rect 4528 21836 4580 21888
rect 4988 21879 5040 21888
rect 4988 21845 4997 21879
rect 4997 21845 5031 21879
rect 5031 21845 5040 21879
rect 4988 21836 5040 21845
rect 5632 22015 5684 22024
rect 5632 21981 5641 22015
rect 5641 21981 5675 22015
rect 5675 21981 5684 22015
rect 5632 21972 5684 21981
rect 6644 22108 6696 22160
rect 5908 22083 5960 22092
rect 5908 22049 5917 22083
rect 5917 22049 5951 22083
rect 5951 22049 5960 22083
rect 5908 22040 5960 22049
rect 6184 22040 6236 22092
rect 5540 21947 5592 21956
rect 5540 21913 5549 21947
rect 5549 21913 5583 21947
rect 5583 21913 5592 21947
rect 5540 21904 5592 21913
rect 6000 21947 6052 21956
rect 6000 21913 6009 21947
rect 6009 21913 6043 21947
rect 6043 21913 6052 21947
rect 6000 21904 6052 21913
rect 7196 21972 7248 22024
rect 7104 21904 7156 21956
rect 6644 21836 6696 21888
rect 11980 22176 12032 22228
rect 8300 22108 8352 22160
rect 8576 22108 8628 22160
rect 15384 22108 15436 22160
rect 8392 21972 8444 22024
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 9312 22083 9364 22092
rect 9312 22049 9321 22083
rect 9321 22049 9355 22083
rect 9355 22049 9364 22083
rect 9312 22040 9364 22049
rect 11520 22083 11572 22092
rect 11520 22049 11529 22083
rect 11529 22049 11563 22083
rect 11563 22049 11572 22083
rect 11520 22040 11572 22049
rect 12256 21972 12308 22024
rect 7748 21947 7800 21956
rect 7748 21913 7757 21947
rect 7757 21913 7791 21947
rect 7791 21913 7800 21947
rect 7748 21904 7800 21913
rect 10324 21904 10376 21956
rect 10876 21904 10928 21956
rect 11336 21879 11388 21888
rect 11336 21845 11345 21879
rect 11345 21845 11379 21879
rect 11379 21845 11388 21879
rect 11336 21836 11388 21845
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 12900 22015 12952 22024
rect 12900 21981 12909 22015
rect 12909 21981 12943 22015
rect 12943 21981 12952 22015
rect 12900 21972 12952 21981
rect 15200 21972 15252 22024
rect 14924 21836 14976 21888
rect 15844 22083 15896 22092
rect 15844 22049 15853 22083
rect 15853 22049 15887 22083
rect 15887 22049 15896 22083
rect 15844 22040 15896 22049
rect 16764 22108 16816 22160
rect 18696 22108 18748 22160
rect 20352 22176 20404 22228
rect 20812 22176 20864 22228
rect 20996 22219 21048 22228
rect 20996 22185 21005 22219
rect 21005 22185 21039 22219
rect 21039 22185 21048 22219
rect 20996 22176 21048 22185
rect 21824 22176 21876 22228
rect 25504 22176 25556 22228
rect 22192 22108 22244 22160
rect 22376 22108 22428 22160
rect 24400 22151 24452 22160
rect 24400 22117 24409 22151
rect 24409 22117 24443 22151
rect 24443 22117 24452 22151
rect 24400 22108 24452 22117
rect 24952 22108 25004 22160
rect 28356 22176 28408 22228
rect 29460 22176 29512 22228
rect 30380 22176 30432 22228
rect 31484 22176 31536 22228
rect 27620 22108 27672 22160
rect 28172 22108 28224 22160
rect 17592 22040 17644 22092
rect 16764 21972 16816 22024
rect 16856 22015 16908 22024
rect 16856 21981 16865 22015
rect 16865 21981 16899 22015
rect 16899 21981 16908 22015
rect 16856 21972 16908 21981
rect 17132 22015 17184 22024
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 18144 21972 18196 22024
rect 19064 22040 19116 22092
rect 20260 22040 20312 22092
rect 21272 21972 21324 22024
rect 23204 22040 23256 22092
rect 21456 21972 21508 22024
rect 21640 21972 21692 22024
rect 22100 21972 22152 22024
rect 22284 22015 22336 22024
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 19432 21836 19484 21888
rect 21456 21836 21508 21888
rect 22192 21836 22244 21888
rect 22376 21904 22428 21956
rect 22836 21904 22888 21956
rect 24860 22015 24912 22024
rect 24860 21981 24869 22015
rect 24869 21981 24903 22015
rect 24903 21981 24912 22015
rect 24860 21972 24912 21981
rect 24952 21972 25004 22024
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 25412 22015 25464 22024
rect 25412 21981 25421 22015
rect 25421 21981 25455 22015
rect 25455 21981 25464 22015
rect 25412 21972 25464 21981
rect 25504 22015 25556 22024
rect 25504 21981 25513 22015
rect 25513 21981 25547 22015
rect 25547 21981 25556 22015
rect 25504 21972 25556 21981
rect 26976 22040 27028 22092
rect 25320 21947 25372 21956
rect 25320 21913 25329 21947
rect 25329 21913 25363 21947
rect 25363 21913 25372 21947
rect 25320 21904 25372 21913
rect 25688 21904 25740 21956
rect 25964 21972 26016 22024
rect 27344 21972 27396 22024
rect 27988 21972 28040 22024
rect 28816 22083 28868 22092
rect 28816 22049 28825 22083
rect 28825 22049 28859 22083
rect 28859 22049 28868 22083
rect 28816 22040 28868 22049
rect 28540 22015 28592 22024
rect 28540 21981 28549 22015
rect 28549 21981 28583 22015
rect 28583 21981 28592 22015
rect 28540 21972 28592 21981
rect 28724 21972 28776 22024
rect 30656 22108 30708 22160
rect 31576 22108 31628 22160
rect 31944 22108 31996 22160
rect 26884 21904 26936 21956
rect 23756 21836 23808 21888
rect 27620 21836 27672 21888
rect 27804 21947 27856 21956
rect 27804 21913 27813 21947
rect 27813 21913 27847 21947
rect 27847 21913 27856 21947
rect 27804 21904 27856 21913
rect 28356 21947 28408 21956
rect 28356 21913 28365 21947
rect 28365 21913 28399 21947
rect 28399 21913 28408 21947
rect 28356 21904 28408 21913
rect 28448 21947 28500 21956
rect 28448 21913 28457 21947
rect 28457 21913 28491 21947
rect 28491 21913 28500 21947
rect 28448 21904 28500 21913
rect 29736 22015 29788 22024
rect 29736 21981 29745 22015
rect 29745 21981 29779 22015
rect 29779 21981 29788 22015
rect 29736 21972 29788 21981
rect 29000 21836 29052 21888
rect 29092 21836 29144 21888
rect 29920 21836 29972 21888
rect 30380 22015 30432 22024
rect 30380 21981 30389 22015
rect 30389 21981 30423 22015
rect 30423 21981 30432 22015
rect 30380 21972 30432 21981
rect 32312 22108 32364 22160
rect 32680 22108 32732 22160
rect 31208 22015 31260 22024
rect 31208 21981 31217 22015
rect 31217 21981 31251 22015
rect 31251 21981 31260 22015
rect 31208 21972 31260 21981
rect 31576 22015 31628 22024
rect 31576 21981 31585 22015
rect 31585 21981 31619 22015
rect 31619 21981 31628 22015
rect 31576 21972 31628 21981
rect 31852 22015 31904 22024
rect 31852 21981 31861 22015
rect 31861 21981 31895 22015
rect 31895 21981 31904 22015
rect 31852 21972 31904 21981
rect 32036 22015 32088 22024
rect 32036 21981 32045 22015
rect 32045 21981 32079 22015
rect 32079 21981 32088 22015
rect 32036 21972 32088 21981
rect 32128 21972 32180 22024
rect 32404 21972 32456 22024
rect 30472 21879 30524 21888
rect 30472 21845 30481 21879
rect 30481 21845 30515 21879
rect 30515 21845 30524 21879
rect 30472 21836 30524 21845
rect 31300 21836 31352 21888
rect 32864 22015 32916 22024
rect 32864 21981 32873 22015
rect 32873 21981 32907 22015
rect 32907 21981 32916 22015
rect 32864 21972 32916 21981
rect 33140 21972 33192 22024
rect 32496 21836 32548 21888
rect 32772 21836 32824 21888
rect 33508 22040 33560 22092
rect 34612 22040 34664 22092
rect 33876 21904 33928 21956
rect 34336 22015 34388 22024
rect 34336 21981 34345 22015
rect 34345 21981 34379 22015
rect 34379 21981 34388 22015
rect 34336 21972 34388 21981
rect 35440 22108 35492 22160
rect 35808 22040 35860 22092
rect 35900 21947 35952 21956
rect 35900 21913 35909 21947
rect 35909 21913 35943 21947
rect 35943 21913 35952 21947
rect 35900 21904 35952 21913
rect 34152 21836 34204 21888
rect 34796 21836 34848 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2596 21632 2648 21684
rect 5908 21632 5960 21684
rect 7012 21632 7064 21684
rect 8208 21632 8260 21684
rect 2504 21564 2556 21616
rect 5264 21564 5316 21616
rect 2412 21539 2464 21548
rect 2412 21505 2421 21539
rect 2421 21505 2455 21539
rect 2455 21505 2464 21539
rect 2412 21496 2464 21505
rect 3884 21496 3936 21548
rect 3976 21496 4028 21548
rect 4528 21496 4580 21548
rect 2964 21471 3016 21480
rect 2964 21437 2973 21471
rect 2973 21437 3007 21471
rect 3007 21437 3016 21471
rect 2964 21428 3016 21437
rect 3056 21471 3108 21480
rect 3056 21437 3065 21471
rect 3065 21437 3099 21471
rect 3099 21437 3108 21471
rect 3056 21428 3108 21437
rect 6000 21564 6052 21616
rect 6644 21564 6696 21616
rect 8852 21564 8904 21616
rect 13360 21675 13412 21684
rect 13360 21641 13369 21675
rect 13369 21641 13403 21675
rect 13403 21641 13412 21675
rect 13360 21632 13412 21641
rect 15476 21632 15528 21684
rect 16764 21632 16816 21684
rect 17684 21632 17736 21684
rect 19984 21632 20036 21684
rect 22100 21632 22152 21684
rect 25136 21632 25188 21684
rect 25964 21632 26016 21684
rect 27896 21675 27948 21684
rect 27896 21641 27905 21675
rect 27905 21641 27939 21675
rect 27939 21641 27948 21675
rect 27896 21632 27948 21641
rect 29736 21632 29788 21684
rect 30104 21632 30156 21684
rect 31208 21632 31260 21684
rect 32128 21632 32180 21684
rect 32404 21632 32456 21684
rect 32864 21675 32916 21684
rect 32864 21641 32873 21675
rect 32873 21641 32907 21675
rect 32907 21641 32916 21675
rect 32864 21632 32916 21641
rect 34152 21632 34204 21684
rect 34336 21632 34388 21684
rect 6184 21496 6236 21548
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 7748 21360 7800 21412
rect 2504 21335 2556 21344
rect 2504 21301 2513 21335
rect 2513 21301 2547 21335
rect 2547 21301 2556 21335
rect 2504 21292 2556 21301
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 5540 21292 5592 21301
rect 5724 21335 5776 21344
rect 5724 21301 5733 21335
rect 5733 21301 5767 21335
rect 5767 21301 5776 21335
rect 5724 21292 5776 21301
rect 9312 21539 9364 21548
rect 9312 21505 9321 21539
rect 9321 21505 9355 21539
rect 9355 21505 9364 21539
rect 9312 21496 9364 21505
rect 9772 21496 9824 21548
rect 9864 21539 9916 21548
rect 9864 21505 9873 21539
rect 9873 21505 9907 21539
rect 9907 21505 9916 21539
rect 9864 21496 9916 21505
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 10692 21496 10744 21548
rect 10324 21428 10376 21480
rect 12900 21564 12952 21616
rect 13360 21539 13412 21548
rect 13360 21505 13369 21539
rect 13369 21505 13403 21539
rect 13403 21505 13412 21539
rect 13360 21496 13412 21505
rect 12900 21428 12952 21480
rect 15200 21564 15252 21616
rect 16396 21607 16448 21616
rect 16396 21573 16405 21607
rect 16405 21573 16439 21607
rect 16439 21573 16448 21607
rect 16396 21564 16448 21573
rect 14924 21496 14976 21548
rect 15016 21496 15068 21548
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 16212 21539 16264 21548
rect 16212 21505 16221 21539
rect 16221 21505 16255 21539
rect 16255 21505 16264 21539
rect 16212 21496 16264 21505
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 9404 21360 9456 21412
rect 9772 21292 9824 21344
rect 16764 21360 16816 21412
rect 17224 21360 17276 21412
rect 17592 21496 17644 21548
rect 17776 21496 17828 21548
rect 17960 21539 18012 21548
rect 17960 21505 17969 21539
rect 17969 21505 18003 21539
rect 18003 21505 18012 21539
rect 17960 21496 18012 21505
rect 18880 21564 18932 21616
rect 19064 21496 19116 21548
rect 17960 21360 18012 21412
rect 19432 21428 19484 21480
rect 18880 21360 18932 21412
rect 20720 21564 20772 21616
rect 21272 21564 21324 21616
rect 22652 21564 22704 21616
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 22376 21496 22428 21548
rect 22836 21496 22888 21548
rect 24676 21564 24728 21616
rect 20720 21428 20772 21480
rect 20812 21428 20864 21480
rect 21364 21428 21416 21480
rect 22284 21428 22336 21480
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 19708 21360 19760 21412
rect 20168 21360 20220 21412
rect 21088 21360 21140 21412
rect 22008 21360 22060 21412
rect 25136 21496 25188 21548
rect 25228 21496 25280 21548
rect 25320 21496 25372 21548
rect 25780 21496 25832 21548
rect 25964 21539 26016 21548
rect 25964 21505 25973 21539
rect 25973 21505 26007 21539
rect 26007 21505 26016 21539
rect 25964 21496 26016 21505
rect 26792 21496 26844 21548
rect 27344 21539 27396 21548
rect 27344 21505 27353 21539
rect 27353 21505 27387 21539
rect 27387 21505 27396 21539
rect 27344 21496 27396 21505
rect 26976 21428 27028 21480
rect 27712 21539 27764 21548
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 27804 21428 27856 21480
rect 28448 21428 28500 21480
rect 17592 21292 17644 21344
rect 17684 21292 17736 21344
rect 17868 21292 17920 21344
rect 22284 21292 22336 21344
rect 22376 21292 22428 21344
rect 23020 21292 23072 21344
rect 28724 21496 28776 21548
rect 29184 21539 29236 21548
rect 29184 21505 29193 21539
rect 29193 21505 29227 21539
rect 29227 21505 29236 21539
rect 29184 21496 29236 21505
rect 29920 21428 29972 21480
rect 30196 21496 30248 21548
rect 31484 21496 31536 21548
rect 31852 21539 31904 21548
rect 31852 21505 31861 21539
rect 31861 21505 31895 21539
rect 31895 21505 31904 21539
rect 31852 21496 31904 21505
rect 32036 21496 32088 21548
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 32588 21539 32640 21548
rect 32588 21505 32597 21539
rect 32597 21505 32631 21539
rect 32631 21505 32640 21539
rect 32588 21496 32640 21505
rect 32772 21539 32824 21548
rect 32772 21505 32781 21539
rect 32781 21505 32815 21539
rect 32815 21505 32824 21539
rect 32772 21496 32824 21505
rect 33140 21496 33192 21548
rect 34060 21539 34112 21548
rect 34060 21505 34069 21539
rect 34069 21505 34103 21539
rect 34103 21505 34112 21539
rect 34060 21496 34112 21505
rect 34704 21539 34756 21548
rect 34704 21505 34713 21539
rect 34713 21505 34747 21539
rect 34747 21505 34756 21539
rect 34704 21496 34756 21505
rect 33324 21428 33376 21480
rect 24952 21292 25004 21344
rect 25228 21335 25280 21344
rect 25228 21301 25237 21335
rect 25237 21301 25271 21335
rect 25271 21301 25280 21335
rect 25228 21292 25280 21301
rect 29460 21292 29512 21344
rect 29920 21292 29972 21344
rect 30472 21360 30524 21412
rect 30932 21292 30984 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1676 21088 1728 21140
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 3884 20952 3936 21004
rect 4068 20952 4120 21004
rect 4620 21088 4672 21140
rect 5540 21088 5592 21140
rect 9220 21088 9272 21140
rect 10784 21131 10836 21140
rect 10784 21097 10793 21131
rect 10793 21097 10827 21131
rect 10827 21097 10836 21131
rect 10784 21088 10836 21097
rect 12440 21088 12492 21140
rect 14740 21131 14792 21140
rect 14740 21097 14749 21131
rect 14749 21097 14783 21131
rect 14783 21097 14792 21131
rect 14740 21088 14792 21097
rect 16580 21088 16632 21140
rect 17316 21131 17368 21140
rect 17316 21097 17325 21131
rect 17325 21097 17359 21131
rect 17359 21097 17368 21131
rect 17316 21088 17368 21097
rect 17500 21088 17552 21140
rect 17776 21088 17828 21140
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 3240 20816 3292 20868
rect 4160 20816 4212 20868
rect 5632 20927 5684 20936
rect 5632 20893 5641 20927
rect 5641 20893 5675 20927
rect 5675 20893 5684 20927
rect 5632 20884 5684 20893
rect 10324 21020 10376 21072
rect 9128 20884 9180 20936
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 10324 20884 10376 20936
rect 10416 20927 10468 20936
rect 10416 20893 10425 20927
rect 10425 20893 10459 20927
rect 10459 20893 10468 20927
rect 10416 20884 10468 20893
rect 10692 20884 10744 20936
rect 11152 20884 11204 20936
rect 12256 20927 12308 20936
rect 12256 20893 12265 20927
rect 12265 20893 12299 20927
rect 12299 20893 12308 20927
rect 12256 20884 12308 20893
rect 17868 21020 17920 21072
rect 12716 20927 12768 20936
rect 12716 20893 12719 20927
rect 12719 20893 12768 20927
rect 12716 20884 12768 20893
rect 13360 20884 13412 20936
rect 14464 20952 14516 21004
rect 9404 20816 9456 20868
rect 9864 20859 9916 20868
rect 9864 20825 9873 20859
rect 9873 20825 9907 20859
rect 9907 20825 9916 20859
rect 9864 20816 9916 20825
rect 10140 20816 10192 20868
rect 12164 20816 12216 20868
rect 3700 20748 3752 20800
rect 4436 20748 4488 20800
rect 5264 20791 5316 20800
rect 5264 20757 5273 20791
rect 5273 20757 5307 20791
rect 5307 20757 5316 20791
rect 5264 20748 5316 20757
rect 9680 20748 9732 20800
rect 9956 20748 10008 20800
rect 10416 20748 10468 20800
rect 13820 20748 13872 20800
rect 15016 20884 15068 20936
rect 14740 20816 14792 20868
rect 14372 20748 14424 20800
rect 15200 20748 15252 20800
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 16488 20884 16540 20936
rect 17592 20952 17644 21004
rect 18880 21020 18932 21072
rect 19432 20952 19484 21004
rect 21916 21020 21968 21072
rect 20168 20952 20220 21004
rect 22376 20952 22428 21004
rect 17776 20927 17828 20936
rect 15752 20816 15804 20868
rect 16580 20816 16632 20868
rect 17776 20893 17783 20927
rect 17783 20893 17817 20927
rect 17817 20893 17828 20927
rect 17776 20884 17828 20893
rect 17960 20884 18012 20936
rect 18328 20927 18380 20936
rect 18328 20893 18337 20927
rect 18337 20893 18371 20927
rect 18371 20893 18380 20927
rect 18328 20884 18380 20893
rect 15660 20748 15712 20800
rect 16028 20748 16080 20800
rect 17684 20748 17736 20800
rect 18604 20859 18656 20868
rect 18604 20825 18613 20859
rect 18613 20825 18647 20859
rect 18647 20825 18656 20859
rect 18604 20816 18656 20825
rect 18880 20884 18932 20936
rect 19064 20884 19116 20936
rect 18972 20791 19024 20800
rect 18972 20757 18981 20791
rect 18981 20757 19015 20791
rect 19015 20757 19024 20791
rect 18972 20748 19024 20757
rect 19432 20859 19484 20868
rect 19432 20825 19441 20859
rect 19441 20825 19475 20859
rect 19475 20825 19484 20859
rect 19432 20816 19484 20825
rect 19708 20748 19760 20800
rect 20720 20884 20772 20936
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 21088 20884 21140 20936
rect 21456 20884 21508 20936
rect 23756 21131 23808 21140
rect 23756 21097 23765 21131
rect 23765 21097 23799 21131
rect 23799 21097 23808 21131
rect 23756 21088 23808 21097
rect 26884 21088 26936 21140
rect 27160 21088 27212 21140
rect 27620 21088 27672 21140
rect 24124 20952 24176 21004
rect 24492 20884 24544 20936
rect 24124 20816 24176 20868
rect 24860 20816 24912 20868
rect 25044 20995 25096 21004
rect 25044 20961 25053 20995
rect 25053 20961 25087 20995
rect 25087 20961 25096 20995
rect 25044 20952 25096 20961
rect 25136 20952 25188 21004
rect 25412 20995 25464 21004
rect 25412 20961 25421 20995
rect 25421 20961 25455 20995
rect 25455 20961 25464 20995
rect 25412 20952 25464 20961
rect 28356 21020 28408 21072
rect 34796 21088 34848 21140
rect 26792 20884 26844 20936
rect 27160 20884 27212 20936
rect 27252 20884 27304 20936
rect 29828 20927 29880 20936
rect 29828 20893 29837 20927
rect 29837 20893 29871 20927
rect 29871 20893 29880 20927
rect 29828 20884 29880 20893
rect 29920 20884 29972 20936
rect 26056 20816 26108 20868
rect 26332 20816 26384 20868
rect 26976 20859 27028 20868
rect 26976 20825 26985 20859
rect 26985 20825 27019 20859
rect 27019 20825 27028 20859
rect 26976 20816 27028 20825
rect 20168 20748 20220 20800
rect 24216 20791 24268 20800
rect 24216 20757 24225 20791
rect 24225 20757 24259 20791
rect 24259 20757 24268 20791
rect 24216 20748 24268 20757
rect 31300 20884 31352 20936
rect 32496 20952 32548 21004
rect 34704 20952 34756 21004
rect 35900 20952 35952 21004
rect 34520 20884 34572 20936
rect 35164 20927 35216 20936
rect 35164 20893 35173 20927
rect 35173 20893 35207 20927
rect 35207 20893 35216 20927
rect 35164 20884 35216 20893
rect 31116 20748 31168 20800
rect 33048 20748 33100 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 38384 20680 38436 20732
rect 940 20544 992 20596
rect 1676 20544 1728 20596
rect 2504 20544 2556 20596
rect 2964 20544 3016 20596
rect 3608 20544 3660 20596
rect 1768 20476 1820 20528
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 4896 20544 4948 20596
rect 8576 20587 8628 20596
rect 8576 20553 8585 20587
rect 8585 20553 8619 20587
rect 8619 20553 8628 20587
rect 8576 20544 8628 20553
rect 9496 20544 9548 20596
rect 1492 20204 1544 20256
rect 3240 20383 3292 20392
rect 3240 20349 3249 20383
rect 3249 20349 3283 20383
rect 3283 20349 3292 20383
rect 3240 20340 3292 20349
rect 3700 20451 3752 20460
rect 3700 20417 3709 20451
rect 3709 20417 3743 20451
rect 3743 20417 3752 20451
rect 3700 20408 3752 20417
rect 4068 20451 4120 20460
rect 4068 20417 4077 20451
rect 4077 20417 4111 20451
rect 4111 20417 4120 20451
rect 4068 20408 4120 20417
rect 4436 20476 4488 20528
rect 4252 20408 4304 20460
rect 4896 20408 4948 20460
rect 7104 20383 7156 20392
rect 7104 20349 7113 20383
rect 7113 20349 7147 20383
rect 7147 20349 7156 20383
rect 7104 20340 7156 20349
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 9312 20451 9364 20460
rect 9312 20417 9321 20451
rect 9321 20417 9355 20451
rect 9355 20417 9364 20451
rect 9312 20408 9364 20417
rect 10508 20544 10560 20596
rect 10876 20587 10928 20596
rect 10876 20553 10885 20587
rect 10885 20553 10919 20587
rect 10919 20553 10928 20587
rect 10876 20544 10928 20553
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 9772 20476 9824 20528
rect 10232 20476 10284 20528
rect 9956 20451 10008 20460
rect 9956 20417 9965 20451
rect 9965 20417 9999 20451
rect 9999 20417 10008 20451
rect 9956 20408 10008 20417
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 10416 20408 10468 20460
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 14188 20544 14240 20596
rect 14280 20544 14332 20596
rect 14740 20544 14792 20596
rect 15108 20544 15160 20596
rect 16764 20544 16816 20596
rect 16580 20476 16632 20528
rect 17316 20476 17368 20528
rect 17684 20476 17736 20528
rect 18328 20476 18380 20528
rect 18604 20476 18656 20528
rect 19064 20476 19116 20528
rect 5816 20204 5868 20256
rect 6920 20204 6972 20256
rect 8300 20204 8352 20256
rect 11244 20272 11296 20324
rect 13728 20408 13780 20460
rect 9772 20204 9824 20256
rect 10416 20204 10468 20256
rect 12440 20204 12492 20256
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 14096 20408 14148 20417
rect 14372 20408 14424 20460
rect 14556 20408 14608 20460
rect 14464 20340 14516 20392
rect 15108 20451 15160 20460
rect 15108 20417 15122 20451
rect 15122 20417 15156 20451
rect 15156 20417 15160 20451
rect 15108 20408 15160 20417
rect 15476 20408 15528 20460
rect 15660 20408 15712 20460
rect 17224 20408 17276 20460
rect 24124 20544 24176 20596
rect 23664 20476 23716 20528
rect 20076 20451 20128 20460
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20260 20408 20312 20417
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 20812 20451 20864 20460
rect 20812 20417 20821 20451
rect 20821 20417 20855 20451
rect 20855 20417 20864 20451
rect 20812 20408 20864 20417
rect 21272 20451 21324 20460
rect 21272 20417 21281 20451
rect 21281 20417 21315 20451
rect 21315 20417 21324 20451
rect 21272 20408 21324 20417
rect 22284 20408 22336 20460
rect 23020 20408 23072 20460
rect 23940 20408 23992 20460
rect 33968 20544 34020 20596
rect 35900 20544 35952 20596
rect 25044 20408 25096 20460
rect 25412 20451 25464 20460
rect 25412 20417 25421 20451
rect 25421 20417 25455 20451
rect 25455 20417 25464 20451
rect 25412 20408 25464 20417
rect 25504 20451 25556 20460
rect 25504 20417 25513 20451
rect 25513 20417 25547 20451
rect 25547 20417 25556 20451
rect 25504 20408 25556 20417
rect 25688 20408 25740 20460
rect 25780 20408 25832 20460
rect 29000 20476 29052 20528
rect 28908 20451 28960 20460
rect 28908 20417 28917 20451
rect 28917 20417 28951 20451
rect 28951 20417 28960 20451
rect 28908 20408 28960 20417
rect 14740 20272 14792 20324
rect 15200 20272 15252 20324
rect 14556 20204 14608 20256
rect 17040 20383 17092 20392
rect 17040 20349 17049 20383
rect 17049 20349 17083 20383
rect 17083 20349 17092 20383
rect 17040 20340 17092 20349
rect 17684 20340 17736 20392
rect 18052 20340 18104 20392
rect 18696 20340 18748 20392
rect 23756 20340 23808 20392
rect 29368 20408 29420 20460
rect 29460 20408 29512 20460
rect 29552 20408 29604 20460
rect 30104 20408 30156 20460
rect 34796 20408 34848 20460
rect 29920 20383 29972 20392
rect 15844 20272 15896 20324
rect 19984 20272 20036 20324
rect 23388 20315 23440 20324
rect 23388 20281 23397 20315
rect 23397 20281 23431 20315
rect 23431 20281 23440 20315
rect 23388 20272 23440 20281
rect 24952 20272 25004 20324
rect 27528 20272 27580 20324
rect 29920 20349 29929 20383
rect 29929 20349 29963 20383
rect 29963 20349 29972 20383
rect 29920 20340 29972 20349
rect 33876 20340 33928 20392
rect 34428 20340 34480 20392
rect 35440 20383 35492 20392
rect 35440 20349 35449 20383
rect 35449 20349 35483 20383
rect 35483 20349 35492 20383
rect 35440 20340 35492 20349
rect 35348 20272 35400 20324
rect 36176 20451 36228 20460
rect 36176 20417 36185 20451
rect 36185 20417 36219 20451
rect 36219 20417 36228 20451
rect 36176 20408 36228 20417
rect 36268 20451 36320 20460
rect 36268 20417 36277 20451
rect 36277 20417 36311 20451
rect 36311 20417 36320 20451
rect 36268 20408 36320 20417
rect 16212 20204 16264 20256
rect 18972 20204 19024 20256
rect 21088 20204 21140 20256
rect 23204 20247 23256 20256
rect 23204 20213 23213 20247
rect 23213 20213 23247 20247
rect 23247 20213 23256 20247
rect 23204 20204 23256 20213
rect 28448 20204 28500 20256
rect 28632 20247 28684 20256
rect 28632 20213 28641 20247
rect 28641 20213 28675 20247
rect 28675 20213 28684 20247
rect 28632 20204 28684 20213
rect 29092 20204 29144 20256
rect 29276 20204 29328 20256
rect 29460 20247 29512 20256
rect 29460 20213 29469 20247
rect 29469 20213 29503 20247
rect 29503 20213 29512 20247
rect 29460 20204 29512 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7104 20000 7156 20052
rect 9312 20000 9364 20052
rect 14004 20000 14056 20052
rect 14096 20000 14148 20052
rect 15108 20000 15160 20052
rect 17408 20000 17460 20052
rect 18420 20043 18472 20052
rect 18420 20009 18429 20043
rect 18429 20009 18463 20043
rect 18463 20009 18472 20043
rect 18420 20000 18472 20009
rect 18972 20043 19024 20052
rect 18972 20009 18981 20043
rect 18981 20009 19015 20043
rect 19015 20009 19024 20043
rect 18972 20000 19024 20009
rect 20352 20000 20404 20052
rect 21456 20043 21508 20052
rect 21456 20009 21465 20043
rect 21465 20009 21499 20043
rect 21499 20009 21508 20043
rect 21456 20000 21508 20009
rect 23204 20000 23256 20052
rect 26608 20000 26660 20052
rect 11612 19932 11664 19984
rect 11796 19932 11848 19984
rect 14372 19975 14424 19984
rect 14372 19941 14381 19975
rect 14381 19941 14415 19975
rect 14415 19941 14424 19975
rect 14372 19932 14424 19941
rect 3884 19864 3936 19916
rect 5724 19907 5776 19916
rect 5724 19873 5733 19907
rect 5733 19873 5767 19907
rect 5767 19873 5776 19907
rect 5724 19864 5776 19873
rect 8024 19864 8076 19916
rect 8576 19864 8628 19916
rect 11888 19864 11940 19916
rect 12256 19864 12308 19916
rect 14740 19864 14792 19916
rect 15200 19864 15252 19916
rect 15660 19932 15712 19984
rect 3148 19796 3200 19848
rect 4160 19796 4212 19848
rect 5448 19796 5500 19848
rect 5816 19796 5868 19848
rect 3240 19728 3292 19780
rect 2688 19703 2740 19712
rect 2688 19669 2697 19703
rect 2697 19669 2731 19703
rect 2731 19669 2740 19703
rect 2688 19660 2740 19669
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 3884 19703 3936 19712
rect 3884 19669 3893 19703
rect 3893 19669 3927 19703
rect 3927 19669 3936 19703
rect 3884 19660 3936 19669
rect 5908 19660 5960 19712
rect 6000 19703 6052 19712
rect 6000 19669 6009 19703
rect 6009 19669 6043 19703
rect 6043 19669 6052 19703
rect 6000 19660 6052 19669
rect 9864 19728 9916 19780
rect 11152 19728 11204 19780
rect 9312 19660 9364 19712
rect 9588 19660 9640 19712
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 12808 19728 12860 19780
rect 13452 19728 13504 19780
rect 15476 19728 15528 19780
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 15844 19932 15896 19984
rect 16028 19839 16080 19848
rect 16028 19805 16037 19839
rect 16037 19805 16071 19839
rect 16071 19805 16080 19839
rect 16028 19796 16080 19805
rect 17040 19864 17092 19916
rect 16488 19796 16540 19848
rect 16856 19796 16908 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 20076 19932 20128 19984
rect 24216 19932 24268 19984
rect 17868 19864 17920 19916
rect 19432 19864 19484 19916
rect 20168 19864 20220 19916
rect 28264 20000 28316 20052
rect 28908 20000 28960 20052
rect 34796 20000 34848 20052
rect 36176 20000 36228 20052
rect 29276 19932 29328 19984
rect 12624 19660 12676 19712
rect 18696 19796 18748 19848
rect 19248 19796 19300 19848
rect 17868 19728 17920 19780
rect 18420 19728 18472 19780
rect 19064 19660 19116 19712
rect 22560 19796 22612 19848
rect 24032 19839 24084 19848
rect 20536 19660 20588 19712
rect 20628 19660 20680 19712
rect 22928 19728 22980 19780
rect 24032 19805 24041 19839
rect 24041 19805 24075 19839
rect 24075 19805 24084 19839
rect 24032 19796 24084 19805
rect 24676 19839 24728 19848
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 24952 19796 25004 19848
rect 25596 19796 25648 19848
rect 25872 19839 25924 19848
rect 25872 19805 25881 19839
rect 25881 19805 25915 19839
rect 25915 19805 25924 19839
rect 25872 19796 25924 19805
rect 25964 19796 26016 19848
rect 26884 19796 26936 19848
rect 27896 19864 27948 19916
rect 25688 19771 25740 19780
rect 25688 19737 25697 19771
rect 25697 19737 25731 19771
rect 25731 19737 25740 19771
rect 25688 19728 25740 19737
rect 25780 19771 25832 19780
rect 25780 19737 25789 19771
rect 25789 19737 25823 19771
rect 25823 19737 25832 19771
rect 25780 19728 25832 19737
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 28448 19864 28500 19916
rect 29000 19864 29052 19916
rect 28724 19796 28776 19848
rect 29552 19839 29604 19848
rect 29552 19805 29561 19839
rect 29561 19805 29595 19839
rect 29595 19805 29604 19839
rect 29552 19796 29604 19805
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 30104 19839 30156 19848
rect 30104 19805 30113 19839
rect 30113 19805 30147 19839
rect 30147 19805 30156 19839
rect 30104 19796 30156 19805
rect 33232 19796 33284 19848
rect 34704 19932 34756 19984
rect 35348 19932 35400 19984
rect 23940 19703 23992 19712
rect 23940 19669 23949 19703
rect 23949 19669 23983 19703
rect 23983 19669 23992 19703
rect 23940 19660 23992 19669
rect 24400 19660 24452 19712
rect 25596 19660 25648 19712
rect 30288 19771 30340 19780
rect 30288 19737 30297 19771
rect 30297 19737 30331 19771
rect 30331 19737 30340 19771
rect 30288 19728 30340 19737
rect 30840 19728 30892 19780
rect 28172 19703 28224 19712
rect 28172 19669 28181 19703
rect 28181 19669 28215 19703
rect 28215 19669 28224 19703
rect 28172 19660 28224 19669
rect 28264 19660 28316 19712
rect 29184 19660 29236 19712
rect 30472 19660 30524 19712
rect 33232 19703 33284 19712
rect 33232 19669 33241 19703
rect 33241 19669 33275 19703
rect 33275 19669 33284 19703
rect 33232 19660 33284 19669
rect 34244 19703 34296 19712
rect 34244 19669 34253 19703
rect 34253 19669 34287 19703
rect 34287 19669 34296 19703
rect 34244 19660 34296 19669
rect 34520 19660 34572 19712
rect 35072 19839 35124 19848
rect 35072 19805 35081 19839
rect 35081 19805 35115 19839
rect 35115 19805 35124 19839
rect 35072 19796 35124 19805
rect 35900 19796 35952 19848
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 2688 19456 2740 19508
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 4712 19456 4764 19508
rect 6920 19456 6972 19508
rect 9312 19499 9364 19508
rect 9312 19465 9321 19499
rect 9321 19465 9355 19499
rect 9355 19465 9364 19499
rect 9312 19456 9364 19465
rect 6000 19388 6052 19440
rect 10876 19388 10928 19440
rect 11152 19456 11204 19508
rect 15108 19456 15160 19508
rect 15200 19456 15252 19508
rect 15568 19456 15620 19508
rect 16580 19456 16632 19508
rect 11060 19388 11112 19440
rect 5908 19320 5960 19372
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 4620 19252 4672 19304
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 7196 19320 7248 19372
rect 7564 19320 7616 19372
rect 8668 19320 8720 19372
rect 9588 19320 9640 19372
rect 10968 19320 11020 19372
rect 12992 19320 13044 19372
rect 8944 19295 8996 19304
rect 8944 19261 8953 19295
rect 8953 19261 8987 19295
rect 8987 19261 8996 19295
rect 8944 19252 8996 19261
rect 10784 19252 10836 19304
rect 11520 19252 11572 19304
rect 12532 19252 12584 19304
rect 6828 19184 6880 19236
rect 11888 19184 11940 19236
rect 12716 19184 12768 19236
rect 13820 19320 13872 19372
rect 13636 19295 13688 19304
rect 13636 19261 13645 19295
rect 13645 19261 13679 19295
rect 13679 19261 13688 19295
rect 13636 19252 13688 19261
rect 14924 19320 14976 19372
rect 15476 19320 15528 19372
rect 17592 19431 17644 19440
rect 17592 19397 17601 19431
rect 17601 19397 17635 19431
rect 17635 19397 17644 19431
rect 17592 19388 17644 19397
rect 20168 19388 20220 19440
rect 24768 19456 24820 19508
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 15108 19252 15160 19304
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 2044 19116 2096 19168
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 5816 19116 5868 19168
rect 6000 19159 6052 19168
rect 6000 19125 6009 19159
rect 6009 19125 6043 19159
rect 6043 19125 6052 19159
rect 6000 19116 6052 19125
rect 7012 19116 7064 19168
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 9312 19116 9364 19168
rect 13084 19116 13136 19168
rect 13176 19159 13228 19168
rect 13176 19125 13185 19159
rect 13185 19125 13219 19159
rect 13219 19125 13228 19159
rect 13176 19116 13228 19125
rect 17132 19184 17184 19236
rect 17776 19227 17828 19236
rect 17776 19193 17785 19227
rect 17785 19193 17819 19227
rect 17819 19193 17828 19227
rect 17776 19184 17828 19193
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 19064 19320 19116 19372
rect 19432 19320 19484 19372
rect 19984 19320 20036 19372
rect 18972 19252 19024 19304
rect 20260 19252 20312 19304
rect 14924 19116 14976 19168
rect 17500 19116 17552 19168
rect 18972 19116 19024 19168
rect 19892 19116 19944 19168
rect 24216 19388 24268 19440
rect 25964 19456 26016 19508
rect 26424 19456 26476 19508
rect 27344 19456 27396 19508
rect 28172 19456 28224 19508
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22560 19320 22612 19372
rect 22928 19320 22980 19372
rect 23480 19320 23532 19372
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 23848 19320 23900 19372
rect 20904 19227 20956 19236
rect 20904 19193 20913 19227
rect 20913 19193 20947 19227
rect 20947 19193 20956 19227
rect 20904 19184 20956 19193
rect 23296 19227 23348 19236
rect 23296 19193 23305 19227
rect 23305 19193 23339 19227
rect 23339 19193 23348 19227
rect 23296 19184 23348 19193
rect 23848 19116 23900 19168
rect 24400 19363 24452 19372
rect 24400 19329 24409 19363
rect 24409 19329 24443 19363
rect 24443 19329 24452 19363
rect 24400 19320 24452 19329
rect 25688 19363 25740 19372
rect 25688 19329 25697 19363
rect 25697 19329 25731 19363
rect 25731 19329 25740 19363
rect 25688 19320 25740 19329
rect 26056 19363 26108 19372
rect 26056 19329 26065 19363
rect 26065 19329 26099 19363
rect 26099 19329 26108 19363
rect 26056 19320 26108 19329
rect 26332 19363 26384 19372
rect 26332 19329 26341 19363
rect 26341 19329 26375 19363
rect 26375 19329 26384 19363
rect 26332 19320 26384 19329
rect 26608 19320 26660 19372
rect 26792 19320 26844 19372
rect 24124 19184 24176 19236
rect 27252 19320 27304 19372
rect 27896 19320 27948 19372
rect 30012 19456 30064 19508
rect 30288 19456 30340 19508
rect 30472 19456 30524 19508
rect 33232 19456 33284 19508
rect 34428 19499 34480 19508
rect 34428 19465 34437 19499
rect 34437 19465 34471 19499
rect 34471 19465 34480 19499
rect 34428 19456 34480 19465
rect 35072 19456 35124 19508
rect 29184 19388 29236 19440
rect 28632 19320 28684 19372
rect 29000 19363 29052 19372
rect 29000 19329 29009 19363
rect 29009 19329 29043 19363
rect 29043 19329 29052 19363
rect 29000 19320 29052 19329
rect 29276 19320 29328 19372
rect 29460 19363 29512 19372
rect 29460 19329 29469 19363
rect 29469 19329 29503 19363
rect 29503 19329 29512 19363
rect 29460 19320 29512 19329
rect 24308 19184 24360 19236
rect 24860 19116 24912 19168
rect 30748 19388 30800 19440
rect 31208 19388 31260 19440
rect 30472 19363 30524 19372
rect 30472 19329 30481 19363
rect 30481 19329 30515 19363
rect 30515 19329 30524 19363
rect 30472 19320 30524 19329
rect 31944 19320 31996 19372
rect 32404 19320 32456 19372
rect 32588 19363 32640 19372
rect 32588 19329 32597 19363
rect 32597 19329 32631 19363
rect 32631 19329 32640 19363
rect 32588 19320 32640 19329
rect 30932 19252 30984 19304
rect 25136 19116 25188 19168
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 29184 19159 29236 19168
rect 29184 19125 29193 19159
rect 29193 19125 29227 19159
rect 29227 19125 29236 19159
rect 29184 19116 29236 19125
rect 29368 19116 29420 19168
rect 30472 19116 30524 19168
rect 31300 19116 31352 19168
rect 32220 19295 32272 19304
rect 32220 19261 32229 19295
rect 32229 19261 32263 19295
rect 32263 19261 32272 19295
rect 34244 19320 34296 19372
rect 32220 19252 32272 19261
rect 34520 19184 34572 19236
rect 35348 19184 35400 19236
rect 33324 19116 33376 19168
rect 34796 19116 34848 19168
rect 35716 19116 35768 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 3792 18955 3844 18964
rect 3792 18921 3801 18955
rect 3801 18921 3835 18955
rect 3835 18921 3844 18955
rect 3792 18912 3844 18921
rect 4620 18912 4672 18964
rect 7012 18912 7064 18964
rect 8668 18955 8720 18964
rect 8668 18921 8677 18955
rect 8677 18921 8711 18955
rect 8711 18921 8720 18955
rect 8668 18912 8720 18921
rect 10692 18912 10744 18964
rect 12164 18912 12216 18964
rect 12532 18955 12584 18964
rect 12532 18921 12541 18955
rect 12541 18921 12575 18955
rect 12575 18921 12584 18955
rect 12532 18912 12584 18921
rect 1768 18708 1820 18760
rect 2044 18751 2096 18760
rect 2044 18717 2053 18751
rect 2053 18717 2087 18751
rect 2087 18717 2096 18751
rect 2044 18708 2096 18717
rect 3240 18776 3292 18828
rect 8760 18844 8812 18896
rect 10416 18844 10468 18896
rect 10968 18887 11020 18896
rect 10968 18853 10977 18887
rect 10977 18853 11011 18887
rect 11011 18853 11020 18887
rect 10968 18844 11020 18853
rect 17592 18912 17644 18964
rect 17776 18912 17828 18964
rect 18144 18912 18196 18964
rect 19432 18912 19484 18964
rect 20168 18912 20220 18964
rect 20628 18955 20680 18964
rect 20628 18921 20637 18955
rect 20637 18921 20671 18955
rect 20671 18921 20680 18955
rect 20628 18912 20680 18921
rect 21916 18955 21968 18964
rect 21916 18921 21925 18955
rect 21925 18921 21959 18955
rect 21959 18921 21968 18955
rect 21916 18912 21968 18921
rect 3516 18708 3568 18760
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 4252 18751 4304 18760
rect 4252 18717 4261 18751
rect 4261 18717 4295 18751
rect 4295 18717 4304 18751
rect 4252 18708 4304 18717
rect 2964 18640 3016 18692
rect 5356 18640 5408 18692
rect 940 18572 992 18624
rect 2780 18615 2832 18624
rect 2780 18581 2789 18615
rect 2789 18581 2823 18615
rect 2823 18581 2832 18615
rect 2780 18572 2832 18581
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 6920 18819 6972 18828
rect 6920 18785 6929 18819
rect 6929 18785 6963 18819
rect 6963 18785 6972 18819
rect 13084 18844 13136 18896
rect 23296 18912 23348 18964
rect 23388 18955 23440 18964
rect 23388 18921 23397 18955
rect 23397 18921 23431 18955
rect 23431 18921 23440 18955
rect 23388 18912 23440 18921
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 23756 18955 23808 18964
rect 23756 18921 23765 18955
rect 23765 18921 23799 18955
rect 23799 18921 23808 18955
rect 23756 18912 23808 18921
rect 23940 18912 23992 18964
rect 24124 18912 24176 18964
rect 6920 18776 6972 18785
rect 8300 18708 8352 18760
rect 9128 18708 9180 18760
rect 10600 18708 10652 18760
rect 6000 18572 6052 18624
rect 6920 18572 6972 18624
rect 7472 18640 7524 18692
rect 10140 18640 10192 18692
rect 10968 18708 11020 18760
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 13084 18708 13136 18760
rect 16580 18776 16632 18828
rect 16764 18776 16816 18828
rect 18144 18776 18196 18828
rect 13820 18708 13872 18760
rect 10416 18615 10468 18624
rect 10416 18581 10425 18615
rect 10425 18581 10459 18615
rect 10459 18581 10468 18615
rect 10416 18572 10468 18581
rect 10600 18615 10652 18624
rect 10600 18581 10609 18615
rect 10609 18581 10643 18615
rect 10643 18581 10652 18615
rect 10600 18572 10652 18581
rect 11980 18572 12032 18624
rect 12808 18683 12860 18692
rect 12808 18649 12817 18683
rect 12817 18649 12851 18683
rect 12851 18649 12860 18683
rect 12808 18640 12860 18649
rect 12992 18683 13044 18692
rect 12992 18649 13001 18683
rect 13001 18649 13035 18683
rect 13035 18649 13044 18683
rect 12992 18640 13044 18649
rect 13268 18683 13320 18692
rect 13268 18649 13277 18683
rect 13277 18649 13311 18683
rect 13311 18649 13320 18683
rect 13268 18640 13320 18649
rect 13728 18640 13780 18692
rect 14372 18640 14424 18692
rect 14924 18683 14976 18692
rect 14924 18649 14933 18683
rect 14933 18649 14967 18683
rect 14967 18649 14976 18683
rect 14924 18640 14976 18649
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 16028 18640 16080 18692
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 13084 18572 13136 18624
rect 13636 18572 13688 18624
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 17592 18708 17644 18760
rect 19248 18708 19300 18760
rect 20536 18776 20588 18828
rect 21824 18776 21876 18828
rect 22468 18819 22520 18828
rect 22468 18785 22477 18819
rect 22477 18785 22511 18819
rect 22511 18785 22520 18819
rect 22468 18776 22520 18785
rect 17868 18640 17920 18692
rect 18052 18683 18104 18692
rect 18052 18649 18061 18683
rect 18061 18649 18095 18683
rect 18095 18649 18104 18683
rect 18052 18640 18104 18649
rect 18328 18640 18380 18692
rect 19064 18640 19116 18692
rect 20812 18708 20864 18760
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 22928 18844 22980 18896
rect 23112 18844 23164 18896
rect 24400 18844 24452 18896
rect 23020 18776 23072 18828
rect 23204 18776 23256 18828
rect 23848 18776 23900 18828
rect 24216 18819 24268 18828
rect 24216 18785 24231 18819
rect 24231 18785 24265 18819
rect 24265 18785 24268 18819
rect 26792 18912 26844 18964
rect 28724 18955 28776 18964
rect 28724 18921 28733 18955
rect 28733 18921 28767 18955
rect 28767 18921 28776 18955
rect 28724 18912 28776 18921
rect 24216 18776 24268 18785
rect 24768 18776 24820 18828
rect 22836 18751 22888 18760
rect 22836 18717 22845 18751
rect 22845 18717 22879 18751
rect 22879 18717 22888 18751
rect 22836 18708 22888 18717
rect 22928 18751 22980 18760
rect 22928 18717 22937 18751
rect 22937 18717 22971 18751
rect 22971 18717 22980 18751
rect 22928 18708 22980 18717
rect 20076 18640 20128 18692
rect 21364 18640 21416 18692
rect 20628 18572 20680 18624
rect 21272 18572 21324 18624
rect 22468 18572 22520 18624
rect 23388 18708 23440 18760
rect 24032 18708 24084 18760
rect 24124 18751 24176 18760
rect 24124 18717 24133 18751
rect 24133 18717 24167 18751
rect 24167 18717 24176 18751
rect 24124 18708 24176 18717
rect 25044 18708 25096 18760
rect 25780 18708 25832 18760
rect 26608 18776 26660 18828
rect 31760 18844 31812 18896
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 24860 18640 24912 18692
rect 25596 18640 25648 18692
rect 26424 18683 26476 18692
rect 26424 18649 26433 18683
rect 26433 18649 26467 18683
rect 26467 18649 26476 18683
rect 26424 18640 26476 18649
rect 25872 18572 25924 18624
rect 28816 18751 28868 18760
rect 28816 18717 28825 18751
rect 28825 18717 28859 18751
rect 28859 18717 28868 18751
rect 28816 18708 28868 18717
rect 29184 18708 29236 18760
rect 34704 18887 34756 18896
rect 34704 18853 34713 18887
rect 34713 18853 34747 18887
rect 34747 18853 34756 18887
rect 34704 18844 34756 18853
rect 31208 18751 31260 18760
rect 31208 18717 31217 18751
rect 31217 18717 31251 18751
rect 31251 18717 31260 18751
rect 31208 18708 31260 18717
rect 31944 18640 31996 18692
rect 32220 18708 32272 18760
rect 32588 18751 32640 18760
rect 32588 18717 32597 18751
rect 32597 18717 32631 18751
rect 32631 18717 32640 18751
rect 32588 18708 32640 18717
rect 32956 18640 33008 18692
rect 35532 18887 35584 18896
rect 35532 18853 35541 18887
rect 35541 18853 35575 18887
rect 35575 18853 35584 18887
rect 35532 18844 35584 18853
rect 35164 18819 35216 18828
rect 35164 18785 35173 18819
rect 35173 18785 35207 18819
rect 35207 18785 35216 18819
rect 35164 18776 35216 18785
rect 35440 18776 35492 18828
rect 32036 18572 32088 18624
rect 32312 18572 32364 18624
rect 32404 18572 32456 18624
rect 32772 18572 32824 18624
rect 35716 18683 35768 18692
rect 35716 18649 35725 18683
rect 35725 18649 35759 18683
rect 35759 18649 35768 18683
rect 35716 18640 35768 18649
rect 36268 18572 36320 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2412 18368 2464 18420
rect 2780 18368 2832 18420
rect 3516 18368 3568 18420
rect 4252 18368 4304 18420
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 4068 18232 4120 18284
rect 4160 18232 4212 18284
rect 6920 18343 6972 18352
rect 6920 18309 6929 18343
rect 6929 18309 6963 18343
rect 6963 18309 6972 18343
rect 6920 18300 6972 18309
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 8760 18300 8812 18352
rect 10600 18368 10652 18420
rect 12716 18368 12768 18420
rect 15568 18368 15620 18420
rect 16028 18368 16080 18420
rect 16304 18368 16356 18420
rect 16488 18368 16540 18420
rect 17132 18368 17184 18420
rect 18696 18411 18748 18420
rect 18696 18377 18705 18411
rect 18705 18377 18739 18411
rect 18739 18377 18748 18411
rect 18696 18368 18748 18377
rect 20720 18368 20772 18420
rect 21824 18368 21876 18420
rect 25136 18368 25188 18420
rect 25320 18368 25372 18420
rect 6828 18232 6880 18284
rect 7196 18232 7248 18284
rect 3884 18164 3936 18216
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2320 18071 2372 18080
rect 2320 18037 2329 18071
rect 2329 18037 2363 18071
rect 2363 18037 2372 18071
rect 2320 18028 2372 18037
rect 6736 18164 6788 18216
rect 8576 18232 8628 18284
rect 9036 18232 9088 18284
rect 9588 18232 9640 18284
rect 10140 18275 10192 18284
rect 10140 18241 10149 18275
rect 10149 18241 10183 18275
rect 10183 18241 10192 18275
rect 10140 18232 10192 18241
rect 10692 18232 10744 18284
rect 10968 18275 11020 18284
rect 10968 18241 10977 18275
rect 10977 18241 11011 18275
rect 11011 18241 11020 18275
rect 10968 18232 11020 18241
rect 10416 18164 10468 18216
rect 10600 18164 10652 18216
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 11796 18232 11848 18284
rect 19708 18300 19760 18352
rect 20904 18300 20956 18352
rect 21916 18300 21968 18352
rect 23848 18300 23900 18352
rect 24492 18300 24544 18352
rect 28356 18300 28408 18352
rect 32036 18368 32088 18420
rect 35164 18368 35216 18420
rect 35532 18368 35584 18420
rect 12532 18232 12584 18284
rect 13636 18232 13688 18284
rect 11980 18164 12032 18216
rect 12072 18164 12124 18216
rect 13084 18164 13136 18216
rect 13820 18164 13872 18216
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 15936 18232 15988 18284
rect 16120 18232 16172 18284
rect 17592 18232 17644 18284
rect 16488 18164 16540 18216
rect 16580 18164 16632 18216
rect 16764 18164 16816 18216
rect 17500 18164 17552 18216
rect 18512 18275 18564 18284
rect 18512 18241 18521 18275
rect 18521 18241 18555 18275
rect 18555 18241 18564 18275
rect 18512 18232 18564 18241
rect 18604 18232 18656 18284
rect 18972 18232 19024 18284
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 20076 18232 20128 18284
rect 20260 18232 20312 18284
rect 20812 18232 20864 18284
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 18420 18164 18472 18216
rect 23388 18232 23440 18284
rect 27160 18232 27212 18284
rect 22192 18164 22244 18216
rect 26700 18164 26752 18216
rect 27712 18164 27764 18216
rect 28356 18207 28408 18216
rect 28356 18173 28365 18207
rect 28365 18173 28399 18207
rect 28399 18173 28408 18207
rect 28356 18164 28408 18173
rect 30196 18232 30248 18284
rect 30104 18164 30156 18216
rect 31116 18164 31168 18216
rect 31760 18164 31812 18216
rect 32404 18164 32456 18216
rect 9588 18096 9640 18148
rect 9680 18096 9732 18148
rect 11060 18096 11112 18148
rect 12992 18096 13044 18148
rect 15568 18096 15620 18148
rect 32220 18096 32272 18148
rect 34704 18275 34756 18284
rect 34704 18241 34713 18275
rect 34713 18241 34747 18275
rect 34747 18241 34756 18275
rect 34704 18232 34756 18241
rect 34796 18207 34848 18216
rect 34796 18173 34805 18207
rect 34805 18173 34839 18207
rect 34839 18173 34848 18207
rect 34796 18164 34848 18173
rect 33416 18096 33468 18148
rect 11888 18028 11940 18080
rect 13728 18028 13780 18080
rect 15752 18028 15804 18080
rect 16304 18028 16356 18080
rect 17132 18028 17184 18080
rect 17868 18028 17920 18080
rect 18788 18028 18840 18080
rect 19064 18071 19116 18080
rect 19064 18037 19073 18071
rect 19073 18037 19107 18071
rect 19107 18037 19116 18071
rect 19064 18028 19116 18037
rect 21824 18028 21876 18080
rect 23388 18028 23440 18080
rect 26608 18028 26660 18080
rect 30472 18028 30524 18080
rect 30656 18028 30708 18080
rect 32772 18028 32824 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 38384 17960 38436 18012
rect 7564 17824 7616 17876
rect 9588 17824 9640 17876
rect 10140 17824 10192 17876
rect 10692 17824 10744 17876
rect 11336 17824 11388 17876
rect 11428 17867 11480 17876
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 11796 17824 11848 17876
rect 3056 17731 3108 17740
rect 3056 17697 3065 17731
rect 3065 17697 3099 17731
rect 3099 17697 3108 17731
rect 3056 17688 3108 17697
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 4252 17688 4304 17740
rect 6644 17756 6696 17808
rect 7472 17731 7524 17740
rect 7472 17697 7481 17731
rect 7481 17697 7515 17731
rect 7515 17697 7524 17731
rect 7472 17688 7524 17697
rect 8024 17688 8076 17740
rect 8668 17688 8720 17740
rect 9680 17688 9732 17740
rect 4436 17663 4488 17672
rect 4436 17629 4445 17663
rect 4445 17629 4479 17663
rect 4479 17629 4488 17663
rect 4436 17620 4488 17629
rect 5172 17620 5224 17672
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 4896 17552 4948 17604
rect 5080 17552 5132 17604
rect 6000 17552 6052 17604
rect 7196 17552 7248 17604
rect 10784 17731 10836 17740
rect 10784 17697 10793 17731
rect 10793 17697 10827 17731
rect 10827 17697 10836 17731
rect 10784 17688 10836 17697
rect 11152 17688 11204 17740
rect 5448 17484 5500 17536
rect 8668 17552 8720 17604
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 15384 17824 15436 17876
rect 16948 17824 17000 17876
rect 18512 17824 18564 17876
rect 20996 17824 21048 17876
rect 27160 17824 27212 17876
rect 30380 17824 30432 17876
rect 31208 17824 31260 17876
rect 32312 17824 32364 17876
rect 11520 17620 11572 17672
rect 11704 17620 11756 17672
rect 15292 17756 15344 17808
rect 15568 17756 15620 17808
rect 9772 17552 9824 17604
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 9588 17484 9640 17536
rect 10416 17484 10468 17536
rect 10968 17484 11020 17536
rect 11704 17484 11756 17536
rect 13084 17552 13136 17604
rect 13268 17552 13320 17604
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14556 17620 14608 17629
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 15200 17620 15252 17672
rect 12164 17484 12216 17536
rect 14004 17484 14056 17536
rect 14188 17484 14240 17536
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 15660 17620 15712 17672
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 16672 17731 16724 17740
rect 16672 17697 16681 17731
rect 16681 17697 16715 17731
rect 16715 17697 16724 17731
rect 16672 17688 16724 17697
rect 18696 17756 18748 17808
rect 20720 17756 20772 17808
rect 23296 17756 23348 17808
rect 18512 17688 18564 17740
rect 19800 17688 19852 17740
rect 19892 17688 19944 17740
rect 20260 17688 20312 17740
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 18420 17620 18472 17672
rect 19340 17663 19392 17672
rect 19340 17629 19349 17663
rect 19349 17629 19383 17663
rect 19383 17629 19392 17663
rect 19340 17620 19392 17629
rect 16580 17552 16632 17604
rect 16948 17552 17000 17604
rect 20076 17620 20128 17672
rect 20536 17620 20588 17672
rect 20904 17620 20956 17672
rect 15936 17484 15988 17536
rect 16028 17484 16080 17536
rect 18420 17484 18472 17536
rect 19616 17484 19668 17536
rect 20260 17552 20312 17604
rect 23848 17731 23900 17740
rect 23848 17697 23857 17731
rect 23857 17697 23891 17731
rect 23891 17697 23900 17731
rect 23848 17688 23900 17697
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 24216 17620 24268 17672
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 24952 17799 25004 17808
rect 24952 17765 24961 17799
rect 24961 17765 24995 17799
rect 24995 17765 25004 17799
rect 24952 17756 25004 17765
rect 25136 17688 25188 17740
rect 28908 17756 28960 17808
rect 30012 17756 30064 17808
rect 32220 17756 32272 17808
rect 25596 17620 25648 17672
rect 21272 17552 21324 17604
rect 24768 17552 24820 17604
rect 24952 17552 25004 17604
rect 26608 17552 26660 17604
rect 23940 17484 23992 17536
rect 27620 17688 27672 17740
rect 27988 17663 28040 17672
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 29460 17688 29512 17740
rect 29828 17663 29880 17672
rect 29828 17629 29837 17663
rect 29837 17629 29871 17663
rect 29871 17629 29880 17663
rect 29828 17620 29880 17629
rect 29920 17620 29972 17672
rect 30196 17552 30248 17604
rect 31392 17731 31444 17740
rect 31392 17697 31401 17731
rect 31401 17697 31435 17731
rect 31435 17697 31444 17731
rect 31392 17688 31444 17697
rect 31760 17731 31812 17740
rect 31760 17697 31770 17731
rect 31770 17697 31804 17731
rect 31804 17697 31812 17731
rect 33784 17824 33836 17876
rect 31760 17688 31812 17697
rect 30472 17663 30524 17672
rect 30472 17629 30481 17663
rect 30481 17629 30515 17663
rect 30515 17629 30524 17663
rect 30472 17620 30524 17629
rect 31576 17663 31628 17672
rect 31576 17629 31585 17663
rect 31585 17629 31619 17663
rect 31619 17629 31628 17663
rect 31576 17620 31628 17629
rect 31668 17663 31720 17672
rect 31668 17629 31677 17663
rect 31677 17629 31711 17663
rect 31711 17629 31720 17663
rect 31668 17620 31720 17629
rect 31852 17663 31904 17672
rect 31852 17629 31861 17663
rect 31861 17629 31895 17663
rect 31895 17629 31904 17663
rect 31852 17620 31904 17629
rect 32496 17620 32548 17672
rect 32864 17620 32916 17672
rect 33140 17688 33192 17740
rect 32772 17595 32824 17604
rect 32772 17561 32781 17595
rect 32781 17561 32815 17595
rect 32815 17561 32824 17595
rect 32772 17552 32824 17561
rect 33140 17595 33192 17604
rect 28724 17484 28776 17536
rect 31668 17484 31720 17536
rect 32680 17484 32732 17536
rect 33140 17561 33149 17595
rect 33149 17561 33183 17595
rect 33183 17561 33192 17595
rect 33140 17552 33192 17561
rect 33416 17620 33468 17672
rect 33784 17552 33836 17604
rect 34060 17527 34112 17536
rect 34060 17493 34069 17527
rect 34069 17493 34103 17527
rect 34103 17493 34112 17527
rect 34060 17484 34112 17493
rect 34428 17527 34480 17536
rect 34428 17493 34437 17527
rect 34437 17493 34471 17527
rect 34471 17493 34480 17527
rect 34428 17484 34480 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 5172 17280 5224 17332
rect 3976 17212 4028 17264
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 2780 17144 2832 17196
rect 1676 17119 1728 17128
rect 1676 17085 1685 17119
rect 1685 17085 1719 17119
rect 1719 17085 1728 17119
rect 1676 17076 1728 17085
rect 4712 17255 4764 17264
rect 4712 17221 4737 17255
rect 4737 17221 4764 17255
rect 4712 17212 4764 17221
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 5448 17280 5500 17332
rect 10784 17280 10836 17332
rect 11060 17280 11112 17332
rect 11152 17280 11204 17332
rect 11428 17280 11480 17332
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 13360 17280 13412 17332
rect 14372 17280 14424 17332
rect 16120 17280 16172 17332
rect 16488 17280 16540 17332
rect 16672 17280 16724 17332
rect 3976 17008 4028 17060
rect 4160 17008 4212 17060
rect 4804 17076 4856 17128
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 9772 17212 9824 17264
rect 5816 17119 5868 17128
rect 5816 17085 5825 17119
rect 5825 17085 5859 17119
rect 5859 17085 5868 17119
rect 5816 17076 5868 17085
rect 2872 16940 2924 16992
rect 4896 17051 4948 17060
rect 4896 17017 4905 17051
rect 4905 17017 4939 17051
rect 4939 17017 4948 17051
rect 4896 17008 4948 17017
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 5448 16940 5500 16992
rect 5540 16940 5592 16992
rect 6092 17076 6144 17128
rect 9680 17144 9732 17196
rect 10968 17144 11020 17196
rect 11244 17144 11296 17196
rect 11428 17144 11480 17196
rect 12348 17212 12400 17264
rect 13452 17255 13504 17264
rect 13452 17221 13461 17255
rect 13461 17221 13495 17255
rect 13495 17221 13504 17255
rect 13452 17212 13504 17221
rect 15292 17212 15344 17264
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 12164 17144 12216 17196
rect 6644 17008 6696 17060
rect 9956 17008 10008 17060
rect 12440 17144 12492 17196
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 9220 16940 9272 16992
rect 11428 16940 11480 16992
rect 12256 17008 12308 17060
rect 14188 16940 14240 16992
rect 14372 16940 14424 16992
rect 15384 17144 15436 17196
rect 15844 17212 15896 17264
rect 15752 17187 15804 17196
rect 15752 17153 15765 17187
rect 15765 17153 15804 17187
rect 15752 17144 15804 17153
rect 16028 17187 16080 17196
rect 16028 17153 16037 17187
rect 16037 17153 16071 17187
rect 16071 17153 16080 17187
rect 16028 17144 16080 17153
rect 16396 17212 16448 17264
rect 17500 17280 17552 17332
rect 16488 17144 16540 17196
rect 16948 17144 17000 17196
rect 18236 17212 18288 17264
rect 18420 17212 18472 17264
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 16304 16940 16356 16992
rect 16672 17076 16724 17128
rect 18328 17144 18380 17196
rect 18696 17280 18748 17332
rect 18880 17323 18932 17332
rect 18880 17289 18889 17323
rect 18889 17289 18923 17323
rect 18923 17289 18932 17323
rect 18880 17280 18932 17289
rect 19892 17280 19944 17332
rect 20260 17323 20312 17332
rect 20260 17289 20269 17323
rect 20269 17289 20303 17323
rect 20303 17289 20312 17323
rect 20260 17280 20312 17289
rect 17960 17076 18012 17128
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 18880 17076 18932 17128
rect 19892 17187 19944 17196
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 20076 17187 20128 17196
rect 20628 17280 20680 17332
rect 20720 17255 20772 17264
rect 20720 17221 20729 17255
rect 20729 17221 20763 17255
rect 20763 17221 20772 17255
rect 20720 17212 20772 17221
rect 21364 17280 21416 17332
rect 20076 17153 20090 17187
rect 20090 17153 20124 17187
rect 20124 17153 20128 17187
rect 20076 17144 20128 17153
rect 17132 16983 17184 16992
rect 17132 16949 17141 16983
rect 17141 16949 17175 16983
rect 17175 16949 17184 16983
rect 17132 16940 17184 16949
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 19892 17008 19944 17060
rect 20628 17187 20680 17196
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 20904 17144 20956 17196
rect 20996 17144 21048 17196
rect 21180 17144 21232 17196
rect 21088 17119 21140 17128
rect 21088 17085 21097 17119
rect 21097 17085 21131 17119
rect 21131 17085 21140 17119
rect 21088 17076 21140 17085
rect 23388 17144 23440 17196
rect 24584 17280 24636 17332
rect 25596 17280 25648 17332
rect 28080 17280 28132 17332
rect 28356 17323 28408 17332
rect 28356 17289 28365 17323
rect 28365 17289 28399 17323
rect 28399 17289 28408 17323
rect 28356 17280 28408 17289
rect 29460 17323 29512 17332
rect 29460 17289 29469 17323
rect 29469 17289 29503 17323
rect 29503 17289 29512 17323
rect 29460 17280 29512 17289
rect 31392 17280 31444 17332
rect 31576 17323 31628 17332
rect 31576 17289 31585 17323
rect 31585 17289 31619 17323
rect 31619 17289 31628 17323
rect 31576 17280 31628 17289
rect 31668 17280 31720 17332
rect 34060 17280 34112 17332
rect 24308 17144 24360 17196
rect 29092 17255 29144 17264
rect 29092 17221 29101 17255
rect 29101 17221 29135 17255
rect 29135 17221 29144 17255
rect 29092 17212 29144 17221
rect 29184 17212 29236 17264
rect 30472 17212 30524 17264
rect 34428 17280 34480 17332
rect 21548 17119 21600 17128
rect 21548 17085 21557 17119
rect 21557 17085 21591 17119
rect 21591 17085 21600 17119
rect 21548 17076 21600 17085
rect 23020 17076 23072 17128
rect 24216 17076 24268 17128
rect 25688 17076 25740 17128
rect 27068 17076 27120 17128
rect 28632 17187 28684 17196
rect 28632 17153 28641 17187
rect 28641 17153 28675 17187
rect 28675 17153 28684 17187
rect 28632 17144 28684 17153
rect 28724 17187 28776 17196
rect 28724 17153 28733 17187
rect 28733 17153 28767 17187
rect 28767 17153 28776 17187
rect 28724 17144 28776 17153
rect 28816 17187 28868 17196
rect 28816 17153 28825 17187
rect 28825 17153 28859 17187
rect 28859 17153 28868 17187
rect 28816 17144 28868 17153
rect 29000 17187 29052 17196
rect 29000 17153 29009 17187
rect 29009 17153 29043 17187
rect 29043 17153 29052 17187
rect 29000 17144 29052 17153
rect 31208 17187 31260 17196
rect 31208 17153 31217 17187
rect 31217 17153 31251 17187
rect 31251 17153 31260 17187
rect 31208 17144 31260 17153
rect 31576 17144 31628 17196
rect 31760 17144 31812 17196
rect 34520 17255 34572 17264
rect 34520 17221 34545 17255
rect 34545 17221 34572 17255
rect 34520 17212 34572 17221
rect 20352 17008 20404 17060
rect 20444 17008 20496 17060
rect 21180 16940 21232 16992
rect 22652 17051 22704 17060
rect 22652 17017 22661 17051
rect 22661 17017 22695 17051
rect 22695 17017 22704 17051
rect 22652 17008 22704 17017
rect 27988 17051 28040 17060
rect 27988 17017 27997 17051
rect 27997 17017 28031 17051
rect 28031 17017 28040 17051
rect 27988 17008 28040 17017
rect 24124 16940 24176 16992
rect 29184 16940 29236 16992
rect 34336 17076 34388 17128
rect 34520 17076 34572 17128
rect 34704 17076 34756 17128
rect 34980 17076 35032 17128
rect 35532 17255 35584 17264
rect 35532 17221 35541 17255
rect 35541 17221 35575 17255
rect 35575 17221 35584 17255
rect 35532 17212 35584 17221
rect 32404 17051 32456 17060
rect 32404 17017 32413 17051
rect 32413 17017 32447 17051
rect 32447 17017 32456 17051
rect 32404 17008 32456 17017
rect 34428 16940 34480 16992
rect 34520 16983 34572 16992
rect 34520 16949 34529 16983
rect 34529 16949 34563 16983
rect 34563 16949 34572 16983
rect 34520 16940 34572 16949
rect 34612 16940 34664 16992
rect 34980 16940 35032 16992
rect 35348 16940 35400 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1676 16736 1728 16788
rect 2504 16736 2556 16788
rect 3056 16736 3108 16788
rect 4528 16600 4580 16652
rect 4712 16668 4764 16720
rect 5172 16736 5224 16788
rect 5540 16668 5592 16720
rect 5816 16711 5868 16720
rect 5816 16677 5825 16711
rect 5825 16677 5859 16711
rect 5859 16677 5868 16711
rect 5816 16668 5868 16677
rect 7196 16736 7248 16788
rect 8484 16668 8536 16720
rect 6736 16600 6788 16652
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 9220 16600 9272 16652
rect 10048 16600 10100 16652
rect 15384 16736 15436 16788
rect 16488 16736 16540 16788
rect 18144 16736 18196 16788
rect 12808 16600 12860 16652
rect 4804 16532 4856 16584
rect 8300 16532 8352 16584
rect 9036 16532 9088 16584
rect 9496 16532 9548 16584
rect 13728 16600 13780 16652
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 15476 16600 15528 16652
rect 7196 16507 7248 16516
rect 7196 16473 7205 16507
rect 7205 16473 7239 16507
rect 7239 16473 7248 16507
rect 7196 16464 7248 16473
rect 13084 16464 13136 16516
rect 6184 16439 6236 16448
rect 6184 16405 6193 16439
rect 6193 16405 6227 16439
rect 6227 16405 6236 16439
rect 6184 16396 6236 16405
rect 9128 16396 9180 16448
rect 9404 16396 9456 16448
rect 9588 16396 9640 16448
rect 12624 16396 12676 16448
rect 12900 16439 12952 16448
rect 12900 16405 12909 16439
rect 12909 16405 12943 16439
rect 12943 16405 12952 16439
rect 12900 16396 12952 16405
rect 15292 16532 15344 16584
rect 16488 16532 16540 16584
rect 16764 16532 16816 16584
rect 18512 16600 18564 16652
rect 20444 16736 20496 16788
rect 20536 16736 20588 16788
rect 20996 16779 21048 16788
rect 20996 16745 21005 16779
rect 21005 16745 21039 16779
rect 21039 16745 21048 16779
rect 20996 16736 21048 16745
rect 21180 16779 21232 16788
rect 21180 16745 21189 16779
rect 21189 16745 21223 16779
rect 21223 16745 21232 16779
rect 21180 16736 21232 16745
rect 19616 16668 19668 16720
rect 20352 16668 20404 16720
rect 26884 16736 26936 16788
rect 24952 16668 25004 16720
rect 32404 16736 32456 16788
rect 34704 16736 34756 16788
rect 35348 16736 35400 16788
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 18788 16532 18840 16584
rect 19064 16532 19116 16584
rect 19432 16532 19484 16584
rect 19800 16532 19852 16584
rect 19984 16532 20036 16584
rect 14832 16507 14884 16516
rect 14832 16473 14841 16507
rect 14841 16473 14875 16507
rect 14875 16473 14884 16507
rect 14832 16464 14884 16473
rect 15660 16464 15712 16516
rect 14464 16396 14516 16448
rect 14556 16396 14608 16448
rect 17316 16396 17368 16448
rect 17592 16439 17644 16448
rect 17592 16405 17601 16439
rect 17601 16405 17635 16439
rect 17635 16405 17644 16439
rect 17592 16396 17644 16405
rect 17960 16507 18012 16516
rect 17960 16473 17969 16507
rect 17969 16473 18003 16507
rect 18003 16473 18012 16507
rect 17960 16464 18012 16473
rect 19616 16464 19668 16516
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 20444 16532 20496 16584
rect 20720 16532 20772 16584
rect 21180 16532 21232 16584
rect 23112 16643 23164 16652
rect 23112 16609 23121 16643
rect 23121 16609 23155 16643
rect 23155 16609 23164 16643
rect 23112 16600 23164 16609
rect 24124 16600 24176 16652
rect 27252 16600 27304 16652
rect 28632 16600 28684 16652
rect 32496 16600 32548 16652
rect 34796 16643 34848 16652
rect 34796 16609 34805 16643
rect 34805 16609 34839 16643
rect 34839 16609 34848 16643
rect 34796 16600 34848 16609
rect 21272 16464 21324 16516
rect 22008 16507 22060 16516
rect 22008 16473 22017 16507
rect 22017 16473 22051 16507
rect 22051 16473 22060 16507
rect 22008 16464 22060 16473
rect 22560 16507 22612 16516
rect 22560 16473 22569 16507
rect 22569 16473 22603 16507
rect 22603 16473 22612 16507
rect 22560 16464 22612 16473
rect 25872 16532 25924 16584
rect 32128 16532 32180 16584
rect 33324 16532 33376 16584
rect 24860 16464 24912 16516
rect 22928 16439 22980 16448
rect 22928 16405 22937 16439
rect 22937 16405 22971 16439
rect 22971 16405 22980 16439
rect 22928 16396 22980 16405
rect 30380 16396 30432 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1492 16167 1544 16176
rect 1492 16133 1501 16167
rect 1501 16133 1535 16167
rect 1535 16133 1544 16167
rect 1492 16124 1544 16133
rect 3976 16099 4028 16108
rect 3976 16065 3985 16099
rect 3985 16065 4019 16099
rect 4019 16065 4028 16099
rect 3976 16056 4028 16065
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 4528 16099 4580 16108
rect 4528 16065 4537 16099
rect 4537 16065 4571 16099
rect 4571 16065 4580 16099
rect 4528 16056 4580 16065
rect 6184 16192 6236 16244
rect 7196 16192 7248 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 8576 16192 8628 16244
rect 940 15852 992 15904
rect 4712 15920 4764 15972
rect 6828 16124 6880 16176
rect 9128 16056 9180 16108
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 8484 15920 8536 15972
rect 8760 15920 8812 15972
rect 9036 15963 9088 15972
rect 9036 15929 9045 15963
rect 9045 15929 9079 15963
rect 9079 15929 9088 15963
rect 9036 15920 9088 15929
rect 9128 15920 9180 15972
rect 12164 16124 12216 16176
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 13912 16167 13964 16176
rect 13912 16133 13921 16167
rect 13921 16133 13955 16167
rect 13955 16133 13964 16167
rect 13912 16124 13964 16133
rect 18880 16192 18932 16244
rect 30104 16235 30156 16244
rect 30104 16201 30113 16235
rect 30113 16201 30147 16235
rect 30147 16201 30156 16235
rect 30104 16192 30156 16201
rect 34336 16235 34388 16244
rect 34336 16201 34345 16235
rect 34345 16201 34379 16235
rect 34379 16201 34388 16235
rect 34336 16192 34388 16201
rect 16948 16167 17000 16176
rect 16948 16133 16957 16167
rect 16957 16133 16991 16167
rect 16991 16133 17000 16167
rect 16948 16124 17000 16133
rect 12808 15988 12860 16040
rect 13084 16031 13136 16040
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 16028 15988 16080 16040
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 16212 15852 16264 15861
rect 16856 15920 16908 15972
rect 17500 16056 17552 16108
rect 17684 16056 17736 16108
rect 17776 16099 17828 16108
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 17868 16056 17920 16108
rect 18972 16099 19024 16108
rect 18972 16065 18981 16099
rect 18981 16065 19015 16099
rect 19015 16065 19024 16099
rect 18972 16056 19024 16065
rect 20628 16124 20680 16176
rect 20444 16056 20496 16108
rect 20904 16056 20956 16108
rect 24308 16099 24360 16108
rect 24308 16065 24317 16099
rect 24317 16065 24351 16099
rect 24351 16065 24360 16099
rect 24308 16056 24360 16065
rect 24584 16056 24636 16108
rect 24952 16056 25004 16108
rect 25136 16056 25188 16108
rect 27160 16124 27212 16176
rect 29368 16167 29420 16176
rect 29368 16133 29377 16167
rect 29377 16133 29411 16167
rect 29411 16133 29420 16167
rect 29368 16124 29420 16133
rect 29092 16056 29144 16108
rect 30288 16056 30340 16108
rect 26240 15988 26292 16040
rect 26424 15988 26476 16040
rect 32864 16056 32916 16108
rect 33968 16099 34020 16108
rect 33968 16065 33977 16099
rect 33977 16065 34011 16099
rect 34011 16065 34020 16099
rect 33968 16056 34020 16065
rect 37648 16099 37700 16108
rect 37648 16065 37657 16099
rect 37657 16065 37691 16099
rect 37691 16065 37700 16099
rect 37648 16056 37700 16065
rect 33876 16031 33928 16040
rect 33876 15997 33885 16031
rect 33885 15997 33919 16031
rect 33919 15997 33928 16031
rect 33876 15988 33928 15997
rect 20628 15920 20680 15972
rect 26516 15920 26568 15972
rect 26884 15920 26936 15972
rect 27896 15920 27948 15972
rect 30380 15920 30432 15972
rect 30748 15920 30800 15972
rect 18696 15852 18748 15904
rect 24676 15852 24728 15904
rect 27160 15852 27212 15904
rect 29552 15895 29604 15904
rect 29552 15861 29561 15895
rect 29561 15861 29595 15895
rect 29595 15861 29604 15895
rect 29552 15852 29604 15861
rect 29828 15852 29880 15904
rect 37832 15895 37884 15904
rect 37832 15861 37841 15895
rect 37841 15861 37875 15895
rect 37875 15861 37884 15895
rect 37832 15852 37884 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2964 15648 3016 15700
rect 3976 15648 4028 15700
rect 4712 15648 4764 15700
rect 6736 15648 6788 15700
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 4620 15512 4672 15564
rect 2780 15444 2832 15496
rect 9588 15648 9640 15700
rect 14556 15648 14608 15700
rect 14740 15648 14792 15700
rect 17132 15648 17184 15700
rect 17408 15648 17460 15700
rect 17776 15648 17828 15700
rect 18052 15648 18104 15700
rect 20904 15648 20956 15700
rect 21548 15648 21600 15700
rect 12992 15580 13044 15632
rect 22560 15648 22612 15700
rect 25136 15648 25188 15700
rect 9312 15512 9364 15564
rect 6920 15444 6972 15496
rect 8760 15487 8812 15496
rect 8760 15453 8769 15487
rect 8769 15453 8803 15487
rect 8803 15453 8812 15487
rect 8760 15444 8812 15453
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 1676 15419 1728 15428
rect 1676 15385 1685 15419
rect 1685 15385 1719 15419
rect 1719 15385 1728 15419
rect 1676 15376 1728 15385
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 9956 15308 10008 15360
rect 11336 15419 11388 15428
rect 11336 15385 11345 15419
rect 11345 15385 11379 15419
rect 11379 15385 11388 15419
rect 11336 15376 11388 15385
rect 14464 15555 14516 15564
rect 14464 15521 14473 15555
rect 14473 15521 14507 15555
rect 14507 15521 14516 15555
rect 14464 15512 14516 15521
rect 14740 15512 14792 15564
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 13268 15444 13320 15496
rect 16212 15512 16264 15564
rect 16488 15512 16540 15564
rect 24400 15580 24452 15632
rect 26424 15580 26476 15632
rect 13084 15376 13136 15428
rect 11980 15308 12032 15360
rect 12900 15308 12952 15360
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 18880 15512 18932 15564
rect 20996 15512 21048 15564
rect 14372 15308 14424 15360
rect 15660 15308 15712 15360
rect 15844 15308 15896 15360
rect 16856 15444 16908 15496
rect 18052 15444 18104 15496
rect 18972 15444 19024 15496
rect 20444 15487 20496 15496
rect 20444 15453 20453 15487
rect 20453 15453 20487 15487
rect 20487 15453 20496 15487
rect 20444 15444 20496 15453
rect 20628 15444 20680 15496
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 21916 15512 21968 15564
rect 26884 15623 26936 15632
rect 26884 15589 26893 15623
rect 26893 15589 26927 15623
rect 26927 15589 26936 15623
rect 26884 15580 26936 15589
rect 27160 15580 27212 15632
rect 21272 15444 21324 15496
rect 16120 15419 16172 15428
rect 16120 15385 16129 15419
rect 16129 15385 16163 15419
rect 16163 15385 16172 15419
rect 16120 15376 16172 15385
rect 16304 15376 16356 15428
rect 17776 15376 17828 15428
rect 16580 15308 16632 15360
rect 17316 15351 17368 15360
rect 17316 15317 17341 15351
rect 17341 15317 17368 15351
rect 17316 15308 17368 15317
rect 20720 15351 20772 15360
rect 20720 15317 20729 15351
rect 20729 15317 20763 15351
rect 20763 15317 20772 15351
rect 20720 15308 20772 15317
rect 22284 15419 22336 15428
rect 22284 15385 22293 15419
rect 22293 15385 22327 15419
rect 22327 15385 22336 15419
rect 22284 15376 22336 15385
rect 23204 15487 23256 15496
rect 23204 15453 23213 15487
rect 23213 15453 23247 15487
rect 23247 15453 23256 15487
rect 23204 15444 23256 15453
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 23572 15444 23624 15496
rect 24676 15444 24728 15496
rect 24952 15444 25004 15496
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 26332 15444 26384 15496
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 29552 15648 29604 15700
rect 30656 15648 30708 15700
rect 28172 15512 28224 15564
rect 30380 15623 30432 15632
rect 30380 15589 30389 15623
rect 30389 15589 30423 15623
rect 30423 15589 30432 15623
rect 30380 15580 30432 15589
rect 30748 15512 30800 15564
rect 23940 15308 23992 15360
rect 26240 15376 26292 15428
rect 27712 15376 27764 15428
rect 27896 15444 27948 15496
rect 29092 15444 29144 15496
rect 29828 15444 29880 15496
rect 32036 15555 32088 15564
rect 32036 15521 32045 15555
rect 32045 15521 32079 15555
rect 32079 15521 32088 15555
rect 32036 15512 32088 15521
rect 28908 15376 28960 15428
rect 27804 15308 27856 15360
rect 27988 15308 28040 15360
rect 28724 15351 28776 15360
rect 28724 15317 28733 15351
rect 28733 15317 28767 15351
rect 28767 15317 28776 15351
rect 28724 15308 28776 15317
rect 30104 15351 30156 15360
rect 30104 15317 30113 15351
rect 30113 15317 30147 15351
rect 30147 15317 30156 15351
rect 30104 15308 30156 15317
rect 32404 15444 32456 15496
rect 33876 15648 33928 15700
rect 32956 15308 33008 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1676 15104 1728 15156
rect 2964 15147 3016 15156
rect 2964 15113 2973 15147
rect 2973 15113 3007 15147
rect 3007 15113 3016 15147
rect 2964 15104 3016 15113
rect 3792 15104 3844 15156
rect 6828 15104 6880 15156
rect 7380 15104 7432 15156
rect 8760 15104 8812 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 11336 15104 11388 15156
rect 6920 15036 6972 15088
rect 8300 15036 8352 15088
rect 9312 15036 9364 15088
rect 3884 14968 3936 15020
rect 3056 14900 3108 14952
rect 4712 14968 4764 15020
rect 6368 15011 6420 15020
rect 6368 14977 6377 15011
rect 6377 14977 6411 15011
rect 6411 14977 6420 15011
rect 6368 14968 6420 14977
rect 9404 14968 9456 15020
rect 11796 15104 11848 15156
rect 12992 15104 13044 15156
rect 16120 15104 16172 15156
rect 16212 15147 16264 15156
rect 16212 15113 16221 15147
rect 16221 15113 16255 15147
rect 16255 15113 16264 15147
rect 16212 15104 16264 15113
rect 16396 15104 16448 15156
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 13268 14968 13320 15020
rect 14832 14968 14884 15020
rect 15660 15036 15712 15088
rect 15752 14968 15804 15020
rect 6644 14943 6696 14952
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 6644 14900 6696 14909
rect 11336 14900 11388 14952
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 12532 14900 12584 14952
rect 18236 15104 18288 15156
rect 20168 15147 20220 15156
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 17040 15036 17092 15088
rect 17500 15036 17552 15088
rect 16948 14968 17000 15020
rect 17868 14968 17920 15020
rect 19984 15036 20036 15088
rect 18052 14968 18104 15020
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 7656 14832 7708 14884
rect 9864 14832 9916 14884
rect 17224 14900 17276 14952
rect 18236 14900 18288 14952
rect 15384 14832 15436 14884
rect 16672 14832 16724 14884
rect 20444 14968 20496 15020
rect 20720 15036 20772 15088
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 24308 15104 24360 15156
rect 25504 15104 25556 15156
rect 26976 15104 27028 15156
rect 27068 15104 27120 15156
rect 23388 15011 23440 15020
rect 23388 14977 23397 15011
rect 23397 14977 23431 15011
rect 23431 14977 23440 15011
rect 23388 14968 23440 14977
rect 24584 15011 24636 15020
rect 24584 14977 24593 15011
rect 24593 14977 24627 15011
rect 24627 14977 24636 15011
rect 24584 14968 24636 14977
rect 26240 15079 26292 15088
rect 26240 15045 26249 15079
rect 26249 15045 26283 15079
rect 26283 15045 26292 15079
rect 26240 15036 26292 15045
rect 26516 15036 26568 15088
rect 27988 15036 28040 15088
rect 28356 15036 28408 15088
rect 23480 14900 23532 14952
rect 24124 14900 24176 14952
rect 25872 14900 25924 14952
rect 27896 15011 27948 15020
rect 27896 14977 27905 15011
rect 27905 14977 27939 15011
rect 27939 14977 27948 15011
rect 27896 14968 27948 14977
rect 28264 15011 28316 15020
rect 28264 14977 28273 15011
rect 28273 14977 28307 15011
rect 28307 14977 28316 15011
rect 28264 14968 28316 14977
rect 30656 15036 30708 15088
rect 5448 14764 5500 14816
rect 7288 14764 7340 14816
rect 15016 14807 15068 14816
rect 15016 14773 15025 14807
rect 15025 14773 15059 14807
rect 15059 14773 15068 14807
rect 15016 14764 15068 14773
rect 15200 14764 15252 14816
rect 16488 14764 16540 14816
rect 20168 14832 20220 14884
rect 20996 14832 21048 14884
rect 25044 14832 25096 14884
rect 18328 14764 18380 14816
rect 19616 14764 19668 14816
rect 20260 14764 20312 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 21088 14764 21140 14816
rect 25596 14807 25648 14816
rect 25596 14773 25605 14807
rect 25605 14773 25639 14807
rect 25639 14773 25648 14807
rect 25596 14764 25648 14773
rect 25780 14807 25832 14816
rect 25780 14773 25789 14807
rect 25789 14773 25823 14807
rect 25823 14773 25832 14807
rect 25780 14764 25832 14773
rect 26700 14807 26752 14816
rect 26700 14773 26709 14807
rect 26709 14773 26743 14807
rect 26743 14773 26752 14807
rect 26700 14764 26752 14773
rect 27988 14875 28040 14884
rect 27988 14841 27997 14875
rect 27997 14841 28031 14875
rect 28031 14841 28040 14875
rect 27988 14832 28040 14841
rect 28632 14943 28684 14952
rect 28632 14909 28641 14943
rect 28641 14909 28675 14943
rect 28675 14909 28684 14943
rect 28632 14900 28684 14909
rect 29092 14968 29144 15020
rect 29368 15011 29420 15020
rect 29368 14977 29377 15011
rect 29377 14977 29411 15011
rect 29411 14977 29420 15011
rect 29368 14968 29420 14977
rect 29552 14900 29604 14952
rect 30012 14900 30064 14952
rect 30564 14968 30616 15020
rect 32864 15036 32916 15088
rect 33048 15079 33100 15088
rect 33048 15045 33057 15079
rect 33057 15045 33091 15079
rect 33091 15045 33100 15079
rect 33048 15036 33100 15045
rect 31760 14968 31812 15020
rect 33416 14968 33468 15020
rect 32956 14900 33008 14952
rect 30288 14832 30340 14884
rect 28632 14764 28684 14816
rect 30932 14764 30984 14816
rect 33232 14807 33284 14816
rect 33232 14773 33241 14807
rect 33241 14773 33275 14807
rect 33275 14773 33284 14807
rect 33232 14764 33284 14773
rect 33600 14807 33652 14816
rect 33600 14773 33609 14807
rect 33609 14773 33643 14807
rect 33643 14773 33652 14807
rect 33600 14764 33652 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 6460 14560 6512 14612
rect 6644 14560 6696 14612
rect 13268 14603 13320 14612
rect 13268 14569 13277 14603
rect 13277 14569 13311 14603
rect 13311 14569 13320 14603
rect 13268 14560 13320 14569
rect 13912 14560 13964 14612
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 15476 14560 15528 14612
rect 16764 14603 16816 14612
rect 16764 14569 16773 14603
rect 16773 14569 16807 14603
rect 16807 14569 16816 14603
rect 16764 14560 16816 14569
rect 19156 14560 19208 14612
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 20076 14603 20128 14612
rect 20076 14569 20085 14603
rect 20085 14569 20119 14603
rect 20119 14569 20128 14603
rect 20076 14560 20128 14569
rect 23388 14560 23440 14612
rect 27252 14560 27304 14612
rect 27988 14560 28040 14612
rect 28172 14603 28224 14612
rect 28172 14569 28181 14603
rect 28181 14569 28215 14603
rect 28215 14569 28224 14603
rect 28172 14560 28224 14569
rect 28356 14560 28408 14612
rect 6828 14492 6880 14544
rect 6368 14424 6420 14476
rect 3792 14356 3844 14408
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 6000 14356 6052 14408
rect 7380 14467 7432 14476
rect 7380 14433 7389 14467
rect 7389 14433 7423 14467
rect 7423 14433 7432 14467
rect 7380 14424 7432 14433
rect 7564 14467 7616 14476
rect 7564 14433 7573 14467
rect 7573 14433 7607 14467
rect 7607 14433 7616 14467
rect 7564 14424 7616 14433
rect 8668 14424 8720 14476
rect 4804 14288 4856 14340
rect 4896 14331 4948 14340
rect 4896 14297 4905 14331
rect 4905 14297 4939 14331
rect 4939 14297 4948 14331
rect 4896 14288 4948 14297
rect 3976 14263 4028 14272
rect 3976 14229 3985 14263
rect 3985 14229 4019 14263
rect 4019 14229 4028 14263
rect 3976 14220 4028 14229
rect 4068 14220 4120 14272
rect 8300 14356 8352 14408
rect 11060 14356 11112 14408
rect 15752 14535 15804 14544
rect 15752 14501 15761 14535
rect 15761 14501 15795 14535
rect 15795 14501 15804 14535
rect 15752 14492 15804 14501
rect 14924 14356 14976 14408
rect 15016 14356 15068 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 11796 14331 11848 14340
rect 11796 14297 11805 14331
rect 11805 14297 11839 14331
rect 11839 14297 11848 14331
rect 11796 14288 11848 14297
rect 13084 14288 13136 14340
rect 13452 14288 13504 14340
rect 10140 14220 10192 14272
rect 11704 14220 11756 14272
rect 12440 14220 12492 14272
rect 14832 14263 14884 14272
rect 14832 14229 14841 14263
rect 14841 14229 14875 14263
rect 14875 14229 14884 14263
rect 14832 14220 14884 14229
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 16580 14424 16632 14476
rect 20720 14492 20772 14544
rect 16212 14356 16264 14408
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 17684 14424 17736 14476
rect 18788 14424 18840 14476
rect 19064 14424 19116 14476
rect 17224 14356 17276 14408
rect 15844 14288 15896 14340
rect 17868 14356 17920 14408
rect 15936 14220 15988 14272
rect 16120 14220 16172 14272
rect 17960 14288 18012 14340
rect 18512 14331 18564 14340
rect 18512 14297 18521 14331
rect 18521 14297 18555 14331
rect 18555 14297 18564 14331
rect 18512 14288 18564 14297
rect 18236 14220 18288 14272
rect 19248 14331 19300 14340
rect 19248 14297 19257 14331
rect 19257 14297 19291 14331
rect 19291 14297 19300 14331
rect 19248 14288 19300 14297
rect 20168 14356 20220 14408
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 20904 14424 20956 14476
rect 21180 14467 21232 14476
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 24952 14424 25004 14476
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 22192 14288 22244 14340
rect 24216 14356 24268 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 25044 14356 25096 14408
rect 22744 14220 22796 14272
rect 23480 14220 23532 14272
rect 27988 14288 28040 14340
rect 28172 14288 28224 14340
rect 28724 14356 28776 14408
rect 30656 14492 30708 14544
rect 30840 14356 30892 14408
rect 31484 14399 31536 14408
rect 31484 14365 31493 14399
rect 31493 14365 31527 14399
rect 31527 14365 31536 14399
rect 31484 14356 31536 14365
rect 31576 14399 31628 14408
rect 31576 14365 31585 14399
rect 31585 14365 31619 14399
rect 31619 14365 31628 14399
rect 32036 14560 32088 14612
rect 33048 14560 33100 14612
rect 33324 14603 33376 14612
rect 33324 14569 33333 14603
rect 33333 14569 33367 14603
rect 33367 14569 33376 14603
rect 33324 14560 33376 14569
rect 32956 14424 33008 14476
rect 33600 14424 33652 14476
rect 31576 14356 31628 14365
rect 30472 14220 30524 14272
rect 30748 14331 30800 14340
rect 30748 14297 30757 14331
rect 30757 14297 30791 14331
rect 30791 14297 30800 14331
rect 30748 14288 30800 14297
rect 30932 14331 30984 14340
rect 30932 14297 30941 14331
rect 30941 14297 30975 14331
rect 30975 14297 30984 14331
rect 30932 14288 30984 14297
rect 31300 14288 31352 14340
rect 34060 14356 34112 14408
rect 32680 14288 32732 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 3976 14016 4028 14068
rect 4620 14059 4672 14068
rect 4620 14025 4645 14059
rect 4645 14025 4672 14059
rect 4620 14016 4672 14025
rect 4804 14059 4856 14068
rect 4804 14025 4813 14059
rect 4813 14025 4847 14059
rect 4847 14025 4856 14059
rect 4804 14016 4856 14025
rect 4896 14016 4948 14068
rect 3884 13948 3936 14000
rect 2780 13880 2832 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 4068 13812 4120 13864
rect 4528 13812 4580 13864
rect 4804 13812 4856 13864
rect 11152 14016 11204 14068
rect 11704 14016 11756 14068
rect 11796 14016 11848 14068
rect 12532 14016 12584 14068
rect 13360 14016 13412 14068
rect 14832 14016 14884 14068
rect 14924 14059 14976 14068
rect 14924 14025 14939 14059
rect 14939 14025 14973 14059
rect 14973 14025 14976 14059
rect 14924 14016 14976 14025
rect 15292 14016 15344 14068
rect 15844 14016 15896 14068
rect 15936 14016 15988 14068
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 2964 13744 3016 13796
rect 6368 13744 6420 13796
rect 9312 13948 9364 14000
rect 9772 13948 9824 14000
rect 9956 13948 10008 14000
rect 10140 13948 10192 14000
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 7564 13812 7616 13864
rect 9036 13812 9088 13864
rect 11888 13880 11940 13932
rect 12440 13880 12492 13932
rect 14740 13880 14792 13932
rect 15016 13923 15068 13932
rect 15016 13889 15025 13923
rect 15025 13889 15059 13923
rect 15059 13889 15068 13923
rect 15016 13880 15068 13889
rect 11336 13812 11388 13864
rect 15476 13880 15528 13932
rect 16120 13923 16172 13932
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 16120 13880 16172 13889
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 17960 14016 18012 14068
rect 17684 13880 17736 13932
rect 17776 13923 17828 13932
rect 17776 13889 17785 13923
rect 17785 13889 17819 13923
rect 17819 13889 17828 13923
rect 17776 13880 17828 13889
rect 16580 13812 16632 13864
rect 18328 13923 18380 13932
rect 18328 13889 18337 13923
rect 18337 13889 18371 13923
rect 18371 13889 18380 13923
rect 18328 13880 18380 13889
rect 18788 14059 18840 14068
rect 18788 14025 18797 14059
rect 18797 14025 18831 14059
rect 18831 14025 18840 14059
rect 18788 14016 18840 14025
rect 19248 14016 19300 14068
rect 20536 14016 20588 14068
rect 22192 14016 22244 14068
rect 23020 14016 23072 14068
rect 24952 14016 25004 14068
rect 25044 14059 25096 14068
rect 25044 14025 25053 14059
rect 25053 14025 25087 14059
rect 25087 14025 25096 14059
rect 25044 14016 25096 14025
rect 25320 14016 25372 14068
rect 25872 14016 25924 14068
rect 28264 14016 28316 14068
rect 28632 14016 28684 14068
rect 18604 13880 18656 13932
rect 18788 13812 18840 13864
rect 18972 13812 19024 13864
rect 2872 13676 2924 13728
rect 4712 13676 4764 13728
rect 8208 13676 8260 13728
rect 8576 13676 8628 13728
rect 17868 13744 17920 13796
rect 19432 13744 19484 13796
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 9588 13676 9640 13728
rect 12072 13676 12124 13728
rect 16028 13676 16080 13728
rect 22008 13948 22060 14000
rect 20904 13880 20956 13932
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 22836 13991 22888 14000
rect 22836 13957 22845 13991
rect 22845 13957 22879 13991
rect 22879 13957 22888 13991
rect 22836 13948 22888 13957
rect 22560 13812 22612 13864
rect 22744 13676 22796 13728
rect 23388 13744 23440 13796
rect 23664 13880 23716 13932
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24860 13880 24912 13932
rect 25136 13880 25188 13932
rect 24124 13812 24176 13864
rect 25504 13923 25556 13932
rect 25504 13889 25513 13923
rect 25513 13889 25547 13923
rect 25547 13889 25556 13923
rect 25504 13880 25556 13889
rect 25688 13923 25740 13932
rect 25688 13889 25697 13923
rect 25697 13889 25731 13923
rect 25731 13889 25740 13923
rect 25688 13880 25740 13889
rect 30748 14016 30800 14068
rect 31576 14016 31628 14068
rect 33324 14016 33376 14068
rect 26700 13880 26752 13932
rect 26884 13880 26936 13932
rect 28172 13880 28224 13932
rect 23664 13719 23716 13728
rect 23664 13685 23673 13719
rect 23673 13685 23707 13719
rect 23707 13685 23716 13719
rect 23664 13676 23716 13685
rect 24032 13676 24084 13728
rect 25872 13744 25924 13796
rect 28632 13923 28684 13932
rect 28632 13889 28641 13923
rect 28641 13889 28675 13923
rect 28675 13889 28684 13923
rect 28632 13880 28684 13889
rect 31852 13880 31904 13932
rect 33140 13923 33192 13932
rect 33140 13889 33149 13923
rect 33149 13889 33183 13923
rect 33183 13889 33192 13923
rect 33140 13880 33192 13889
rect 33232 13880 33284 13932
rect 33876 13948 33928 14000
rect 30564 13812 30616 13864
rect 31760 13812 31812 13864
rect 32588 13812 32640 13864
rect 33784 13880 33836 13932
rect 33968 13880 34020 13932
rect 25964 13676 26016 13728
rect 26240 13719 26292 13728
rect 26240 13685 26249 13719
rect 26249 13685 26283 13719
rect 26283 13685 26292 13719
rect 26240 13676 26292 13685
rect 27252 13676 27304 13728
rect 28540 13744 28592 13796
rect 29920 13744 29972 13796
rect 31668 13676 31720 13728
rect 32956 13676 33008 13728
rect 33600 13676 33652 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 940 13472 992 13524
rect 1676 13472 1728 13524
rect 3792 13515 3844 13524
rect 3792 13481 3801 13515
rect 3801 13481 3835 13515
rect 3835 13481 3844 13515
rect 3792 13472 3844 13481
rect 6368 13472 6420 13524
rect 6828 13472 6880 13524
rect 8208 13515 8260 13524
rect 8208 13481 8217 13515
rect 8217 13481 8251 13515
rect 8251 13481 8260 13515
rect 8208 13472 8260 13481
rect 9588 13472 9640 13524
rect 2964 13379 3016 13388
rect 2964 13345 2973 13379
rect 2973 13345 3007 13379
rect 3007 13345 3016 13379
rect 2964 13336 3016 13345
rect 3056 13379 3108 13388
rect 3056 13345 3065 13379
rect 3065 13345 3099 13379
rect 3099 13345 3108 13379
rect 3056 13336 3108 13345
rect 3884 13268 3936 13320
rect 4712 13268 4764 13320
rect 10324 13472 10376 13524
rect 11152 13472 11204 13524
rect 12532 13472 12584 13524
rect 14556 13472 14608 13524
rect 15016 13472 15068 13524
rect 18328 13472 18380 13524
rect 20444 13472 20496 13524
rect 20720 13472 20772 13524
rect 22560 13472 22612 13524
rect 23204 13472 23256 13524
rect 9864 13336 9916 13388
rect 10048 13336 10100 13388
rect 10416 13336 10468 13388
rect 12808 13336 12860 13388
rect 13360 13336 13412 13388
rect 7840 13200 7892 13252
rect 9128 13200 9180 13252
rect 9496 13200 9548 13252
rect 12532 13200 12584 13252
rect 3056 13132 3108 13184
rect 4620 13132 4672 13184
rect 6736 13132 6788 13184
rect 8668 13132 8720 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 9588 13132 9640 13184
rect 12440 13132 12492 13184
rect 13176 13268 13228 13320
rect 14556 13268 14608 13320
rect 15016 13268 15068 13320
rect 15476 13404 15528 13456
rect 16672 13404 16724 13456
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15660 13268 15712 13320
rect 16764 13268 16816 13320
rect 17500 13268 17552 13320
rect 22100 13404 22152 13456
rect 25504 13472 25556 13524
rect 27252 13472 27304 13524
rect 24860 13404 24912 13456
rect 27896 13472 27948 13524
rect 18696 13336 18748 13388
rect 20168 13336 20220 13388
rect 20812 13336 20864 13388
rect 20352 13200 20404 13252
rect 20720 13268 20772 13320
rect 20996 13243 21048 13252
rect 20996 13209 21005 13243
rect 21005 13209 21039 13243
rect 21039 13209 21048 13243
rect 20996 13200 21048 13209
rect 21180 13243 21232 13252
rect 21180 13209 21205 13243
rect 21205 13209 21232 13243
rect 21180 13200 21232 13209
rect 22192 13268 22244 13320
rect 22376 13311 22428 13320
rect 22376 13277 22385 13311
rect 22385 13277 22419 13311
rect 22419 13277 22428 13311
rect 22376 13268 22428 13277
rect 21732 13132 21784 13184
rect 21824 13132 21876 13184
rect 23112 13200 23164 13252
rect 23388 13311 23440 13320
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 23480 13311 23532 13320
rect 23480 13277 23489 13311
rect 23489 13277 23523 13311
rect 23523 13277 23532 13311
rect 23480 13268 23532 13277
rect 23664 13268 23716 13320
rect 23756 13200 23808 13252
rect 23388 13132 23440 13184
rect 25044 13268 25096 13320
rect 25780 13311 25832 13320
rect 25780 13277 25789 13311
rect 25789 13277 25823 13311
rect 25823 13277 25832 13311
rect 25780 13268 25832 13277
rect 25964 13268 26016 13320
rect 26240 13311 26292 13320
rect 26240 13277 26249 13311
rect 26249 13277 26283 13311
rect 26283 13277 26292 13311
rect 26240 13268 26292 13277
rect 26424 13311 26476 13320
rect 26424 13277 26433 13311
rect 26433 13277 26467 13311
rect 26467 13277 26476 13311
rect 26424 13268 26476 13277
rect 26516 13268 26568 13320
rect 26976 13268 27028 13320
rect 26792 13243 26844 13252
rect 26792 13209 26801 13243
rect 26801 13209 26835 13243
rect 26835 13209 26844 13243
rect 26792 13200 26844 13209
rect 25872 13132 25924 13184
rect 26332 13132 26384 13184
rect 27252 13268 27304 13320
rect 28632 13404 28684 13456
rect 30104 13472 30156 13524
rect 31944 13515 31996 13524
rect 31944 13481 31953 13515
rect 31953 13481 31987 13515
rect 31987 13481 31996 13515
rect 31944 13472 31996 13481
rect 32128 13515 32180 13524
rect 32128 13481 32137 13515
rect 32137 13481 32171 13515
rect 32171 13481 32180 13515
rect 32128 13472 32180 13481
rect 33692 13472 33744 13524
rect 29828 13404 29880 13456
rect 28448 13311 28500 13320
rect 28448 13277 28457 13311
rect 28457 13277 28491 13311
rect 28491 13277 28500 13311
rect 28448 13268 28500 13277
rect 28540 13311 28592 13320
rect 28540 13277 28549 13311
rect 28549 13277 28583 13311
rect 28583 13277 28592 13311
rect 28540 13268 28592 13277
rect 29000 13268 29052 13320
rect 27528 13132 27580 13184
rect 29000 13132 29052 13184
rect 29368 13175 29420 13184
rect 29368 13141 29377 13175
rect 29377 13141 29411 13175
rect 29411 13141 29420 13175
rect 29368 13132 29420 13141
rect 29644 13200 29696 13252
rect 30656 13311 30708 13320
rect 30656 13277 30665 13311
rect 30665 13277 30699 13311
rect 30699 13277 30708 13311
rect 30656 13268 30708 13277
rect 31760 13336 31812 13388
rect 30104 13200 30156 13252
rect 30380 13200 30432 13252
rect 31668 13268 31720 13320
rect 32956 13311 33008 13320
rect 32956 13277 32965 13311
rect 32965 13277 32999 13311
rect 32999 13277 33008 13311
rect 32956 13268 33008 13277
rect 33508 13311 33560 13320
rect 33508 13277 33517 13311
rect 33517 13277 33551 13311
rect 33551 13277 33560 13311
rect 33508 13268 33560 13277
rect 33048 13200 33100 13252
rect 33324 13243 33376 13252
rect 33324 13209 33333 13243
rect 33333 13209 33367 13243
rect 33367 13209 33376 13243
rect 33324 13200 33376 13209
rect 33784 13268 33836 13320
rect 33876 13311 33928 13320
rect 33876 13277 33885 13311
rect 33885 13277 33919 13311
rect 33919 13277 33928 13311
rect 33876 13268 33928 13277
rect 30472 13132 30524 13184
rect 30840 13132 30892 13184
rect 33600 13132 33652 13184
rect 34244 13175 34296 13184
rect 34244 13141 34253 13175
rect 34253 13141 34287 13175
rect 34287 13141 34296 13175
rect 34244 13132 34296 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 2872 12928 2924 12980
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 3884 12792 3936 12844
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 4804 12860 4856 12912
rect 5172 12860 5224 12912
rect 4620 12724 4672 12776
rect 6552 12928 6604 12980
rect 7196 12928 7248 12980
rect 9220 12928 9272 12980
rect 8760 12903 8812 12912
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 8760 12860 8812 12869
rect 8208 12792 8260 12844
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 10416 12792 10468 12844
rect 10876 12928 10928 12980
rect 11980 12928 12032 12980
rect 12256 12928 12308 12980
rect 15016 12928 15068 12980
rect 16120 12928 16172 12980
rect 18144 12928 18196 12980
rect 8668 12724 8720 12776
rect 9312 12724 9364 12776
rect 9588 12724 9640 12776
rect 14096 12860 14148 12912
rect 16028 12903 16080 12912
rect 16028 12869 16037 12903
rect 16037 12869 16071 12903
rect 16071 12869 16080 12903
rect 16028 12860 16080 12869
rect 11336 12792 11388 12844
rect 12348 12792 12400 12844
rect 14924 12792 14976 12844
rect 16856 12792 16908 12844
rect 17500 12792 17552 12844
rect 18604 12860 18656 12912
rect 13636 12724 13688 12776
rect 15384 12724 15436 12776
rect 15568 12724 15620 12776
rect 9036 12656 9088 12708
rect 12256 12656 12308 12708
rect 3884 12631 3936 12640
rect 3884 12597 3893 12631
rect 3893 12597 3927 12631
rect 3927 12597 3936 12631
rect 3884 12588 3936 12597
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 8392 12588 8444 12640
rect 10416 12588 10468 12640
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 17776 12724 17828 12776
rect 15752 12656 15804 12708
rect 18328 12792 18380 12844
rect 19064 12792 19116 12844
rect 20812 12792 20864 12844
rect 20996 12860 21048 12912
rect 23020 12928 23072 12980
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 25136 12928 25188 12980
rect 25596 12928 25648 12980
rect 20904 12656 20956 12708
rect 22468 12792 22520 12844
rect 21732 12724 21784 12776
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22100 12724 22152 12733
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 22376 12767 22428 12776
rect 22376 12733 22385 12767
rect 22385 12733 22419 12767
rect 22419 12733 22428 12767
rect 22376 12724 22428 12733
rect 22744 12656 22796 12708
rect 23756 12656 23808 12708
rect 24584 12860 24636 12912
rect 25688 12860 25740 12912
rect 24400 12792 24452 12844
rect 25320 12792 25372 12844
rect 26332 12835 26384 12844
rect 26332 12801 26341 12835
rect 26341 12801 26375 12835
rect 26375 12801 26384 12835
rect 26332 12792 26384 12801
rect 26792 12928 26844 12980
rect 28632 12928 28684 12980
rect 26608 12792 26660 12844
rect 26976 12792 27028 12844
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 28908 12860 28960 12912
rect 31484 12928 31536 12980
rect 33048 12971 33100 12980
rect 33048 12937 33057 12971
rect 33057 12937 33091 12971
rect 33091 12937 33100 12971
rect 33048 12928 33100 12937
rect 33140 12928 33192 12980
rect 33508 12928 33560 12980
rect 34244 12928 34296 12980
rect 24860 12724 24912 12776
rect 25044 12724 25096 12776
rect 26332 12656 26384 12708
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 29092 12792 29144 12844
rect 29276 12835 29328 12844
rect 29276 12801 29285 12835
rect 29285 12801 29319 12835
rect 29319 12801 29328 12835
rect 29276 12792 29328 12801
rect 29000 12724 29052 12776
rect 30564 12792 30616 12844
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 21088 12631 21140 12640
rect 21088 12597 21097 12631
rect 21097 12597 21131 12631
rect 21131 12597 21140 12631
rect 21088 12588 21140 12597
rect 22652 12588 22704 12640
rect 24492 12588 24544 12640
rect 25688 12588 25740 12640
rect 26608 12588 26660 12640
rect 29644 12656 29696 12708
rect 29828 12656 29880 12708
rect 31484 12835 31536 12844
rect 31484 12801 31493 12835
rect 31493 12801 31527 12835
rect 31527 12801 31536 12835
rect 33324 12860 33376 12912
rect 31484 12792 31536 12801
rect 31760 12724 31812 12776
rect 32956 12835 33008 12844
rect 32956 12801 32965 12835
rect 32965 12801 32999 12835
rect 32999 12801 33008 12835
rect 32956 12792 33008 12801
rect 32496 12724 32548 12776
rect 33968 12835 34020 12844
rect 33968 12801 33977 12835
rect 33977 12801 34011 12835
rect 34011 12801 34020 12835
rect 33968 12792 34020 12801
rect 30472 12656 30524 12708
rect 29552 12588 29604 12640
rect 30380 12588 30432 12640
rect 31944 12699 31996 12708
rect 31944 12665 31953 12699
rect 31953 12665 31987 12699
rect 31987 12665 31996 12699
rect 31944 12656 31996 12665
rect 34336 12656 34388 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 8852 12384 8904 12436
rect 11612 12384 11664 12436
rect 15108 12384 15160 12436
rect 19340 12384 19392 12436
rect 1400 12316 1452 12368
rect 3240 12248 3292 12300
rect 3792 12248 3844 12300
rect 8024 12316 8076 12368
rect 9404 12316 9456 12368
rect 6092 12248 6144 12300
rect 6828 12248 6880 12300
rect 11060 12248 11112 12300
rect 11980 12248 12032 12300
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 3884 12180 3936 12232
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 2780 12112 2832 12164
rect 3424 12112 3476 12164
rect 5724 12112 5776 12164
rect 7380 12112 7432 12164
rect 8760 12180 8812 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 13268 12248 13320 12300
rect 15200 12248 15252 12300
rect 15568 12291 15620 12300
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 18788 12248 18840 12300
rect 19524 12316 19576 12368
rect 20168 12316 20220 12368
rect 22468 12384 22520 12436
rect 12808 12180 12860 12232
rect 18144 12223 18196 12232
rect 8668 12044 8720 12096
rect 10508 12155 10560 12164
rect 10508 12121 10517 12155
rect 10517 12121 10551 12155
rect 10551 12121 10560 12155
rect 10508 12112 10560 12121
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 9496 12044 9548 12096
rect 11520 12044 11572 12096
rect 16212 12155 16264 12164
rect 16212 12121 16221 12155
rect 16221 12121 16255 12155
rect 16255 12121 16264 12155
rect 16212 12112 16264 12121
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 12900 12044 12952 12053
rect 15200 12044 15252 12096
rect 15292 12087 15344 12096
rect 15292 12053 15301 12087
rect 15301 12053 15335 12087
rect 15335 12053 15344 12087
rect 15292 12044 15344 12053
rect 15568 12044 15620 12096
rect 19340 12112 19392 12164
rect 19432 12155 19484 12164
rect 19432 12121 19462 12155
rect 19462 12121 19484 12155
rect 21824 12248 21876 12300
rect 22652 12316 22704 12368
rect 22376 12248 22428 12300
rect 23296 12316 23348 12368
rect 24032 12384 24084 12436
rect 24400 12427 24452 12436
rect 24400 12393 24409 12427
rect 24409 12393 24443 12427
rect 24443 12393 24452 12427
rect 24400 12384 24452 12393
rect 23572 12291 23624 12300
rect 23572 12257 23581 12291
rect 23581 12257 23615 12291
rect 23615 12257 23624 12291
rect 23572 12248 23624 12257
rect 27620 12384 27672 12436
rect 28816 12384 28868 12436
rect 29460 12384 29512 12436
rect 29552 12427 29604 12436
rect 29552 12393 29561 12427
rect 29561 12393 29595 12427
rect 29595 12393 29604 12427
rect 29552 12384 29604 12393
rect 30196 12384 30248 12436
rect 29000 12316 29052 12368
rect 25136 12291 25188 12300
rect 25136 12257 25145 12291
rect 25145 12257 25179 12291
rect 25179 12257 25188 12291
rect 25136 12248 25188 12257
rect 25320 12291 25372 12300
rect 25320 12257 25329 12291
rect 25329 12257 25363 12291
rect 25363 12257 25372 12291
rect 25320 12248 25372 12257
rect 25872 12248 25924 12300
rect 26700 12248 26752 12300
rect 26884 12248 26936 12300
rect 27988 12248 28040 12300
rect 30012 12316 30064 12368
rect 30472 12316 30524 12368
rect 23204 12180 23256 12232
rect 23388 12180 23440 12232
rect 24308 12180 24360 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 19432 12112 19484 12121
rect 22468 12112 22520 12164
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 18696 12044 18748 12096
rect 20076 12087 20128 12096
rect 20076 12053 20085 12087
rect 20085 12053 20119 12087
rect 20119 12053 20128 12087
rect 20076 12044 20128 12053
rect 21456 12044 21508 12096
rect 21824 12087 21876 12096
rect 21824 12053 21849 12087
rect 21849 12053 21876 12087
rect 21824 12044 21876 12053
rect 22560 12044 22612 12096
rect 22928 12044 22980 12096
rect 24860 12112 24912 12164
rect 25688 12180 25740 12232
rect 26332 12180 26384 12232
rect 28908 12223 28960 12232
rect 28908 12189 28917 12223
rect 28917 12189 28951 12223
rect 28951 12189 28960 12223
rect 28908 12180 28960 12189
rect 25964 12112 26016 12164
rect 29460 12180 29512 12232
rect 30196 12223 30248 12232
rect 30196 12189 30205 12223
rect 30205 12189 30239 12223
rect 30239 12189 30248 12223
rect 30196 12180 30248 12189
rect 30564 12223 30616 12232
rect 30564 12189 30573 12223
rect 30573 12189 30607 12223
rect 30607 12189 30616 12223
rect 30564 12180 30616 12189
rect 25780 12044 25832 12096
rect 26700 12087 26752 12096
rect 26700 12053 26709 12087
rect 26709 12053 26743 12087
rect 26743 12053 26752 12087
rect 26700 12044 26752 12053
rect 29276 12044 29328 12096
rect 29828 12044 29880 12096
rect 30104 12087 30156 12096
rect 30104 12053 30113 12087
rect 30113 12053 30147 12087
rect 30147 12053 30156 12087
rect 30104 12044 30156 12053
rect 30656 12087 30708 12096
rect 30656 12053 30665 12087
rect 30665 12053 30699 12087
rect 30699 12053 30708 12087
rect 30656 12044 30708 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 1768 11840 1820 11892
rect 3424 11840 3476 11892
rect 8668 11840 8720 11892
rect 9404 11840 9456 11892
rect 12900 11840 12952 11892
rect 7380 11772 7432 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 2964 11704 3016 11756
rect 3792 11704 3844 11756
rect 6092 11704 6144 11756
rect 6184 11747 6236 11756
rect 6184 11713 6193 11747
rect 6193 11713 6227 11747
rect 6227 11713 6236 11747
rect 6184 11704 6236 11713
rect 9220 11772 9272 11824
rect 9956 11772 10008 11824
rect 12348 11815 12400 11824
rect 12348 11781 12357 11815
rect 12357 11781 12391 11815
rect 12391 11781 12400 11815
rect 12348 11772 12400 11781
rect 13268 11772 13320 11824
rect 15016 11840 15068 11892
rect 15200 11840 15252 11892
rect 16212 11840 16264 11892
rect 14924 11815 14976 11824
rect 14924 11781 14933 11815
rect 14933 11781 14967 11815
rect 14967 11781 14976 11815
rect 14924 11772 14976 11781
rect 8852 11704 8904 11756
rect 9588 11704 9640 11756
rect 11152 11704 11204 11756
rect 12072 11704 12124 11756
rect 17684 11772 17736 11824
rect 21180 11840 21232 11892
rect 21456 11840 21508 11892
rect 24768 11840 24820 11892
rect 25320 11840 25372 11892
rect 25780 11840 25832 11892
rect 7104 11636 7156 11688
rect 8116 11636 8168 11688
rect 9772 11636 9824 11688
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 19616 11747 19668 11756
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 9496 11568 9548 11620
rect 8668 11500 8720 11552
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 8760 11500 8812 11509
rect 8944 11500 8996 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10416 11500 10468 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12256 11500 12308 11552
rect 12808 11500 12860 11552
rect 13912 11636 13964 11688
rect 19984 11704 20036 11756
rect 28632 11840 28684 11892
rect 28908 11840 28960 11892
rect 29276 11840 29328 11892
rect 29828 11840 29880 11892
rect 31208 11840 31260 11892
rect 32956 11883 33008 11892
rect 32956 11849 32965 11883
rect 32965 11849 32999 11883
rect 32999 11849 33008 11883
rect 32956 11840 33008 11849
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 21824 11636 21876 11688
rect 22284 11636 22336 11688
rect 19248 11611 19300 11620
rect 19248 11577 19257 11611
rect 19257 11577 19291 11611
rect 19291 11577 19300 11611
rect 19248 11568 19300 11577
rect 22468 11568 22520 11620
rect 23388 11704 23440 11756
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 24308 11704 24360 11713
rect 24492 11772 24544 11824
rect 24676 11772 24728 11824
rect 26792 11772 26844 11824
rect 26976 11815 27028 11824
rect 26976 11781 26985 11815
rect 26985 11781 27019 11815
rect 27019 11781 27028 11815
rect 26976 11772 27028 11781
rect 27252 11772 27304 11824
rect 26884 11704 26936 11756
rect 27344 11704 27396 11756
rect 24860 11568 24912 11620
rect 25320 11568 25372 11620
rect 14648 11500 14700 11552
rect 15016 11500 15068 11552
rect 15568 11500 15620 11552
rect 17960 11543 18012 11552
rect 17960 11509 17969 11543
rect 17969 11509 18003 11543
rect 18003 11509 18012 11543
rect 17960 11500 18012 11509
rect 19984 11500 20036 11552
rect 22008 11500 22060 11552
rect 22928 11500 22980 11552
rect 27528 11568 27580 11620
rect 27804 11568 27856 11620
rect 29092 11747 29144 11756
rect 29092 11713 29101 11747
rect 29101 11713 29135 11747
rect 29135 11713 29144 11747
rect 29092 11704 29144 11713
rect 29552 11704 29604 11756
rect 26976 11500 27028 11552
rect 27160 11543 27212 11552
rect 27160 11509 27169 11543
rect 27169 11509 27203 11543
rect 27203 11509 27212 11543
rect 27160 11500 27212 11509
rect 28724 11500 28776 11552
rect 30012 11636 30064 11688
rect 31392 11704 31444 11756
rect 30564 11636 30616 11688
rect 30656 11636 30708 11688
rect 31116 11679 31168 11688
rect 31116 11645 31125 11679
rect 31125 11645 31159 11679
rect 31159 11645 31168 11679
rect 31116 11636 31168 11645
rect 33784 11747 33836 11756
rect 33784 11713 33793 11747
rect 33793 11713 33827 11747
rect 33827 11713 33836 11747
rect 33784 11704 33836 11713
rect 33232 11636 33284 11688
rect 30472 11500 30524 11552
rect 32036 11500 32088 11552
rect 33876 11611 33928 11620
rect 33876 11577 33885 11611
rect 33885 11577 33919 11611
rect 33919 11577 33928 11611
rect 33876 11568 33928 11577
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4068 11296 4120 11348
rect 5264 11296 5316 11348
rect 6184 11296 6236 11348
rect 8208 11296 8260 11348
rect 940 11092 992 11144
rect 2780 11160 2832 11212
rect 2964 11024 3016 11076
rect 3884 11160 3936 11212
rect 4436 11092 4488 11144
rect 4528 11092 4580 11144
rect 4712 11092 4764 11144
rect 7104 11203 7156 11212
rect 7104 11169 7113 11203
rect 7113 11169 7147 11203
rect 7147 11169 7156 11203
rect 7104 11160 7156 11169
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 5356 11092 5408 11144
rect 7380 11092 7432 11144
rect 12256 11296 12308 11348
rect 12440 11296 12492 11348
rect 13268 11339 13320 11348
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 9036 11228 9088 11280
rect 12808 11228 12860 11280
rect 15292 11296 15344 11348
rect 20168 11296 20220 11348
rect 8668 11092 8720 11144
rect 9588 11092 9640 11144
rect 10048 11092 10100 11144
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 4620 10956 4672 11008
rect 4712 10999 4764 11008
rect 4712 10965 4721 10999
rect 4721 10965 4755 10999
rect 4755 10965 4764 10999
rect 4712 10956 4764 10965
rect 4896 10956 4948 11008
rect 8668 10956 8720 11008
rect 11060 11092 11112 11144
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 15384 11160 15436 11212
rect 13360 11092 13412 11144
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 12808 11024 12860 11076
rect 13728 11024 13780 11076
rect 14924 11092 14976 11144
rect 15476 11092 15528 11144
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 18052 11092 18104 11144
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 17592 11024 17644 11076
rect 19432 11092 19484 11144
rect 20628 11296 20680 11348
rect 20260 11228 20312 11280
rect 20904 11228 20956 11280
rect 21640 11228 21692 11280
rect 25320 11296 25372 11348
rect 27160 11296 27212 11348
rect 27252 11296 27304 11348
rect 27436 11296 27488 11348
rect 23572 11092 23624 11144
rect 19340 11024 19392 11076
rect 12440 10956 12492 11008
rect 14096 10956 14148 11008
rect 15660 10956 15712 11008
rect 18972 10956 19024 11008
rect 20168 10956 20220 11008
rect 23296 11024 23348 11076
rect 24952 11092 25004 11144
rect 25596 11135 25648 11144
rect 25596 11101 25605 11135
rect 25605 11101 25639 11135
rect 25639 11101 25648 11135
rect 25596 11092 25648 11101
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 25872 11092 25924 11101
rect 26700 11228 26752 11280
rect 26792 11203 26844 11212
rect 26792 11169 26801 11203
rect 26801 11169 26835 11203
rect 26835 11169 26844 11203
rect 26792 11160 26844 11169
rect 27344 11228 27396 11280
rect 27160 11092 27212 11144
rect 27344 11092 27396 11144
rect 27620 11092 27672 11144
rect 29736 11296 29788 11348
rect 31116 11296 31168 11348
rect 32588 11339 32640 11348
rect 32588 11305 32597 11339
rect 32597 11305 32631 11339
rect 32631 11305 32640 11339
rect 32588 11296 32640 11305
rect 28632 11228 28684 11280
rect 33232 11228 33284 11280
rect 32956 11160 33008 11212
rect 23480 10956 23532 11008
rect 23848 10956 23900 11008
rect 24308 10956 24360 11008
rect 25780 11024 25832 11076
rect 25872 10999 25924 11008
rect 25872 10965 25881 10999
rect 25881 10965 25915 10999
rect 25915 10965 25924 10999
rect 25872 10956 25924 10965
rect 26240 10999 26292 11008
rect 26240 10965 26249 10999
rect 26249 10965 26283 10999
rect 26283 10965 26292 10999
rect 26240 10956 26292 10965
rect 27528 10956 27580 11008
rect 27712 10956 27764 11008
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 30564 11092 30616 11144
rect 31392 11092 31444 11144
rect 32036 11135 32088 11144
rect 32036 11101 32045 11135
rect 32045 11101 32079 11135
rect 32079 11101 32088 11135
rect 32036 11092 32088 11101
rect 32312 11135 32364 11144
rect 32312 11101 32321 11135
rect 32321 11101 32355 11135
rect 32355 11101 32364 11135
rect 32312 11092 32364 11101
rect 33140 11092 33192 11144
rect 37280 11092 37332 11144
rect 37924 11067 37976 11076
rect 37924 11033 37933 11067
rect 37933 11033 37967 11067
rect 37967 11033 37976 11067
rect 37924 11024 37976 11033
rect 29828 10956 29880 11008
rect 32588 10956 32640 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3240 10752 3292 10804
rect 4620 10795 4672 10804
rect 4620 10761 4629 10795
rect 4629 10761 4663 10795
rect 4663 10761 4672 10795
rect 4620 10752 4672 10761
rect 4712 10752 4764 10804
rect 10048 10752 10100 10804
rect 1400 10548 1452 10600
rect 3792 10412 3844 10464
rect 5080 10616 5132 10668
rect 5448 10616 5500 10668
rect 4436 10548 4488 10600
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 4896 10480 4948 10532
rect 6092 10548 6144 10600
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 9772 10616 9824 10668
rect 9128 10523 9180 10532
rect 9128 10489 9137 10523
rect 9137 10489 9171 10523
rect 9171 10489 9180 10523
rect 9128 10480 9180 10489
rect 10140 10548 10192 10600
rect 11796 10795 11848 10804
rect 11796 10761 11805 10795
rect 11805 10761 11839 10795
rect 11839 10761 11848 10795
rect 11796 10752 11848 10761
rect 11980 10752 12032 10804
rect 14096 10752 14148 10804
rect 13544 10727 13596 10736
rect 13544 10693 13553 10727
rect 13553 10693 13587 10727
rect 13587 10693 13596 10727
rect 13544 10684 13596 10693
rect 14924 10684 14976 10736
rect 15660 10752 15712 10804
rect 15568 10684 15620 10736
rect 17592 10727 17644 10736
rect 17592 10693 17601 10727
rect 17601 10693 17635 10727
rect 17635 10693 17644 10727
rect 17592 10684 17644 10693
rect 19432 10684 19484 10736
rect 12072 10616 12124 10668
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 13912 10548 13964 10600
rect 14372 10591 14424 10600
rect 14372 10557 14381 10591
rect 14381 10557 14415 10591
rect 14415 10557 14424 10591
rect 14372 10548 14424 10557
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 14648 10616 14700 10668
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 18512 10616 18564 10668
rect 20168 10752 20220 10804
rect 20628 10752 20680 10804
rect 21272 10752 21324 10804
rect 23572 10752 23624 10804
rect 25872 10752 25924 10804
rect 26608 10752 26660 10804
rect 30564 10752 30616 10804
rect 20444 10616 20496 10668
rect 20536 10548 20588 10600
rect 20904 10616 20956 10668
rect 21916 10684 21968 10736
rect 23388 10684 23440 10736
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 21548 10548 21600 10600
rect 5356 10412 5408 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 8760 10412 8812 10464
rect 10140 10412 10192 10464
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 14648 10412 14700 10464
rect 19156 10480 19208 10532
rect 20260 10480 20312 10532
rect 20812 10480 20864 10532
rect 22560 10616 22612 10668
rect 23112 10616 23164 10668
rect 23296 10616 23348 10668
rect 25228 10548 25280 10600
rect 26424 10548 26476 10600
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 27528 10659 27580 10668
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 28448 10616 28500 10668
rect 28540 10659 28592 10668
rect 28540 10625 28549 10659
rect 28549 10625 28583 10659
rect 28583 10625 28592 10659
rect 28540 10616 28592 10625
rect 28724 10616 28776 10668
rect 27252 10591 27304 10600
rect 27252 10557 27261 10591
rect 27261 10557 27295 10591
rect 27295 10557 27304 10591
rect 27252 10548 27304 10557
rect 30472 10616 30524 10668
rect 30748 10659 30800 10668
rect 30748 10625 30757 10659
rect 30757 10625 30791 10659
rect 30791 10625 30800 10659
rect 30748 10616 30800 10625
rect 31944 10616 31996 10668
rect 32312 10616 32364 10668
rect 32496 10616 32548 10668
rect 34888 10795 34940 10804
rect 34888 10761 34897 10795
rect 34897 10761 34931 10795
rect 34931 10761 34940 10795
rect 34888 10752 34940 10761
rect 33876 10684 33928 10736
rect 33692 10616 33744 10668
rect 36544 10659 36596 10668
rect 36544 10625 36553 10659
rect 36553 10625 36587 10659
rect 36587 10625 36596 10659
rect 36544 10616 36596 10625
rect 36636 10616 36688 10668
rect 23572 10480 23624 10532
rect 24860 10480 24912 10532
rect 30656 10548 30708 10600
rect 32588 10591 32640 10600
rect 32588 10557 32597 10591
rect 32597 10557 32631 10591
rect 32631 10557 32640 10591
rect 32588 10548 32640 10557
rect 34612 10591 34664 10600
rect 34612 10557 34621 10591
rect 34621 10557 34655 10591
rect 34655 10557 34664 10591
rect 34612 10548 34664 10557
rect 28632 10480 28684 10532
rect 17316 10412 17368 10464
rect 17868 10412 17920 10464
rect 18420 10412 18472 10464
rect 18788 10412 18840 10464
rect 21640 10412 21692 10464
rect 22376 10455 22428 10464
rect 22376 10421 22385 10455
rect 22385 10421 22419 10455
rect 22419 10421 22428 10455
rect 22376 10412 22428 10421
rect 23756 10455 23808 10464
rect 23756 10421 23765 10455
rect 23765 10421 23799 10455
rect 23799 10421 23808 10455
rect 23756 10412 23808 10421
rect 24216 10412 24268 10464
rect 26884 10412 26936 10464
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 27712 10412 27764 10421
rect 33876 10480 33928 10532
rect 29368 10412 29420 10464
rect 29644 10412 29696 10464
rect 30472 10412 30524 10464
rect 32496 10412 32548 10464
rect 33140 10412 33192 10464
rect 36912 10455 36964 10464
rect 36912 10421 36921 10455
rect 36921 10421 36955 10455
rect 36955 10421 36964 10455
rect 36912 10412 36964 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4620 10251 4672 10260
rect 4620 10217 4629 10251
rect 4629 10217 4663 10251
rect 4663 10217 4672 10251
rect 4620 10208 4672 10217
rect 4804 10208 4856 10260
rect 6368 10208 6420 10260
rect 8668 10208 8720 10260
rect 9128 10208 9180 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 9496 10208 9548 10260
rect 2872 10140 2924 10192
rect 3240 10140 3292 10192
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 3240 10004 3292 10056
rect 6092 10072 6144 10124
rect 6368 10072 6420 10124
rect 7656 10072 7708 10124
rect 8576 10140 8628 10192
rect 4344 10004 4396 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 6276 9936 6328 9988
rect 7380 9936 7432 9988
rect 8392 10115 8444 10124
rect 8392 10081 8401 10115
rect 8401 10081 8435 10115
rect 8435 10081 8444 10115
rect 8392 10072 8444 10081
rect 9036 10072 9088 10124
rect 14188 10208 14240 10260
rect 11060 10072 11112 10124
rect 8760 10004 8812 10056
rect 9128 10004 9180 10056
rect 1492 9868 1544 9920
rect 6920 9868 6972 9920
rect 8852 9936 8904 9988
rect 9036 9936 9088 9988
rect 9312 10004 9364 10056
rect 9588 10004 9640 10056
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 7932 9868 7984 9920
rect 8116 9868 8168 9920
rect 8576 9868 8628 9920
rect 10968 9868 11020 9920
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 12808 9868 12860 9920
rect 13544 9868 13596 9920
rect 14372 10004 14424 10056
rect 14924 10208 14976 10260
rect 14740 10072 14792 10124
rect 15568 10072 15620 10124
rect 16672 10072 16724 10124
rect 14648 10004 14700 10056
rect 17316 10208 17368 10260
rect 17868 10115 17920 10124
rect 17868 10081 17877 10115
rect 17877 10081 17911 10115
rect 17911 10081 17920 10115
rect 17868 10072 17920 10081
rect 17960 10004 18012 10056
rect 18512 10072 18564 10124
rect 18236 10004 18288 10056
rect 14740 9868 14792 9920
rect 15568 9936 15620 9988
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 18788 10047 18840 10056
rect 18788 10013 18798 10047
rect 18798 10013 18832 10047
rect 18832 10013 18840 10047
rect 18788 10004 18840 10013
rect 24492 10208 24544 10260
rect 20260 10140 20312 10192
rect 20812 10140 20864 10192
rect 21088 10183 21140 10192
rect 21088 10149 21097 10183
rect 21097 10149 21131 10183
rect 21131 10149 21140 10183
rect 21088 10140 21140 10149
rect 19248 10115 19300 10124
rect 19248 10081 19257 10115
rect 19257 10081 19291 10115
rect 19291 10081 19300 10115
rect 19248 10072 19300 10081
rect 20628 10115 20680 10124
rect 20628 10081 20637 10115
rect 20637 10081 20671 10115
rect 20671 10081 20680 10115
rect 20628 10072 20680 10081
rect 19892 10004 19944 10056
rect 20444 10004 20496 10056
rect 16120 9868 16172 9920
rect 18236 9868 18288 9920
rect 19432 9868 19484 9920
rect 20260 9868 20312 9920
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 22192 10183 22244 10192
rect 22192 10149 22201 10183
rect 22201 10149 22235 10183
rect 22235 10149 22244 10183
rect 22192 10140 22244 10149
rect 21640 10072 21692 10124
rect 22652 10140 22704 10192
rect 27712 10140 27764 10192
rect 22468 10047 22520 10056
rect 22468 10013 22477 10047
rect 22477 10013 22511 10047
rect 22511 10013 22520 10047
rect 22468 10004 22520 10013
rect 21916 9936 21968 9988
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 23112 10004 23164 10013
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 23756 10004 23808 10056
rect 24124 10004 24176 10056
rect 24584 10004 24636 10056
rect 26240 10004 26292 10056
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 27068 10047 27120 10056
rect 27068 10013 27077 10047
rect 27077 10013 27111 10047
rect 27111 10013 27120 10047
rect 27068 10004 27120 10013
rect 22284 9868 22336 9920
rect 24492 9936 24544 9988
rect 28448 10004 28500 10056
rect 28724 10047 28776 10056
rect 28724 10013 28733 10047
rect 28733 10013 28767 10047
rect 28767 10013 28776 10047
rect 28724 10004 28776 10013
rect 29920 10140 29972 10192
rect 29092 10004 29144 10056
rect 29368 10004 29420 10056
rect 29828 10047 29880 10056
rect 29828 10013 29837 10047
rect 29837 10013 29871 10047
rect 29871 10013 29880 10047
rect 29828 10004 29880 10013
rect 30472 10140 30524 10192
rect 30656 10140 30708 10192
rect 30472 10047 30524 10056
rect 30472 10013 30481 10047
rect 30481 10013 30515 10047
rect 30515 10013 30524 10047
rect 30472 10004 30524 10013
rect 30840 10072 30892 10124
rect 30656 10004 30708 10056
rect 34612 10208 34664 10260
rect 32496 10004 32548 10056
rect 33876 10047 33928 10056
rect 33876 10013 33885 10047
rect 33885 10013 33919 10047
rect 33919 10013 33928 10047
rect 33876 10004 33928 10013
rect 33968 10047 34020 10056
rect 33968 10013 33977 10047
rect 33977 10013 34011 10047
rect 34011 10013 34020 10047
rect 33968 10004 34020 10013
rect 34060 10004 34112 10056
rect 22836 9911 22888 9920
rect 22836 9877 22845 9911
rect 22845 9877 22879 9911
rect 22879 9877 22888 9911
rect 22836 9868 22888 9877
rect 23480 9868 23532 9920
rect 24768 9911 24820 9920
rect 24768 9877 24777 9911
rect 24777 9877 24811 9911
rect 24811 9877 24820 9911
rect 24768 9868 24820 9877
rect 26516 9868 26568 9920
rect 28908 9911 28960 9920
rect 28908 9877 28917 9911
rect 28917 9877 28951 9911
rect 28951 9877 28960 9911
rect 28908 9868 28960 9877
rect 29092 9911 29144 9920
rect 29092 9877 29101 9911
rect 29101 9877 29135 9911
rect 29135 9877 29144 9911
rect 29092 9868 29144 9877
rect 34336 9936 34388 9988
rect 30380 9868 30432 9920
rect 30840 9868 30892 9920
rect 30932 9911 30984 9920
rect 30932 9877 30941 9911
rect 30941 9877 30975 9911
rect 30975 9877 30984 9911
rect 30932 9868 30984 9877
rect 32128 9868 32180 9920
rect 33232 9868 33284 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4344 9664 4396 9716
rect 3056 9596 3108 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 3792 9528 3844 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 4620 9528 4672 9580
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5448 9528 5500 9580
rect 6552 9664 6604 9716
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 7840 9664 7892 9716
rect 8208 9596 8260 9648
rect 8300 9528 8352 9580
rect 8576 9596 8628 9648
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 10232 9664 10284 9716
rect 12072 9664 12124 9716
rect 12440 9664 12492 9716
rect 14280 9664 14332 9716
rect 14740 9664 14792 9716
rect 20076 9664 20128 9716
rect 10876 9596 10928 9648
rect 8852 9571 8904 9580
rect 8852 9537 8867 9571
rect 8867 9537 8901 9571
rect 8901 9537 8904 9571
rect 8852 9528 8904 9537
rect 10232 9528 10284 9580
rect 10600 9528 10652 9580
rect 5356 9392 5408 9444
rect 7288 9460 7340 9512
rect 7840 9460 7892 9512
rect 7932 9460 7984 9512
rect 10140 9460 10192 9512
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 12624 9528 12676 9580
rect 19432 9596 19484 9648
rect 20812 9664 20864 9716
rect 22284 9664 22336 9716
rect 22376 9664 22428 9716
rect 22744 9664 22796 9716
rect 24492 9664 24544 9716
rect 13084 9528 13136 9580
rect 14740 9528 14792 9580
rect 15200 9528 15252 9580
rect 18512 9528 18564 9580
rect 20720 9528 20772 9580
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 4068 9324 4120 9376
rect 4436 9324 4488 9376
rect 4804 9324 4856 9376
rect 4896 9324 4948 9376
rect 5172 9324 5224 9376
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 12532 9392 12584 9444
rect 13820 9460 13872 9512
rect 15016 9460 15068 9512
rect 17960 9460 18012 9512
rect 19984 9460 20036 9512
rect 20536 9460 20588 9512
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 21088 9639 21140 9648
rect 21088 9605 21097 9639
rect 21097 9605 21131 9639
rect 21131 9605 21140 9639
rect 21088 9596 21140 9605
rect 22836 9528 22888 9580
rect 28540 9664 28592 9716
rect 24676 9571 24728 9580
rect 24676 9537 24685 9571
rect 24685 9537 24719 9571
rect 24719 9537 24728 9571
rect 24676 9528 24728 9537
rect 21272 9460 21324 9512
rect 21456 9460 21508 9512
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 14832 9392 14884 9444
rect 19800 9435 19852 9444
rect 19800 9401 19809 9435
rect 19809 9401 19843 9435
rect 19843 9401 19852 9435
rect 19800 9392 19852 9401
rect 17224 9324 17276 9376
rect 18052 9324 18104 9376
rect 21180 9324 21232 9376
rect 23848 9392 23900 9444
rect 24952 9528 25004 9580
rect 25044 9528 25096 9580
rect 25596 9571 25648 9580
rect 25596 9537 25605 9571
rect 25605 9537 25639 9571
rect 25639 9537 25648 9571
rect 25596 9528 25648 9537
rect 25872 9571 25924 9580
rect 25872 9537 25881 9571
rect 25881 9537 25915 9571
rect 25915 9537 25924 9571
rect 25872 9528 25924 9537
rect 25964 9528 26016 9580
rect 27252 9596 27304 9648
rect 27344 9528 27396 9580
rect 27620 9571 27672 9580
rect 27620 9537 27629 9571
rect 27629 9537 27663 9571
rect 27663 9537 27672 9571
rect 27620 9528 27672 9537
rect 29000 9528 29052 9580
rect 29368 9528 29420 9580
rect 27712 9460 27764 9512
rect 28540 9460 28592 9512
rect 30196 9596 30248 9648
rect 30564 9664 30616 9716
rect 32220 9596 32272 9648
rect 33968 9664 34020 9716
rect 32864 9639 32916 9648
rect 32864 9605 32873 9639
rect 32873 9605 32907 9639
rect 32907 9605 32916 9639
rect 32864 9596 32916 9605
rect 33140 9596 33192 9648
rect 30840 9571 30892 9580
rect 30840 9537 30849 9571
rect 30849 9537 30883 9571
rect 30883 9537 30892 9571
rect 30840 9528 30892 9537
rect 30932 9528 30984 9580
rect 32588 9528 32640 9580
rect 25044 9392 25096 9444
rect 29552 9392 29604 9444
rect 21548 9324 21600 9376
rect 21916 9324 21968 9376
rect 22744 9367 22796 9376
rect 22744 9333 22753 9367
rect 22753 9333 22787 9367
rect 22787 9333 22796 9367
rect 22744 9324 22796 9333
rect 22836 9324 22888 9376
rect 23572 9324 23624 9376
rect 23940 9324 23992 9376
rect 24952 9324 25004 9376
rect 26240 9324 26292 9376
rect 26332 9324 26384 9376
rect 26792 9324 26844 9376
rect 28816 9324 28868 9376
rect 29276 9367 29328 9376
rect 29276 9333 29285 9367
rect 29285 9333 29319 9367
rect 29319 9333 29328 9367
rect 29276 9324 29328 9333
rect 30656 9503 30708 9512
rect 30656 9469 30665 9503
rect 30665 9469 30699 9503
rect 30699 9469 30708 9503
rect 30656 9460 30708 9469
rect 31208 9435 31260 9444
rect 31208 9401 31217 9435
rect 31217 9401 31251 9435
rect 31251 9401 31260 9435
rect 31208 9392 31260 9401
rect 31392 9392 31444 9444
rect 31944 9392 31996 9444
rect 33232 9392 33284 9444
rect 34336 9392 34388 9444
rect 32036 9324 32088 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1676 9120 1728 9172
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 3884 8984 3936 9036
rect 4252 8984 4304 9036
rect 4068 8916 4120 8968
rect 4896 9120 4948 9172
rect 4988 9120 5040 9172
rect 5356 9120 5408 9172
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 12072 9120 12124 9172
rect 12440 9120 12492 9172
rect 15016 9120 15068 9172
rect 17684 9163 17736 9172
rect 17684 9129 17693 9163
rect 17693 9129 17727 9163
rect 17727 9129 17736 9163
rect 17684 9120 17736 9129
rect 18512 9120 18564 9172
rect 22468 9120 22520 9172
rect 22744 9163 22796 9172
rect 22744 9129 22753 9163
rect 22753 9129 22787 9163
rect 22787 9129 22796 9163
rect 22744 9120 22796 9129
rect 22836 9120 22888 9172
rect 5080 8984 5132 9036
rect 4712 8916 4764 8968
rect 5448 9052 5500 9104
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 8576 8916 8628 8968
rect 10324 8984 10376 9036
rect 4896 8848 4948 8900
rect 8208 8848 8260 8900
rect 8484 8848 8536 8900
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 11152 8984 11204 9036
rect 13636 9052 13688 9104
rect 12808 8984 12860 9036
rect 13268 8984 13320 9036
rect 17224 9052 17276 9104
rect 11980 8959 12032 8968
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 14280 8916 14332 8968
rect 14464 8916 14516 8968
rect 13544 8848 13596 8900
rect 15016 8848 15068 8900
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 17868 8984 17920 9036
rect 20628 8984 20680 9036
rect 20904 8984 20956 9036
rect 23388 9120 23440 9172
rect 23664 9120 23716 9172
rect 26332 9120 26384 9172
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 18052 8916 18104 8968
rect 19524 8916 19576 8968
rect 20536 8959 20588 8968
rect 20536 8925 20545 8959
rect 20545 8925 20579 8959
rect 20579 8925 20588 8959
rect 20536 8916 20588 8925
rect 20812 8916 20864 8968
rect 16488 8848 16540 8900
rect 18328 8848 18380 8900
rect 23112 8984 23164 9036
rect 22560 8916 22612 8968
rect 22836 8916 22888 8968
rect 24308 9052 24360 9104
rect 23296 9027 23348 9036
rect 23296 8993 23305 9027
rect 23305 8993 23339 9027
rect 23339 8993 23348 9027
rect 23296 8984 23348 8993
rect 23940 8916 23992 8968
rect 24124 8959 24176 8968
rect 24124 8925 24133 8959
rect 24133 8925 24167 8959
rect 24167 8925 24176 8959
rect 24124 8916 24176 8925
rect 940 8780 992 8832
rect 3516 8823 3568 8832
rect 3516 8789 3525 8823
rect 3525 8789 3559 8823
rect 3559 8789 3568 8823
rect 3516 8780 3568 8789
rect 8300 8780 8352 8832
rect 8760 8780 8812 8832
rect 9496 8780 9548 8832
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 12440 8780 12492 8832
rect 12624 8780 12676 8832
rect 14648 8780 14700 8832
rect 15200 8780 15252 8832
rect 20168 8780 20220 8832
rect 20628 8780 20680 8832
rect 23848 8848 23900 8900
rect 24400 8959 24452 8968
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 24768 8984 24820 9036
rect 26424 9052 26476 9104
rect 25780 9027 25832 9036
rect 25780 8993 25789 9027
rect 25789 8993 25823 9027
rect 25823 8993 25832 9027
rect 25780 8984 25832 8993
rect 27160 9120 27212 9172
rect 28724 9120 28776 9172
rect 29276 9120 29328 9172
rect 30840 9120 30892 9172
rect 32588 9163 32640 9172
rect 32588 9129 32597 9163
rect 32597 9129 32631 9163
rect 32631 9129 32640 9163
rect 32588 9120 32640 9129
rect 33140 9120 33192 9172
rect 33600 9120 33652 9172
rect 25596 8959 25648 8968
rect 25596 8925 25605 8959
rect 25605 8925 25639 8959
rect 25639 8925 25648 8959
rect 25596 8916 25648 8925
rect 25688 8916 25740 8968
rect 26240 8959 26292 8968
rect 26240 8925 26249 8959
rect 26249 8925 26283 8959
rect 26283 8925 26292 8959
rect 26240 8916 26292 8925
rect 26332 8959 26384 8968
rect 26332 8925 26341 8959
rect 26341 8925 26375 8959
rect 26375 8925 26384 8959
rect 26332 8916 26384 8925
rect 24676 8891 24728 8900
rect 21364 8823 21416 8832
rect 21364 8789 21373 8823
rect 21373 8789 21407 8823
rect 21407 8789 21416 8823
rect 21364 8780 21416 8789
rect 23020 8780 23072 8832
rect 24676 8857 24685 8891
rect 24685 8857 24719 8891
rect 24719 8857 24728 8891
rect 24676 8848 24728 8857
rect 24492 8780 24544 8832
rect 25136 8780 25188 8832
rect 26792 8916 26844 8968
rect 26884 8959 26936 8968
rect 26884 8925 26893 8959
rect 26893 8925 26927 8959
rect 26927 8925 26936 8959
rect 26884 8916 26936 8925
rect 26976 8916 27028 8968
rect 27804 8984 27856 9036
rect 28448 8959 28500 8968
rect 28448 8925 28471 8959
rect 28471 8925 28500 8959
rect 28448 8916 28500 8925
rect 28816 8959 28868 8968
rect 28816 8925 28825 8959
rect 28825 8925 28859 8959
rect 28859 8925 28868 8959
rect 28816 8916 28868 8925
rect 28724 8848 28776 8900
rect 29092 8984 29144 9036
rect 31392 8984 31444 9036
rect 32036 9052 32088 9104
rect 29552 8959 29604 8968
rect 29552 8925 29561 8959
rect 29561 8925 29595 8959
rect 29595 8925 29604 8959
rect 29552 8916 29604 8925
rect 30104 8916 30156 8968
rect 30380 8916 30432 8968
rect 31392 8848 31444 8900
rect 31852 8916 31904 8968
rect 31944 8959 31996 8968
rect 31944 8925 31953 8959
rect 31953 8925 31987 8959
rect 31987 8925 31996 8959
rect 31944 8916 31996 8925
rect 32956 8984 33008 9036
rect 32496 8916 32548 8968
rect 32220 8848 32272 8900
rect 33140 8959 33192 8968
rect 33140 8925 33149 8959
rect 33149 8925 33183 8959
rect 33183 8925 33192 8959
rect 33140 8916 33192 8925
rect 36636 8984 36688 9036
rect 33784 8916 33836 8968
rect 38108 8916 38160 8968
rect 25688 8780 25740 8832
rect 25964 8823 26016 8832
rect 25964 8789 25973 8823
rect 25973 8789 26007 8823
rect 26007 8789 26016 8823
rect 25964 8780 26016 8789
rect 26240 8780 26292 8832
rect 26976 8780 27028 8832
rect 27252 8780 27304 8832
rect 29184 8780 29236 8832
rect 29920 8823 29972 8832
rect 29920 8789 29929 8823
rect 29929 8789 29963 8823
rect 29963 8789 29972 8823
rect 29920 8780 29972 8789
rect 30840 8780 30892 8832
rect 33140 8780 33192 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2872 8576 2924 8628
rect 3516 8576 3568 8628
rect 4068 8576 4120 8628
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 8760 8576 8812 8628
rect 10048 8576 10100 8628
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 4068 8440 4120 8492
rect 4712 8440 4764 8492
rect 5172 8440 5224 8492
rect 2596 8347 2648 8356
rect 2596 8313 2605 8347
rect 2605 8313 2639 8347
rect 2639 8313 2648 8347
rect 2596 8304 2648 8313
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 7932 8372 7984 8424
rect 8300 8508 8352 8560
rect 13820 8576 13872 8628
rect 14556 8576 14608 8628
rect 8484 8440 8536 8492
rect 4988 8236 5040 8288
rect 7472 8304 7524 8356
rect 11888 8440 11940 8492
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 14648 8508 14700 8560
rect 11980 8372 12032 8424
rect 15200 8372 15252 8424
rect 16672 8576 16724 8628
rect 18328 8508 18380 8560
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 19340 8440 19392 8492
rect 19984 8576 20036 8628
rect 20076 8576 20128 8628
rect 20812 8619 20864 8628
rect 20812 8585 20821 8619
rect 20821 8585 20855 8619
rect 20855 8585 20864 8619
rect 20812 8576 20864 8585
rect 19156 8372 19208 8424
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 20168 8483 20220 8492
rect 20168 8449 20177 8483
rect 20177 8449 20211 8483
rect 20211 8449 20220 8483
rect 20168 8440 20220 8449
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 20904 8483 20956 8492
rect 20904 8449 20913 8483
rect 20913 8449 20947 8483
rect 20947 8449 20956 8483
rect 20904 8440 20956 8449
rect 22836 8576 22888 8628
rect 23204 8576 23256 8628
rect 23572 8576 23624 8628
rect 23848 8576 23900 8628
rect 24124 8576 24176 8628
rect 26240 8576 26292 8628
rect 26884 8576 26936 8628
rect 28172 8576 28224 8628
rect 29552 8576 29604 8628
rect 29920 8576 29972 8628
rect 30656 8576 30708 8628
rect 31760 8576 31812 8628
rect 32956 8576 33008 8628
rect 23296 8551 23348 8560
rect 19984 8415 20036 8424
rect 19984 8381 19993 8415
rect 19993 8381 20027 8415
rect 20027 8381 20036 8415
rect 23296 8517 23305 8551
rect 23305 8517 23339 8551
rect 23339 8517 23348 8551
rect 23296 8508 23348 8517
rect 24952 8508 25004 8560
rect 22652 8440 22704 8492
rect 23112 8483 23164 8492
rect 23112 8449 23119 8483
rect 23119 8449 23164 8483
rect 19984 8372 20036 8381
rect 22744 8415 22796 8424
rect 22744 8381 22753 8415
rect 22753 8381 22787 8415
rect 22787 8381 22796 8415
rect 22744 8372 22796 8381
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 12348 8236 12400 8288
rect 13268 8236 13320 8288
rect 14740 8236 14792 8288
rect 19892 8304 19944 8356
rect 23112 8440 23164 8449
rect 23756 8440 23808 8492
rect 25780 8440 25832 8492
rect 27712 8508 27764 8560
rect 29368 8508 29420 8560
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 23020 8304 23072 8356
rect 23204 8304 23256 8356
rect 24952 8304 25004 8356
rect 20812 8236 20864 8288
rect 23572 8279 23624 8288
rect 23572 8245 23581 8279
rect 23581 8245 23615 8279
rect 23615 8245 23624 8279
rect 23572 8236 23624 8245
rect 23940 8236 23992 8288
rect 25596 8372 25648 8424
rect 26884 8372 26936 8424
rect 28724 8440 28776 8492
rect 28816 8483 28868 8492
rect 28816 8449 28825 8483
rect 28825 8449 28859 8483
rect 28859 8449 28868 8483
rect 28816 8440 28868 8449
rect 30012 8440 30064 8492
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 27620 8304 27672 8356
rect 30564 8372 30616 8424
rect 31760 8415 31812 8424
rect 31760 8381 31769 8415
rect 31769 8381 31803 8415
rect 31803 8381 31812 8415
rect 31760 8372 31812 8381
rect 33784 8440 33836 8492
rect 26516 8236 26568 8288
rect 28264 8236 28316 8288
rect 28356 8279 28408 8288
rect 28356 8245 28365 8279
rect 28365 8245 28399 8279
rect 28399 8245 28408 8279
rect 28356 8236 28408 8245
rect 29368 8304 29420 8356
rect 28632 8236 28684 8288
rect 30840 8304 30892 8356
rect 33324 8372 33376 8424
rect 29552 8236 29604 8288
rect 33232 8304 33284 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 4988 8032 5040 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 6092 7896 6144 7948
rect 7840 7964 7892 8016
rect 9404 8032 9456 8084
rect 12164 8032 12216 8084
rect 12808 8032 12860 8084
rect 14280 8075 14332 8084
rect 14280 8041 14289 8075
rect 14289 8041 14323 8075
rect 14323 8041 14332 8075
rect 14280 8032 14332 8041
rect 25688 8032 25740 8084
rect 26884 8032 26936 8084
rect 27160 8032 27212 8084
rect 27344 8032 27396 8084
rect 4712 7760 4764 7812
rect 6000 7803 6052 7812
rect 6000 7769 6009 7803
rect 6009 7769 6043 7803
rect 6043 7769 6052 7803
rect 6000 7760 6052 7769
rect 7472 7760 7524 7812
rect 9220 7803 9272 7812
rect 9220 7769 9229 7803
rect 9229 7769 9263 7803
rect 9263 7769 9272 7803
rect 9220 7760 9272 7769
rect 11060 7828 11112 7880
rect 11520 7896 11572 7948
rect 12992 7896 13044 7948
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 14372 7964 14424 8016
rect 19432 7964 19484 8016
rect 28724 8032 28776 8084
rect 30012 8032 30064 8084
rect 31852 8032 31904 8084
rect 30564 7964 30616 8016
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 14832 7939 14884 7948
rect 14832 7905 14841 7939
rect 14841 7905 14875 7939
rect 14875 7905 14884 7939
rect 14832 7896 14884 7905
rect 14464 7828 14516 7880
rect 17592 7828 17644 7880
rect 18144 7828 18196 7880
rect 20536 7896 20588 7948
rect 22468 7896 22520 7948
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 20076 7828 20128 7880
rect 20168 7828 20220 7880
rect 28356 7896 28408 7948
rect 28448 7896 28500 7948
rect 20536 7760 20588 7812
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 23480 7828 23532 7837
rect 23572 7828 23624 7880
rect 24032 7828 24084 7880
rect 25964 7828 26016 7880
rect 26976 7871 27028 7880
rect 26976 7837 26985 7871
rect 26985 7837 27019 7871
rect 27019 7837 27028 7871
rect 26976 7828 27028 7837
rect 27160 7871 27212 7880
rect 27160 7837 27169 7871
rect 27169 7837 27203 7871
rect 27203 7837 27212 7871
rect 27160 7828 27212 7837
rect 28172 7828 28224 7880
rect 28816 7871 28868 7880
rect 28816 7837 28825 7871
rect 28825 7837 28859 7871
rect 28859 7837 28868 7871
rect 28816 7828 28868 7837
rect 9496 7692 9548 7744
rect 12164 7735 12216 7744
rect 12164 7701 12173 7735
rect 12173 7701 12207 7735
rect 12207 7701 12216 7735
rect 12164 7692 12216 7701
rect 12256 7692 12308 7744
rect 13268 7692 13320 7744
rect 20352 7692 20404 7744
rect 20628 7692 20680 7744
rect 23020 7735 23072 7744
rect 23020 7701 23029 7735
rect 23029 7701 23063 7735
rect 23063 7701 23072 7735
rect 23020 7692 23072 7701
rect 27344 7692 27396 7744
rect 27436 7692 27488 7744
rect 27528 7735 27580 7744
rect 27528 7701 27537 7735
rect 27537 7701 27571 7735
rect 27571 7701 27580 7735
rect 27528 7692 27580 7701
rect 28540 7760 28592 7812
rect 29552 7871 29604 7880
rect 29552 7837 29561 7871
rect 29561 7837 29595 7871
rect 29595 7837 29604 7871
rect 29552 7828 29604 7837
rect 30288 7828 30340 7880
rect 30564 7871 30616 7880
rect 30564 7837 30573 7871
rect 30573 7837 30607 7871
rect 30607 7837 30616 7871
rect 30564 7828 30616 7837
rect 30656 7828 30708 7880
rect 30840 7828 30892 7880
rect 31300 7828 31352 7880
rect 31668 7964 31720 8016
rect 31760 7896 31812 7948
rect 31668 7760 31720 7812
rect 31300 7735 31352 7744
rect 31300 7701 31309 7735
rect 31309 7701 31343 7735
rect 31343 7701 31352 7735
rect 31300 7692 31352 7701
rect 31484 7692 31536 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4988 7488 5040 7540
rect 6000 7488 6052 7540
rect 6644 7488 6696 7540
rect 9220 7488 9272 7540
rect 13268 7488 13320 7540
rect 15292 7531 15344 7540
rect 15292 7497 15301 7531
rect 15301 7497 15335 7531
rect 15335 7497 15344 7531
rect 15292 7488 15344 7497
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 4712 7352 4764 7404
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 10140 7420 10192 7472
rect 14280 7420 14332 7472
rect 15108 7420 15160 7472
rect 19432 7488 19484 7540
rect 19892 7488 19944 7540
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 10968 7352 11020 7404
rect 11612 7395 11664 7404
rect 11612 7361 11621 7395
rect 11621 7361 11655 7395
rect 11655 7361 11664 7395
rect 11612 7352 11664 7361
rect 17040 7352 17092 7404
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 20536 7531 20588 7540
rect 20536 7497 20545 7531
rect 20545 7497 20579 7531
rect 20579 7497 20588 7531
rect 20536 7488 20588 7497
rect 22376 7488 22428 7540
rect 22744 7488 22796 7540
rect 23020 7488 23072 7540
rect 23480 7488 23532 7540
rect 4620 7327 4672 7336
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 5080 7284 5132 7336
rect 5172 7284 5224 7336
rect 9496 7284 9548 7336
rect 11704 7284 11756 7336
rect 12348 7284 12400 7336
rect 12992 7284 13044 7336
rect 14832 7284 14884 7336
rect 19892 7352 19944 7404
rect 20168 7395 20220 7404
rect 20168 7361 20177 7395
rect 20177 7361 20211 7395
rect 20211 7361 20220 7395
rect 20168 7352 20220 7361
rect 20260 7395 20312 7404
rect 20260 7361 20269 7395
rect 20269 7361 20303 7395
rect 20303 7361 20312 7395
rect 20260 7352 20312 7361
rect 21640 7420 21692 7472
rect 9312 7216 9364 7268
rect 11060 7216 11112 7268
rect 14280 7216 14332 7268
rect 20352 7216 20404 7268
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 22928 7463 22980 7472
rect 22928 7429 22937 7463
rect 22937 7429 22971 7463
rect 22971 7429 22980 7463
rect 22928 7420 22980 7429
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 27344 7488 27396 7540
rect 24952 7420 25004 7472
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 24768 7395 24820 7404
rect 24768 7361 24777 7395
rect 24777 7361 24811 7395
rect 24811 7361 24820 7395
rect 24768 7352 24820 7361
rect 26516 7420 26568 7472
rect 26700 7420 26752 7472
rect 26884 7420 26936 7472
rect 21364 7284 21416 7336
rect 21732 7284 21784 7336
rect 23112 7284 23164 7336
rect 25596 7284 25648 7336
rect 21180 7259 21232 7268
rect 21180 7225 21189 7259
rect 21189 7225 21223 7259
rect 21223 7225 21232 7259
rect 21180 7216 21232 7225
rect 23664 7216 23716 7268
rect 27252 7395 27304 7404
rect 27252 7361 27261 7395
rect 27261 7361 27295 7395
rect 27295 7361 27304 7395
rect 27252 7352 27304 7361
rect 27344 7395 27396 7404
rect 27344 7361 27353 7395
rect 27353 7361 27387 7395
rect 27387 7361 27396 7395
rect 27344 7352 27396 7361
rect 31300 7488 31352 7540
rect 31484 7488 31536 7540
rect 28172 7420 28224 7472
rect 3700 7148 3752 7200
rect 11428 7148 11480 7200
rect 12256 7148 12308 7200
rect 15200 7148 15252 7200
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 19340 7148 19392 7200
rect 20168 7148 20220 7200
rect 20720 7148 20772 7200
rect 24952 7191 25004 7200
rect 24952 7157 24961 7191
rect 24961 7157 24995 7191
rect 24995 7157 25004 7191
rect 24952 7148 25004 7157
rect 25136 7191 25188 7200
rect 25136 7157 25145 7191
rect 25145 7157 25179 7191
rect 25179 7157 25188 7191
rect 25136 7148 25188 7157
rect 25688 7191 25740 7200
rect 25688 7157 25697 7191
rect 25697 7157 25731 7191
rect 25731 7157 25740 7191
rect 25688 7148 25740 7157
rect 26424 7216 26476 7268
rect 28448 7395 28500 7404
rect 28448 7361 28457 7395
rect 28457 7361 28491 7395
rect 28491 7361 28500 7395
rect 28448 7352 28500 7361
rect 31024 7420 31076 7472
rect 29276 7395 29328 7404
rect 29276 7361 29285 7395
rect 29285 7361 29319 7395
rect 29319 7361 29328 7395
rect 29276 7352 29328 7361
rect 29368 7352 29420 7404
rect 29092 7327 29144 7336
rect 29092 7293 29101 7327
rect 29101 7293 29135 7327
rect 29135 7293 29144 7327
rect 29092 7284 29144 7293
rect 30288 7352 30340 7404
rect 31300 7327 31352 7336
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 31852 7352 31904 7404
rect 33692 7531 33744 7540
rect 33692 7497 33701 7531
rect 33701 7497 33735 7531
rect 33735 7497 33744 7531
rect 33692 7488 33744 7497
rect 32128 7284 32180 7336
rect 27160 7148 27212 7200
rect 29368 7148 29420 7200
rect 31760 7148 31812 7200
rect 33324 7216 33376 7268
rect 34060 7148 34112 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 5264 6944 5316 6996
rect 5080 6876 5132 6928
rect 11060 6944 11112 6996
rect 11520 6987 11572 6996
rect 11520 6953 11529 6987
rect 11529 6953 11563 6987
rect 11563 6953 11572 6987
rect 11520 6944 11572 6953
rect 17224 6944 17276 6996
rect 17408 6944 17460 6996
rect 18604 6944 18656 6996
rect 19892 6944 19944 6996
rect 20076 6987 20128 6996
rect 20076 6953 20085 6987
rect 20085 6953 20119 6987
rect 20119 6953 20128 6987
rect 20076 6944 20128 6953
rect 20168 6944 20220 6996
rect 21640 6944 21692 6996
rect 22468 6944 22520 6996
rect 23940 6944 23992 6996
rect 25596 6987 25648 6996
rect 25596 6953 25605 6987
rect 25605 6953 25639 6987
rect 25639 6953 25648 6987
rect 25596 6944 25648 6953
rect 27528 6944 27580 6996
rect 28264 6944 28316 6996
rect 29920 6944 29972 6996
rect 31300 6944 31352 6996
rect 33140 6987 33192 6996
rect 33140 6953 33149 6987
rect 33149 6953 33183 6987
rect 33183 6953 33192 6987
rect 33140 6944 33192 6953
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 7196 6808 7248 6860
rect 8116 6808 8168 6860
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 3700 6740 3752 6792
rect 7472 6740 7524 6792
rect 4712 6604 4764 6656
rect 6460 6715 6512 6724
rect 6460 6681 6469 6715
rect 6469 6681 6503 6715
rect 6503 6681 6512 6715
rect 6460 6672 6512 6681
rect 7932 6740 7984 6792
rect 8208 6740 8260 6792
rect 8300 6672 8352 6724
rect 17040 6919 17092 6928
rect 17040 6885 17049 6919
rect 17049 6885 17083 6919
rect 17083 6885 17092 6919
rect 17040 6876 17092 6885
rect 17592 6876 17644 6928
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 11612 6808 11664 6817
rect 18420 6808 18472 6860
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 10416 6604 10468 6656
rect 11244 6604 11296 6656
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 16580 6672 16632 6724
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 18052 6783 18104 6792
rect 18052 6749 18061 6783
rect 18061 6749 18095 6783
rect 18095 6749 18104 6783
rect 18052 6740 18104 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 19340 6808 19392 6860
rect 18788 6740 18840 6792
rect 20260 6876 20312 6928
rect 21732 6919 21784 6928
rect 21732 6885 21741 6919
rect 21741 6885 21775 6919
rect 21775 6885 21784 6919
rect 21732 6876 21784 6885
rect 22284 6876 22336 6928
rect 21180 6740 21232 6792
rect 21640 6740 21692 6792
rect 22100 6808 22152 6860
rect 21916 6740 21968 6792
rect 23112 6808 23164 6860
rect 23204 6715 23256 6724
rect 23204 6681 23213 6715
rect 23213 6681 23247 6715
rect 23247 6681 23256 6715
rect 23204 6672 23256 6681
rect 23848 6876 23900 6928
rect 27252 6876 27304 6928
rect 24952 6808 25004 6860
rect 25136 6783 25188 6792
rect 25136 6749 25145 6783
rect 25145 6749 25179 6783
rect 25179 6749 25188 6783
rect 25136 6740 25188 6749
rect 25504 6740 25556 6792
rect 27068 6740 27120 6792
rect 27804 6876 27856 6928
rect 27988 6876 28040 6928
rect 27896 6783 27948 6792
rect 27896 6749 27903 6783
rect 27903 6749 27948 6783
rect 27896 6740 27948 6749
rect 29276 6808 29328 6860
rect 30472 6851 30524 6860
rect 30472 6817 30481 6851
rect 30481 6817 30515 6851
rect 30515 6817 30524 6851
rect 30472 6808 30524 6817
rect 28172 6783 28224 6792
rect 28172 6749 28186 6783
rect 28186 6749 28220 6783
rect 28220 6749 28224 6783
rect 28172 6740 28224 6749
rect 28356 6740 28408 6792
rect 28448 6740 28500 6792
rect 18052 6604 18104 6656
rect 18696 6604 18748 6656
rect 21364 6647 21416 6656
rect 21364 6613 21373 6647
rect 21373 6613 21407 6647
rect 21407 6613 21416 6647
rect 21364 6604 21416 6613
rect 22560 6604 22612 6656
rect 22836 6604 22888 6656
rect 25596 6604 25648 6656
rect 28632 6604 28684 6656
rect 29184 6740 29236 6792
rect 30564 6740 30616 6792
rect 30656 6783 30708 6792
rect 30656 6749 30665 6783
rect 30665 6749 30699 6783
rect 30699 6749 30708 6783
rect 30656 6740 30708 6749
rect 31208 6808 31260 6860
rect 32496 6851 32548 6860
rect 32496 6817 32505 6851
rect 32505 6817 32539 6851
rect 32539 6817 32548 6851
rect 32496 6808 32548 6817
rect 31944 6740 31996 6792
rect 32588 6672 32640 6724
rect 31116 6604 31168 6656
rect 31208 6604 31260 6656
rect 33232 6740 33284 6792
rect 33140 6604 33192 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 6460 6400 6512 6452
rect 8024 6400 8076 6452
rect 8208 6400 8260 6452
rect 8300 6400 8352 6452
rect 8392 6400 8444 6452
rect 9036 6400 9088 6452
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 18052 6400 18104 6452
rect 18420 6400 18472 6452
rect 18512 6400 18564 6452
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 12072 6332 12124 6384
rect 12164 6332 12216 6384
rect 12808 6332 12860 6384
rect 8392 6196 8444 6248
rect 9220 6196 9272 6248
rect 8116 6128 8168 6180
rect 8300 6171 8352 6180
rect 8300 6137 8309 6171
rect 8309 6137 8343 6171
rect 8343 6137 8352 6171
rect 8300 6128 8352 6137
rect 8576 6128 8628 6180
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 13728 6264 13780 6316
rect 19340 6400 19392 6452
rect 19432 6400 19484 6452
rect 22376 6400 22428 6452
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 13636 6239 13688 6248
rect 13636 6205 13645 6239
rect 13645 6205 13679 6239
rect 13679 6205 13688 6239
rect 13636 6196 13688 6205
rect 19156 6264 19208 6316
rect 18604 6196 18656 6248
rect 21916 6264 21968 6316
rect 22928 6400 22980 6452
rect 23204 6400 23256 6452
rect 24124 6400 24176 6452
rect 25136 6400 25188 6452
rect 22744 6307 22796 6316
rect 22744 6273 22753 6307
rect 22753 6273 22787 6307
rect 22787 6273 22796 6307
rect 22744 6264 22796 6273
rect 23112 6264 23164 6316
rect 24400 6264 24452 6316
rect 15200 6128 15252 6180
rect 15752 6128 15804 6180
rect 9404 6060 9456 6112
rect 13544 6060 13596 6112
rect 14004 6060 14056 6112
rect 15108 6060 15160 6112
rect 18328 6103 18380 6112
rect 18328 6069 18337 6103
rect 18337 6069 18371 6103
rect 18371 6069 18380 6103
rect 18328 6060 18380 6069
rect 23848 6196 23900 6248
rect 25596 6332 25648 6384
rect 26516 6332 26568 6384
rect 24584 6307 24636 6316
rect 24584 6273 24593 6307
rect 24593 6273 24627 6307
rect 24627 6273 24636 6307
rect 24584 6264 24636 6273
rect 24952 6264 25004 6316
rect 26792 6332 26844 6384
rect 28448 6400 28500 6452
rect 27896 6196 27948 6248
rect 28908 6332 28960 6384
rect 31208 6400 31260 6452
rect 31944 6443 31996 6452
rect 31944 6409 31953 6443
rect 31953 6409 31987 6443
rect 31987 6409 31996 6443
rect 31944 6400 31996 6409
rect 32128 6443 32180 6452
rect 32128 6409 32137 6443
rect 32137 6409 32171 6443
rect 32171 6409 32180 6443
rect 32128 6400 32180 6409
rect 31760 6375 31812 6384
rect 31760 6341 31769 6375
rect 31769 6341 31803 6375
rect 31803 6341 31812 6375
rect 31760 6332 31812 6341
rect 32036 6332 32088 6384
rect 28448 6264 28500 6316
rect 30104 6307 30156 6316
rect 30104 6273 30113 6307
rect 30113 6273 30147 6307
rect 30147 6273 30156 6307
rect 30104 6264 30156 6273
rect 30380 6264 30432 6316
rect 33140 6332 33192 6384
rect 32496 6307 32548 6316
rect 32496 6273 32505 6307
rect 32505 6273 32539 6307
rect 32539 6273 32548 6307
rect 32496 6264 32548 6273
rect 32588 6307 32640 6316
rect 32588 6273 32597 6307
rect 32597 6273 32631 6307
rect 32631 6273 32640 6307
rect 32588 6264 32640 6273
rect 27620 6128 27672 6180
rect 29644 6196 29696 6248
rect 28724 6128 28776 6180
rect 32036 6196 32088 6248
rect 19340 6060 19392 6112
rect 22560 6060 22612 6112
rect 22836 6060 22888 6112
rect 26516 6060 26568 6112
rect 33324 6060 33376 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 7932 5856 7984 5908
rect 8576 5856 8628 5908
rect 9404 5856 9456 5908
rect 9220 5788 9272 5840
rect 8208 5652 8260 5704
rect 8392 5652 8444 5704
rect 9036 5695 9088 5704
rect 9036 5661 9046 5695
rect 9046 5661 9080 5695
rect 9080 5661 9088 5695
rect 9036 5652 9088 5661
rect 9404 5695 9456 5704
rect 9404 5661 9418 5695
rect 9418 5661 9452 5695
rect 9452 5661 9456 5695
rect 11612 5856 11664 5908
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 13176 5856 13228 5908
rect 12716 5788 12768 5840
rect 9404 5652 9456 5661
rect 9772 5652 9824 5704
rect 12164 5652 12216 5704
rect 13544 5763 13596 5772
rect 13544 5729 13553 5763
rect 13553 5729 13587 5763
rect 13587 5729 13596 5763
rect 13544 5720 13596 5729
rect 14004 5652 14056 5704
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 10048 5516 10100 5568
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 12256 5516 12308 5568
rect 12808 5516 12860 5568
rect 15568 5856 15620 5908
rect 19984 5856 20036 5908
rect 22744 5856 22796 5908
rect 24584 5856 24636 5908
rect 28172 5856 28224 5908
rect 28356 5899 28408 5908
rect 28356 5865 28365 5899
rect 28365 5865 28399 5899
rect 28399 5865 28408 5899
rect 28356 5856 28408 5865
rect 29368 5856 29420 5908
rect 30104 5899 30156 5908
rect 30104 5865 30113 5899
rect 30113 5865 30147 5899
rect 30147 5865 30156 5899
rect 30104 5856 30156 5865
rect 31116 5899 31168 5908
rect 31116 5865 31125 5899
rect 31125 5865 31159 5899
rect 31159 5865 31168 5899
rect 31116 5856 31168 5865
rect 32036 5899 32088 5908
rect 32036 5865 32045 5899
rect 32045 5865 32079 5899
rect 32079 5865 32088 5899
rect 32036 5856 32088 5865
rect 32496 5856 32548 5908
rect 15108 5720 15160 5772
rect 22928 5720 22980 5772
rect 14464 5584 14516 5636
rect 15476 5584 15528 5636
rect 20076 5652 20128 5704
rect 22560 5695 22612 5704
rect 22560 5661 22569 5695
rect 22569 5661 22603 5695
rect 22603 5661 22612 5695
rect 22560 5652 22612 5661
rect 23388 5720 23440 5772
rect 27988 5788 28040 5840
rect 29460 5788 29512 5840
rect 29920 5831 29972 5840
rect 29920 5797 29929 5831
rect 29929 5797 29963 5831
rect 29963 5797 29972 5831
rect 29920 5788 29972 5797
rect 30012 5788 30064 5840
rect 20168 5584 20220 5636
rect 20812 5584 20864 5636
rect 23848 5695 23900 5704
rect 23848 5661 23857 5695
rect 23857 5661 23891 5695
rect 23891 5661 23900 5695
rect 23848 5652 23900 5661
rect 23940 5695 23992 5704
rect 23940 5661 23949 5695
rect 23949 5661 23983 5695
rect 23983 5661 23992 5695
rect 23940 5652 23992 5661
rect 24124 5652 24176 5704
rect 24952 5652 25004 5704
rect 25688 5652 25740 5704
rect 27620 5652 27672 5704
rect 28080 5695 28132 5704
rect 28080 5661 28089 5695
rect 28089 5661 28123 5695
rect 28123 5661 28132 5695
rect 28080 5652 28132 5661
rect 29460 5652 29512 5704
rect 29920 5652 29972 5704
rect 30840 5652 30892 5704
rect 31944 5695 31996 5704
rect 31944 5661 31953 5695
rect 31953 5661 31987 5695
rect 31987 5661 31996 5695
rect 31944 5652 31996 5661
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 22836 5559 22888 5568
rect 22836 5525 22845 5559
rect 22845 5525 22879 5559
rect 22879 5525 22888 5559
rect 22836 5516 22888 5525
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 24676 5559 24728 5568
rect 24676 5525 24685 5559
rect 24685 5525 24719 5559
rect 24719 5525 24728 5559
rect 24676 5516 24728 5525
rect 30748 5627 30800 5636
rect 30748 5593 30757 5627
rect 30757 5593 30791 5627
rect 30791 5593 30800 5627
rect 30748 5584 30800 5593
rect 27436 5516 27488 5568
rect 29736 5516 29788 5568
rect 30380 5516 30432 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 7288 5312 7340 5364
rect 7472 5312 7524 5364
rect 6092 5176 6144 5228
rect 8208 5312 8260 5364
rect 9036 5312 9088 5364
rect 8484 5176 8536 5228
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 10048 5244 10100 5296
rect 12532 5312 12584 5364
rect 9404 5176 9456 5228
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 10876 5176 10928 5228
rect 12256 5219 12308 5228
rect 9312 5040 9364 5092
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 13636 5312 13688 5364
rect 14464 5355 14516 5364
rect 14464 5321 14473 5355
rect 14473 5321 14507 5355
rect 14507 5321 14516 5355
rect 14464 5312 14516 5321
rect 13084 5244 13136 5296
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 12164 5108 12216 5160
rect 13728 5176 13780 5228
rect 15292 5312 15344 5364
rect 15476 5312 15528 5364
rect 19340 5312 19392 5364
rect 15108 5176 15160 5228
rect 16396 5176 16448 5228
rect 13452 5040 13504 5092
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 13636 4972 13688 5024
rect 16580 5244 16632 5296
rect 18328 5244 18380 5296
rect 19248 5244 19300 5296
rect 19340 5219 19392 5228
rect 19340 5185 19349 5219
rect 19349 5185 19383 5219
rect 19383 5185 19392 5219
rect 19340 5176 19392 5185
rect 19984 5244 20036 5296
rect 20168 5244 20220 5296
rect 28172 5312 28224 5364
rect 20260 5219 20312 5228
rect 20260 5185 20269 5219
rect 20269 5185 20303 5219
rect 20303 5185 20312 5219
rect 20260 5176 20312 5185
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 23480 5244 23532 5296
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 23204 5219 23256 5228
rect 23204 5185 23213 5219
rect 23213 5185 23247 5219
rect 23247 5185 23256 5219
rect 23204 5176 23256 5185
rect 23388 5176 23440 5228
rect 24308 5287 24360 5296
rect 24308 5253 24317 5287
rect 24317 5253 24351 5287
rect 24351 5253 24360 5287
rect 24308 5244 24360 5253
rect 23848 5176 23900 5228
rect 29552 5176 29604 5228
rect 29736 5219 29788 5228
rect 29736 5185 29745 5219
rect 29745 5185 29779 5219
rect 29779 5185 29788 5219
rect 29736 5176 29788 5185
rect 30840 5312 30892 5364
rect 31944 5312 31996 5364
rect 31760 5244 31812 5296
rect 20352 5151 20404 5160
rect 20352 5117 20361 5151
rect 20361 5117 20395 5151
rect 20395 5117 20404 5151
rect 20352 5108 20404 5117
rect 20076 5040 20128 5092
rect 29828 5151 29880 5160
rect 29828 5117 29837 5151
rect 29837 5117 29871 5151
rect 29871 5117 29880 5151
rect 29828 5108 29880 5117
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 19616 4972 19668 5024
rect 20628 4972 20680 5024
rect 24952 5040 25004 5092
rect 28172 5040 28224 5092
rect 30196 5108 30248 5160
rect 30656 5176 30708 5228
rect 23940 4972 23992 5024
rect 25136 4972 25188 5024
rect 25688 4972 25740 5024
rect 29460 5015 29512 5024
rect 29460 4981 29469 5015
rect 29469 4981 29503 5015
rect 29503 4981 29512 5015
rect 29460 4972 29512 4981
rect 30380 5083 30432 5092
rect 30380 5049 30389 5083
rect 30389 5049 30423 5083
rect 30423 5049 30432 5083
rect 30380 5040 30432 5049
rect 29828 4972 29880 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 8208 4768 8260 4820
rect 8668 4768 8720 4820
rect 9036 4700 9088 4752
rect 13544 4768 13596 4820
rect 13820 4768 13872 4820
rect 15568 4768 15620 4820
rect 19156 4768 19208 4820
rect 20076 4768 20128 4820
rect 20260 4768 20312 4820
rect 21272 4768 21324 4820
rect 23204 4768 23256 4820
rect 24676 4768 24728 4820
rect 25320 4768 25372 4820
rect 25596 4768 25648 4820
rect 25688 4768 25740 4820
rect 25872 4768 25924 4820
rect 26424 4811 26476 4820
rect 26424 4777 26433 4811
rect 26433 4777 26467 4811
rect 26467 4777 26476 4811
rect 26424 4768 26476 4777
rect 6184 4632 6236 4684
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 11704 4632 11756 4684
rect 2596 4564 2648 4616
rect 8300 4564 8352 4616
rect 9312 4564 9364 4616
rect 10876 4564 10928 4616
rect 7472 4496 7524 4548
rect 940 4428 992 4480
rect 9220 4496 9272 4548
rect 11520 4428 11572 4480
rect 12440 4496 12492 4548
rect 13452 4564 13504 4616
rect 13636 4564 13688 4616
rect 19340 4632 19392 4684
rect 19616 4675 19668 4684
rect 19616 4641 19625 4675
rect 19625 4641 19659 4675
rect 19659 4641 19668 4675
rect 19616 4632 19668 4641
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 20444 4632 20496 4684
rect 21364 4632 21416 4684
rect 23388 4632 23440 4684
rect 15016 4496 15068 4548
rect 15292 4428 15344 4480
rect 20076 4428 20128 4480
rect 20352 4539 20404 4548
rect 20352 4505 20377 4539
rect 20377 4505 20404 4539
rect 20352 4496 20404 4505
rect 22928 4607 22980 4616
rect 22928 4573 22937 4607
rect 22937 4573 22971 4607
rect 22971 4573 22980 4607
rect 22928 4564 22980 4573
rect 25228 4700 25280 4752
rect 27712 4768 27764 4820
rect 28448 4768 28500 4820
rect 29460 4768 29512 4820
rect 30012 4811 30064 4820
rect 30012 4777 30021 4811
rect 30021 4777 30055 4811
rect 30055 4777 30064 4811
rect 30012 4768 30064 4777
rect 30196 4768 30248 4820
rect 30748 4768 30800 4820
rect 28080 4700 28132 4752
rect 28724 4700 28776 4752
rect 24032 4496 24084 4548
rect 25228 4607 25280 4616
rect 25228 4573 25237 4607
rect 25237 4573 25271 4607
rect 25271 4573 25280 4607
rect 25228 4564 25280 4573
rect 25504 4564 25556 4616
rect 25596 4607 25648 4616
rect 25596 4573 25605 4607
rect 25605 4573 25639 4607
rect 25639 4573 25648 4607
rect 25596 4564 25648 4573
rect 27068 4632 27120 4684
rect 25964 4607 26016 4616
rect 25964 4573 25973 4607
rect 25973 4573 26007 4607
rect 26007 4573 26016 4607
rect 25964 4564 26016 4573
rect 26792 4607 26844 4616
rect 26792 4573 26801 4607
rect 26801 4573 26835 4607
rect 26835 4573 26844 4607
rect 26792 4564 26844 4573
rect 28540 4675 28592 4684
rect 28540 4641 28549 4675
rect 28549 4641 28583 4675
rect 28583 4641 28592 4675
rect 28540 4632 28592 4641
rect 29276 4675 29328 4684
rect 29276 4641 29285 4675
rect 29285 4641 29319 4675
rect 29319 4641 29328 4675
rect 29276 4632 29328 4641
rect 29920 4564 29972 4616
rect 30656 4564 30708 4616
rect 26516 4496 26568 4548
rect 26884 4496 26936 4548
rect 27436 4539 27488 4548
rect 27436 4505 27445 4539
rect 27445 4505 27479 4539
rect 27479 4505 27488 4539
rect 27436 4496 27488 4505
rect 27896 4428 27948 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 8576 4224 8628 4276
rect 12440 4224 12492 4276
rect 13268 4224 13320 4276
rect 25136 4224 25188 4276
rect 25320 4224 25372 4276
rect 13084 4156 13136 4208
rect 8300 4088 8352 4140
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 20444 4088 20496 4140
rect 20628 4088 20680 4140
rect 24032 4156 24084 4208
rect 25872 4156 25924 4208
rect 25964 4020 26016 4072
rect 24032 3952 24084 4004
rect 25504 3952 25556 4004
rect 26792 4224 26844 4276
rect 27068 4224 27120 4276
rect 27436 4224 27488 4276
rect 27896 4224 27948 4276
rect 28080 4224 28132 4276
rect 26424 4156 26476 4208
rect 26516 4156 26568 4208
rect 27712 4156 27764 4208
rect 28540 4267 28592 4276
rect 28540 4233 28549 4267
rect 28549 4233 28583 4267
rect 28583 4233 28592 4267
rect 28540 4224 28592 4233
rect 27988 4131 28040 4140
rect 27988 4097 27997 4131
rect 27997 4097 28031 4131
rect 28031 4097 28040 4131
rect 27988 4088 28040 4097
rect 28172 4088 28224 4140
rect 29552 4088 29604 4140
rect 26884 4020 26936 4072
rect 27344 3952 27396 4004
rect 22928 3884 22980 3936
rect 28632 3884 28684 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 16488 3136 16540 3188
rect 17684 3136 17736 3188
rect 36912 3136 36964 3188
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 25412 3000 25464 3052
rect 8208 2796 8260 2848
rect 12992 2839 13044 2848
rect 12992 2805 13001 2839
rect 13001 2805 13035 2839
rect 13035 2805 13044 2839
rect 12992 2796 13044 2805
rect 16212 2839 16264 2848
rect 16212 2805 16221 2839
rect 16221 2805 16255 2839
rect 16255 2805 16264 2839
rect 16212 2796 16264 2805
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 17408 2796 17460 2805
rect 21916 2796 21968 2848
rect 37188 2796 37240 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 10232 2456 10284 2508
rect 1492 2431 1544 2440
rect 1492 2397 1501 2431
rect 1501 2397 1535 2431
rect 1535 2397 1544 2431
rect 1492 2388 1544 2397
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 8208 2388 8260 2440
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 9588 2388 9640 2440
rect 11152 2363 11204 2372
rect 11152 2329 11161 2363
rect 11161 2329 11195 2363
rect 11195 2329 11204 2363
rect 11152 2320 11204 2329
rect 12992 2388 13044 2440
rect 16212 2388 16264 2440
rect 17408 2388 17460 2440
rect 21916 2388 21968 2440
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 20 2252 72 2304
rect 1952 2252 2004 2304
rect 3976 2252 4028 2304
rect 6828 2252 6880 2304
rect 12900 2252 12952 2304
rect 15016 2252 15068 2304
rect 17408 2252 17460 2304
rect 19340 2252 19392 2304
rect 26424 2252 26476 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 18 40762 74 41562
rect 1950 40762 2006 41562
rect 4526 40762 4582 41562
rect 6458 40762 6514 41562
rect 9034 40762 9090 41562
rect 10966 40762 11022 41562
rect 12898 40762 12954 41562
rect 15474 40762 15530 41562
rect 17406 40762 17462 41562
rect 19982 40762 20038 41562
rect 21914 40762 21970 41562
rect 24490 40762 24546 41562
rect 26422 40762 26478 41562
rect 28354 40762 28410 41562
rect 30930 40762 30986 41562
rect 32862 40762 32918 41562
rect 35438 40882 35494 41562
rect 35438 40854 35848 40882
rect 35438 40762 35494 40854
rect 32 39098 60 40762
rect 4540 39098 4568 40762
rect 9048 39098 9076 40762
rect 10980 39114 11008 40762
rect 10980 39098 11100 39114
rect 12912 39098 12940 40762
rect 20 39092 72 39098
rect 20 39034 72 39040
rect 4528 39092 4580 39098
rect 4528 39034 4580 39040
rect 9036 39092 9088 39098
rect 10980 39092 11112 39098
rect 10980 39086 11060 39092
rect 9036 39034 9088 39040
rect 11060 39034 11112 39040
rect 12900 39092 12952 39098
rect 12900 39034 12952 39040
rect 15488 39030 15516 40762
rect 17420 39098 17448 40762
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 17408 39092 17460 39098
rect 17408 39034 17460 39040
rect 9128 39024 9180 39030
rect 9128 38966 9180 38972
rect 15476 39024 15528 39030
rect 15476 38966 15528 38972
rect 16028 39024 16080 39030
rect 16028 38966 16080 38972
rect 3792 38956 3844 38962
rect 3792 38898 3844 38904
rect 4804 38956 4856 38962
rect 4804 38898 4856 38904
rect 940 37188 992 37194
rect 940 37130 992 37136
rect 952 36825 980 37130
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 1768 28416 1820 28422
rect 1768 28358 1820 28364
rect 1780 26234 1808 28358
rect 1780 26206 1900 26234
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1582 24984 1638 24993
rect 1582 24919 1584 24928
rect 1636 24919 1638 24928
rect 1584 24890 1636 24896
rect 1688 24886 1716 25230
rect 1676 24880 1728 24886
rect 1676 24822 1728 24828
rect 1492 24812 1544 24818
rect 1492 24754 1544 24760
rect 1504 22778 1532 24754
rect 1688 23798 1716 24822
rect 1676 23792 1728 23798
rect 1676 23734 1728 23740
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 1688 21146 1716 23734
rect 1768 23656 1820 23662
rect 1768 23598 1820 23604
rect 1780 23322 1808 23598
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1872 23202 1900 26206
rect 1952 25220 2004 25226
rect 1952 25162 2004 25168
rect 1964 24954 1992 25162
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 1952 24948 2004 24954
rect 1952 24890 2004 24896
rect 2792 24886 2820 25094
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 1780 23174 1900 23202
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1688 20602 1716 20810
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 952 20505 980 20538
rect 1780 20534 1808 23174
rect 2792 23066 2820 24822
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3700 24744 3752 24750
rect 3700 24686 3752 24692
rect 2884 23322 2912 24686
rect 3160 24138 3188 24686
rect 3712 24410 3740 24686
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3148 24132 3200 24138
rect 3148 24074 3200 24080
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 3160 23186 3188 24074
rect 3332 23520 3384 23526
rect 3332 23462 3384 23468
rect 3148 23180 3200 23186
rect 3148 23122 3200 23128
rect 2700 23038 2820 23066
rect 2700 22778 2728 23038
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 2792 22778 2820 22918
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 3054 22672 3110 22681
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2596 22636 2648 22642
rect 2596 22578 2648 22584
rect 2780 22636 2832 22642
rect 3054 22607 3056 22616
rect 2780 22578 2832 22584
rect 3108 22607 3110 22616
rect 3056 22578 3108 22584
rect 2516 21622 2544 22578
rect 2608 21690 2636 22578
rect 2792 22094 2820 22578
rect 3160 22094 3188 23122
rect 3344 23118 3372 23462
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3252 22098 3280 22374
rect 3344 22166 3372 23054
rect 3608 23044 3660 23050
rect 3608 22986 3660 22992
rect 3620 22778 3648 22986
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3528 22234 3556 22578
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3332 22160 3384 22166
rect 3332 22102 3384 22108
rect 2792 22066 2912 22094
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2504 21616 2556 21622
rect 2410 21584 2466 21593
rect 2504 21558 2556 21564
rect 2410 21519 2412 21528
rect 2464 21519 2466 21528
rect 2412 21490 2464 21496
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2226 20632 2282 20641
rect 2516 20602 2544 21286
rect 2226 20567 2282 20576
rect 2504 20596 2556 20602
rect 1768 20528 1820 20534
rect 938 20496 994 20505
rect 1768 20470 1820 20476
rect 2240 20466 2268 20567
rect 2504 20538 2556 20544
rect 938 20431 994 20440
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 940 18624 992 18630
rect 940 18566 992 18572
rect 952 18465 980 18566
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 952 15745 980 15846
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 1412 15570 1440 17138
rect 1504 16182 1532 20198
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2700 19514 2728 19654
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1780 18766 1808 19110
rect 1964 18970 1992 19314
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2056 18766 2084 19110
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2424 18426 2452 19110
rect 2884 18680 2912 22066
rect 3068 22066 3188 22094
rect 3240 22092 3292 22098
rect 3068 21486 3096 22066
rect 3240 22034 3292 22040
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 2976 20602 3004 21422
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2964 18692 3016 18698
rect 2884 18652 2964 18680
rect 2964 18634 3016 18640
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2792 18426 2820 18566
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 1688 16794 1716 17070
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1492 16176 1544 16182
rect 1492 16118 1544 16124
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1676 15428 1728 15434
rect 1676 15370 1728 15376
rect 1688 15162 1716 15370
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 938 13696 994 13705
rect 938 13631 994 13640
rect 952 13530 980 13631
rect 940 13524 992 13530
rect 940 13466 992 13472
rect 1412 12374 1440 13806
rect 1688 13530 1716 13806
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1400 12368 1452 12374
rect 1400 12310 1452 12316
rect 1412 11762 1440 12310
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 11898 1808 12038
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 952 11150 980 11591
rect 940 11144 992 11150
rect 940 11086 992 11092
rect 1412 10606 1440 11698
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 9586 1440 10542
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1504 8974 1532 9862
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9178 1716 9454
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1492 8968 1544 8974
rect 938 8936 994 8945
rect 1492 8910 1544 8916
rect 938 8871 994 8880
rect 952 8838 980 8871
rect 940 8832 992 8838
rect 940 8774 992 8780
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6905 1532 7346
rect 1964 6914 1992 18022
rect 2332 6914 2360 18022
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2516 16794 2544 17478
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2792 15502 2820 17138
rect 2884 16998 2912 17478
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2976 16810 3004 18634
rect 3068 17746 3096 21422
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3160 19854 3188 20946
rect 3712 20890 3740 22646
rect 3240 20868 3292 20874
rect 3240 20810 3292 20816
rect 3620 20862 3740 20890
rect 3252 20398 3280 20810
rect 3620 20602 3648 20862
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3712 20466 3740 20742
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3252 19786 3280 20334
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 18873 3188 19654
rect 3804 18970 3832 38898
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4816 38554 4844 38898
rect 4804 38548 4856 38554
rect 4804 38490 4856 38496
rect 5170 38448 5226 38457
rect 5170 38383 5226 38392
rect 5184 38350 5212 38383
rect 5172 38344 5224 38350
rect 5172 38286 5224 38292
rect 6458 38312 6514 38321
rect 6458 38247 6514 38256
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 6472 37330 6500 38247
rect 7104 38208 7156 38214
rect 7104 38150 7156 38156
rect 8576 38208 8628 38214
rect 8576 38150 8628 38156
rect 6460 37324 6512 37330
rect 6460 37266 6512 37272
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 5540 36100 5592 36106
rect 5540 36042 5592 36048
rect 5356 36032 5408 36038
rect 5356 35974 5408 35980
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4528 34944 4580 34950
rect 4528 34886 4580 34892
rect 4540 34746 4568 34886
rect 4528 34740 4580 34746
rect 4528 34682 4580 34688
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 34202 4660 34478
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4528 33856 4580 33862
rect 4528 33798 4580 33804
rect 4540 33658 4568 33798
rect 4528 33652 4580 33658
rect 4528 33594 4580 33600
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 33114 4660 33390
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 5368 32434 5396 35974
rect 5552 35834 5580 36042
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 6472 35766 6500 37266
rect 7116 36718 7144 38150
rect 8588 38010 8616 38150
rect 8576 38004 8628 38010
rect 8576 37946 8628 37952
rect 8668 37800 8720 37806
rect 8668 37742 8720 37748
rect 8680 37466 8708 37742
rect 8668 37460 8720 37466
rect 8668 37402 8720 37408
rect 7104 36712 7156 36718
rect 7104 36654 7156 36660
rect 7012 36576 7064 36582
rect 7012 36518 7064 36524
rect 7024 36378 7052 36518
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 6828 36100 6880 36106
rect 6828 36042 6880 36048
rect 6736 36032 6788 36038
rect 6736 35974 6788 35980
rect 5632 35760 5684 35766
rect 5632 35702 5684 35708
rect 6460 35760 6512 35766
rect 6460 35702 6512 35708
rect 5448 35080 5500 35086
rect 5448 35022 5500 35028
rect 5460 33998 5488 35022
rect 5448 33992 5500 33998
rect 5448 33934 5500 33940
rect 5356 32428 5408 32434
rect 5356 32370 5408 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3884 31816 3936 31822
rect 3884 31758 3936 31764
rect 3896 31482 3924 31758
rect 4160 31748 4212 31754
rect 4160 31690 4212 31696
rect 4172 31482 4200 31690
rect 3884 31476 3936 31482
rect 3884 31418 3936 31424
rect 4160 31476 4212 31482
rect 4160 31418 4212 31424
rect 5368 31346 5396 32370
rect 5460 31754 5488 33934
rect 5644 31754 5672 35702
rect 5724 35692 5776 35698
rect 5724 35634 5776 35640
rect 5736 35290 5764 35634
rect 5724 35284 5776 35290
rect 5724 35226 5776 35232
rect 6552 35148 6604 35154
rect 6552 35090 6604 35096
rect 6460 34944 6512 34950
rect 6460 34886 6512 34892
rect 6472 34746 6500 34886
rect 6460 34740 6512 34746
rect 6460 34682 6512 34688
rect 6368 34400 6420 34406
rect 6368 34342 6420 34348
rect 6380 33998 6408 34342
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6184 33312 6236 33318
rect 6184 33254 6236 33260
rect 6196 32774 6224 33254
rect 6184 32768 6236 32774
rect 6184 32710 6236 32716
rect 6196 32502 6224 32710
rect 6184 32496 6236 32502
rect 6184 32438 6236 32444
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 5460 31726 5580 31754
rect 5644 31726 5764 31754
rect 5552 31346 5580 31726
rect 5356 31340 5408 31346
rect 5356 31282 5408 31288
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4528 29504 4580 29510
rect 4528 29446 4580 29452
rect 4540 29306 4568 29446
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4988 28960 5040 28966
rect 4988 28902 5040 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5000 28762 5028 28902
rect 4988 28756 5040 28762
rect 4988 28698 5040 28704
rect 5368 28558 5396 31282
rect 5736 29646 5764 31726
rect 5828 31482 5856 31758
rect 6564 31754 6592 35090
rect 6748 35018 6776 35974
rect 6840 35630 6868 36042
rect 6828 35624 6880 35630
rect 6828 35566 6880 35572
rect 6736 35012 6788 35018
rect 6736 34954 6788 34960
rect 6736 34604 6788 34610
rect 6840 34592 6868 35566
rect 6788 34564 6868 34592
rect 6736 34546 6788 34552
rect 6644 34468 6696 34474
rect 6644 34410 6696 34416
rect 6656 32978 6684 34410
rect 6840 33590 6868 34564
rect 7116 33998 7144 36654
rect 8944 36168 8996 36174
rect 8944 36110 8996 36116
rect 7196 36100 7248 36106
rect 7196 36042 7248 36048
rect 8484 36100 8536 36106
rect 8484 36042 8536 36048
rect 7208 35834 7236 36042
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 8496 35766 8524 36042
rect 8668 36032 8720 36038
rect 8668 35974 8720 35980
rect 8680 35834 8708 35974
rect 8956 35834 8984 36110
rect 8668 35828 8720 35834
rect 8668 35770 8720 35776
rect 8944 35828 8996 35834
rect 8944 35770 8996 35776
rect 8484 35760 8536 35766
rect 8484 35702 8536 35708
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 8024 34944 8076 34950
rect 8024 34886 8076 34892
rect 8036 34678 8064 34886
rect 8024 34672 8076 34678
rect 8024 34614 8076 34620
rect 7748 34536 7800 34542
rect 7748 34478 7800 34484
rect 8116 34536 8168 34542
rect 8116 34478 8168 34484
rect 7760 34066 7788 34478
rect 8128 34202 8156 34478
rect 8116 34196 8168 34202
rect 8116 34138 8168 34144
rect 8220 34082 8248 35430
rect 8680 35290 8708 35770
rect 8944 35624 8996 35630
rect 8944 35566 8996 35572
rect 8668 35284 8720 35290
rect 8668 35226 8720 35232
rect 8956 34746 8984 35566
rect 8944 34740 8996 34746
rect 8944 34682 8996 34688
rect 7748 34060 7800 34066
rect 7748 34002 7800 34008
rect 8128 34054 8248 34082
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 7208 33658 7236 33798
rect 7196 33652 7248 33658
rect 7196 33594 7248 33600
rect 6828 33584 6880 33590
rect 6828 33526 6880 33532
rect 6840 33266 6868 33526
rect 7288 33448 7340 33454
rect 7288 33390 7340 33396
rect 6840 33238 6960 33266
rect 6644 32972 6696 32978
rect 6644 32914 6696 32920
rect 6472 31726 6592 31754
rect 5816 31476 5868 31482
rect 5816 31418 5868 31424
rect 6472 31278 6500 31726
rect 6656 31498 6684 32914
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 6748 31686 6776 32302
rect 6828 32020 6880 32026
rect 6932 32008 6960 33238
rect 7300 33114 7328 33390
rect 8128 33114 8156 34054
rect 8208 33924 8260 33930
rect 8208 33866 8260 33872
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 8116 32972 8168 32978
rect 8116 32914 8168 32920
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 6880 31980 6960 32008
rect 6828 31962 6880 31968
rect 6736 31680 6788 31686
rect 6736 31622 6788 31628
rect 6564 31470 6684 31498
rect 6748 31482 6776 31622
rect 6736 31476 6788 31482
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 6368 30592 6420 30598
rect 6368 30534 6420 30540
rect 6380 30190 6408 30534
rect 6368 30184 6420 30190
rect 6368 30126 6420 30132
rect 5724 29640 5776 29646
rect 5724 29582 5776 29588
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4356 28218 4384 28358
rect 4344 28212 4396 28218
rect 4344 28154 4396 28160
rect 4712 28144 4764 28150
rect 4712 28086 4764 28092
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4724 27674 4752 28086
rect 4712 27668 4764 27674
rect 4712 27610 4764 27616
rect 4066 27296 4122 27305
rect 4066 27231 4122 27240
rect 4080 26450 4108 27231
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5368 26586 5396 28494
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 5368 26330 5396 26522
rect 5276 26314 5396 26330
rect 5460 26314 5488 26726
rect 5264 26308 5396 26314
rect 5316 26302 5396 26308
rect 5448 26308 5500 26314
rect 5264 26250 5316 26256
rect 5448 26250 5500 26256
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 5644 25498 5672 25638
rect 5632 25492 5684 25498
rect 5632 25434 5684 25440
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 4080 24750 4108 25162
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 4080 23798 4108 24686
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4816 24206 4844 24550
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 4160 23112 4212 23118
rect 4620 23112 4672 23118
rect 4160 23054 4212 23060
rect 4618 23080 4620 23089
rect 4672 23080 4674 23089
rect 4816 23066 4844 23122
rect 3988 22778 4016 23054
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 4172 22710 4200 23054
rect 4344 23044 4396 23050
rect 4618 23015 4674 23024
rect 4724 23038 4844 23066
rect 4344 22986 4396 22992
rect 4160 22704 4212 22710
rect 4066 22672 4122 22681
rect 3976 22636 4028 22642
rect 4160 22646 4212 22652
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4066 22607 4068 22616
rect 3976 22578 4028 22584
rect 4120 22607 4122 22616
rect 4068 22578 4120 22584
rect 3988 22137 4016 22578
rect 4264 22438 4292 22646
rect 4356 22574 4384 22986
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4344 22568 4396 22574
rect 4344 22510 4396 22516
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3974 22128 4030 22137
rect 3974 22063 4030 22072
rect 3884 21956 3936 21962
rect 3884 21898 3936 21904
rect 3896 21554 3924 21898
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3896 21010 3924 21490
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3988 20482 4016 21490
rect 4172 21332 4200 21830
rect 4540 21554 4568 21830
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4080 21304 4200 21332
rect 4080 21128 4108 21304
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21146 4660 22578
rect 4620 21140 4672 21146
rect 4080 21100 4200 21128
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4080 20584 4108 20946
rect 4172 20874 4200 21100
rect 4620 21082 4672 21088
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 4080 20556 4292 20584
rect 3896 20454 4016 20482
rect 4066 20496 4122 20505
rect 4264 20466 4292 20556
rect 4448 20534 4476 20742
rect 4436 20528 4488 20534
rect 4436 20470 4488 20476
rect 3896 19922 3924 20454
rect 4066 20431 4068 20440
rect 4120 20431 4122 20440
rect 4252 20460 4304 20466
rect 4068 20402 4120 20408
rect 4252 20402 4304 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3896 19718 3924 19858
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3146 18864 3202 18873
rect 3146 18799 3202 18808
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3252 18290 3280 18770
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3528 18426 3556 18702
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3896 18222 3924 19654
rect 4172 19334 4200 19790
rect 4724 19514 4752 23038
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4816 22030 4844 22374
rect 4908 22098 4936 24006
rect 4988 23044 5040 23050
rect 4988 22986 5040 22992
rect 5080 23044 5132 23050
rect 5080 22986 5132 22992
rect 5000 22166 5028 22986
rect 5092 22778 5120 22986
rect 5080 22772 5132 22778
rect 5080 22714 5132 22720
rect 4988 22160 5040 22166
rect 4988 22102 5040 22108
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4804 22024 4856 22030
rect 5000 21978 5028 22102
rect 4804 21966 4856 21972
rect 4908 21950 5028 21978
rect 4908 20602 4936 21950
rect 4988 21888 5040 21894
rect 4986 21856 4988 21865
rect 5040 21856 5042 21865
rect 4986 21791 5042 21800
rect 5276 21622 5304 24550
rect 5460 24274 5488 24686
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 5460 23186 5488 24210
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 5644 22030 5672 23122
rect 5736 22094 5764 29582
rect 6276 29572 6328 29578
rect 6276 29514 6328 29520
rect 6288 29170 6316 29514
rect 6564 29458 6592 31470
rect 6736 31418 6788 31424
rect 7484 31346 7512 32166
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 7748 31680 7800 31686
rect 7748 31622 7800 31628
rect 7760 31414 7788 31622
rect 7852 31414 7880 31962
rect 8024 31952 8076 31958
rect 8024 31894 8076 31900
rect 7748 31408 7800 31414
rect 7748 31350 7800 31356
rect 7840 31408 7892 31414
rect 7840 31350 7892 31356
rect 6644 31340 6696 31346
rect 6644 31282 6696 31288
rect 7472 31340 7524 31346
rect 7472 31282 7524 31288
rect 6656 30598 6684 31282
rect 6828 31272 6880 31278
rect 6828 31214 6880 31220
rect 6840 30802 6868 31214
rect 8036 30938 8064 31894
rect 8128 31482 8156 32914
rect 8220 32026 8248 33866
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 8772 32910 8800 33254
rect 8956 32910 8984 34682
rect 8760 32904 8812 32910
rect 8760 32846 8812 32852
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 8772 32570 8800 32846
rect 8852 32836 8904 32842
rect 8852 32778 8904 32784
rect 8760 32564 8812 32570
rect 8760 32506 8812 32512
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8668 31680 8720 31686
rect 8668 31622 8720 31628
rect 8116 31476 8168 31482
rect 8116 31418 8168 31424
rect 8024 30932 8076 30938
rect 8024 30874 8076 30880
rect 6828 30796 6880 30802
rect 6828 30738 6880 30744
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 6656 29646 6684 30534
rect 6644 29640 6696 29646
rect 6644 29582 6696 29588
rect 6564 29430 6684 29458
rect 6276 29164 6328 29170
rect 6276 29106 6328 29112
rect 6288 28150 6316 29106
rect 6656 29102 6684 29430
rect 6736 29164 6788 29170
rect 6736 29106 6788 29112
rect 6644 29096 6696 29102
rect 6644 29038 6696 29044
rect 6368 28960 6420 28966
rect 6368 28902 6420 28908
rect 6380 28626 6408 28902
rect 6368 28620 6420 28626
rect 6368 28562 6420 28568
rect 6276 28144 6328 28150
rect 6276 28086 6328 28092
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5920 27470 5948 27814
rect 5908 27464 5960 27470
rect 5908 27406 5960 27412
rect 6748 27402 6776 29106
rect 6840 27538 6868 30738
rect 8128 30682 8156 31418
rect 8680 30734 8708 31622
rect 7944 30666 8156 30682
rect 8208 30728 8260 30734
rect 8208 30670 8260 30676
rect 8668 30728 8720 30734
rect 8864 30716 8892 32778
rect 8944 31884 8996 31890
rect 8944 31826 8996 31832
rect 8956 30938 8984 31826
rect 9140 31754 9168 38966
rect 9312 38956 9364 38962
rect 9312 38898 9364 38904
rect 11612 38956 11664 38962
rect 11612 38898 11664 38904
rect 11980 38956 12032 38962
rect 11980 38898 12032 38904
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 12992 38956 13044 38962
rect 12992 38898 13044 38904
rect 9324 38554 9352 38898
rect 11244 38888 11296 38894
rect 11244 38830 11296 38836
rect 10232 38820 10284 38826
rect 10232 38762 10284 38768
rect 9312 38548 9364 38554
rect 9312 38490 9364 38496
rect 9496 38344 9548 38350
rect 9496 38286 9548 38292
rect 9220 36100 9272 36106
rect 9220 36042 9272 36048
rect 9232 35834 9260 36042
rect 9220 35828 9272 35834
rect 9220 35770 9272 35776
rect 9404 34944 9456 34950
rect 9404 34886 9456 34892
rect 9416 34678 9444 34886
rect 9404 34672 9456 34678
rect 9404 34614 9456 34620
rect 9220 34604 9272 34610
rect 9220 34546 9272 34552
rect 9232 33590 9260 34546
rect 9220 33584 9272 33590
rect 9220 33526 9272 33532
rect 9508 33386 9536 38286
rect 10140 37664 10192 37670
rect 10140 37606 10192 37612
rect 10152 37330 10180 37606
rect 10048 37324 10100 37330
rect 10048 37266 10100 37272
rect 10140 37324 10192 37330
rect 10140 37266 10192 37272
rect 9956 35692 10008 35698
rect 9956 35634 10008 35640
rect 9968 35086 9996 35634
rect 9956 35080 10008 35086
rect 9956 35022 10008 35028
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 9692 33998 9720 34682
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9772 33856 9824 33862
rect 9772 33798 9824 33804
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 9784 33538 9812 33798
rect 9876 33658 9904 33798
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 9784 33510 9904 33538
rect 9772 33448 9824 33454
rect 9772 33390 9824 33396
rect 9496 33380 9548 33386
rect 9496 33322 9548 33328
rect 9784 33114 9812 33390
rect 9772 33108 9824 33114
rect 9772 33050 9824 33056
rect 9496 32904 9548 32910
rect 9496 32846 9548 32852
rect 9404 32768 9456 32774
rect 9404 32710 9456 32716
rect 9416 31958 9444 32710
rect 9404 31952 9456 31958
rect 9404 31894 9456 31900
rect 9048 31726 9168 31754
rect 9508 31754 9536 32846
rect 9508 31726 9628 31754
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 8944 30728 8996 30734
rect 8864 30688 8944 30716
rect 8668 30670 8720 30676
rect 8944 30670 8996 30676
rect 7932 30660 8156 30666
rect 7984 30654 8156 30660
rect 7932 30602 7984 30608
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7668 29238 7696 29446
rect 7656 29232 7708 29238
rect 7656 29174 7708 29180
rect 7380 29096 7432 29102
rect 7380 29038 7432 29044
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7840 29096 7892 29102
rect 7840 29038 7892 29044
rect 6920 28416 6972 28422
rect 6920 28358 6972 28364
rect 6932 28218 6960 28358
rect 6920 28212 6972 28218
rect 6920 28154 6972 28160
rect 7012 28008 7064 28014
rect 7012 27950 7064 27956
rect 7024 27674 7052 27950
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6736 27396 6788 27402
rect 6736 27338 6788 27344
rect 6840 27130 6868 27474
rect 6828 27124 6880 27130
rect 6828 27066 6880 27072
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 5920 26042 5948 26930
rect 6644 26376 6696 26382
rect 6644 26318 6696 26324
rect 5908 26036 5960 26042
rect 5908 25978 5960 25984
rect 6000 25900 6052 25906
rect 6000 25842 6052 25848
rect 6012 25498 6040 25842
rect 6000 25492 6052 25498
rect 6000 25434 6052 25440
rect 6656 25294 6684 26318
rect 6840 25838 6868 27066
rect 7392 26790 7420 29038
rect 7760 28762 7788 29038
rect 7748 28756 7800 28762
rect 7748 28698 7800 28704
rect 7852 28694 7880 29038
rect 7840 28688 7892 28694
rect 7840 28630 7892 28636
rect 7944 28506 7972 30602
rect 8024 30252 8076 30258
rect 8024 30194 8076 30200
rect 8036 29782 8064 30194
rect 8220 30054 8248 30670
rect 8484 30660 8536 30666
rect 8484 30602 8536 30608
rect 8496 30326 8524 30602
rect 8760 30592 8812 30598
rect 8760 30534 8812 30540
rect 8772 30394 8800 30534
rect 8760 30388 8812 30394
rect 8760 30330 8812 30336
rect 8484 30320 8536 30326
rect 8484 30262 8536 30268
rect 8956 30258 8984 30670
rect 8944 30252 8996 30258
rect 8944 30194 8996 30200
rect 8208 30048 8260 30054
rect 8208 29990 8260 29996
rect 8024 29776 8076 29782
rect 8024 29718 8076 29724
rect 8036 28778 8064 29718
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8036 28750 8156 28778
rect 8024 28620 8076 28626
rect 8024 28562 8076 28568
rect 7852 28478 7972 28506
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7748 26784 7800 26790
rect 7748 26726 7800 26732
rect 7104 26444 7156 26450
rect 7104 26386 7156 26392
rect 6828 25832 6880 25838
rect 6828 25774 6880 25780
rect 6644 25288 6696 25294
rect 6644 25230 6696 25236
rect 6656 24886 6684 25230
rect 6644 24880 6696 24886
rect 6644 24822 6696 24828
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 6196 23118 6224 24754
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6748 23866 6776 24074
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6736 23860 6788 23866
rect 6736 23802 6788 23808
rect 6932 23662 6960 24006
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6368 23248 6420 23254
rect 6368 23190 6420 23196
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 5736 22066 5856 22094
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 5552 21434 5580 21898
rect 5552 21406 5672 21434
rect 5540 21344 5592 21350
rect 5644 21332 5672 21406
rect 5724 21344 5776 21350
rect 5644 21304 5724 21332
rect 5540 21286 5592 21292
rect 5724 21286 5776 21292
rect 5552 21146 5580 21286
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5632 20936 5684 20942
rect 5460 20896 5632 20924
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4080 19306 4200 19334
rect 4080 18748 4108 19306
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18970 4660 19246
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4160 18760 4212 18766
rect 4080 18720 4160 18748
rect 4160 18702 4212 18708
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4172 18290 4200 18702
rect 4264 18426 4292 18702
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 2884 16782 3004 16810
rect 3068 16794 3096 17682
rect 3056 16788 3108 16794
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2792 13938 2820 15438
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2884 13818 2912 16782
rect 3056 16730 3108 16736
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2976 15162 3004 15642
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 3068 14958 3096 16730
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15162 3832 15302
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3896 15026 3924 18158
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3988 17270 4016 17614
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 4080 17218 4108 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4252 17740 4304 17746
rect 4304 17700 4384 17728
rect 4252 17682 4304 17688
rect 4080 17190 4200 17218
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 3988 16114 4016 17002
rect 4080 16114 4108 17070
rect 4172 17066 4200 17190
rect 4356 17116 4384 17700
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4448 17241 4476 17614
rect 4908 17610 4936 20402
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4896 17604 4948 17610
rect 4896 17546 4948 17552
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 4712 17264 4764 17270
rect 4434 17232 4490 17241
rect 4712 17206 4764 17212
rect 4434 17167 4490 17176
rect 4356 17088 4660 17116
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4540 16114 4568 16594
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 3988 15706 4016 16050
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2792 13790 2912 13818
rect 2964 13796 3016 13802
rect 2792 12434 2820 13790
rect 2964 13738 3016 13744
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2884 12986 2912 13670
rect 2976 13394 3004 13738
rect 3068 13394 3096 14894
rect 4080 14414 4108 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 17088
rect 4724 16726 4752 17206
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4816 16590 4844 17070
rect 4908 17066 4936 17546
rect 4896 17060 4948 17066
rect 4896 17002 4948 17008
rect 5092 16998 5120 17546
rect 5184 17338 5212 17614
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5184 16794 5212 17274
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4724 15706 4752 15914
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3804 13530 3832 14350
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 4068 14272 4120 14278
rect 4632 14226 4660 15506
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4068 14214 4120 14220
rect 3988 14074 4016 14214
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3068 13274 3096 13330
rect 3896 13326 3924 13942
rect 4080 13870 4108 14214
rect 4540 14198 4660 14226
rect 4540 13870 4568 14198
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3884 13320 3936 13326
rect 3068 13246 3280 13274
rect 3884 13262 3936 13268
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12594 2912 12718
rect 2884 12566 3004 12594
rect 2792 12406 2912 12434
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11218 2820 12106
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2884 10198 2912 12406
rect 2976 11762 3004 12566
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2976 10062 3004 11018
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2884 8634 2912 9998
rect 3068 9654 3096 13126
rect 3252 12306 3280 13246
rect 3896 12850 3924 13262
rect 4632 13190 4660 14010
rect 4724 13734 4752 14962
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 4816 14074 4844 14282
rect 4908 14074 4936 14282
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13326 4752 13670
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3436 12170 3464 12786
rect 4632 12782 4660 13126
rect 4816 12918 4844 13806
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3436 11898 3464 12106
rect 3804 12050 3832 12242
rect 3896 12238 3924 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3804 12022 3924 12050
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3252 10810 3280 10950
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3804 10470 3832 11698
rect 3896 11218 3924 12022
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11348 4120 11354
rect 3988 11308 4068 11336
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3252 10062 3280 10134
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3056 9648 3108 9654
rect 3252 9625 3280 9998
rect 3056 9590 3108 9596
rect 3238 9616 3294 9625
rect 3804 9586 3832 10406
rect 3238 9551 3294 9560
rect 3792 9580 3844 9586
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3252 8498 3280 9551
rect 3792 9522 3844 9528
rect 3896 9042 3924 11154
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8634 3556 8774
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1596 6886 1992 6914
rect 2148 6886 2360 6914
rect 1596 4570 1624 6886
rect 1504 4542 1624 4570
rect 940 4480 992 4486
rect 940 4422 992 4428
rect 952 4185 980 4422
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1504 2446 1532 4542
rect 2148 2446 2176 6886
rect 2608 4622 2636 8298
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3712 6798 3740 7142
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 3988 2774 4016 11308
rect 4068 11290 4120 11296
rect 4632 11234 4660 12718
rect 4540 11206 4660 11234
rect 4540 11150 4568 11206
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4712 11144 4764 11150
rect 4764 11092 4844 11098
rect 4712 11086 4844 11092
rect 4448 10606 4476 11086
rect 4540 10690 4568 11086
rect 4724 11070 4844 11086
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4632 10810 4660 10950
rect 4724 10810 4752 10950
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4540 10662 4660 10690
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10266 4660 10662
rect 4816 10266 4844 11070
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10538 4936 10950
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4908 10062 4936 10474
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4356 9722 4384 9998
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4448 9382 4476 9522
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4080 8974 4108 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8634 4108 8910
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4066 8528 4122 8537
rect 4066 8463 4068 8472
rect 4120 8463 4122 8472
rect 4068 8434 4120 8440
rect 4264 8378 4292 8978
rect 4632 8514 4660 9522
rect 4724 8974 4752 9998
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4816 9024 4844 9318
rect 4908 9178 4936 9318
rect 5000 9178 5028 9522
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5092 9042 5120 10610
rect 5184 10606 5212 12854
rect 5276 11354 5304 20742
rect 5460 19854 5488 20896
rect 5632 20878 5684 20884
rect 5736 19922 5764 21286
rect 5828 20262 5856 22066
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 5920 21690 5948 22034
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 6012 21622 6040 21898
rect 6000 21616 6052 21622
rect 6000 21558 6052 21564
rect 6196 21554 6224 22034
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5828 19174 5856 19790
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5920 19378 5948 19654
rect 6012 19446 6040 19654
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 6380 19378 6408 23190
rect 6932 23186 6960 23598
rect 7116 23594 7144 26386
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 7208 25974 7236 26250
rect 7196 25968 7248 25974
rect 7196 25910 7248 25916
rect 7656 25424 7708 25430
rect 7656 25366 7708 25372
rect 7668 25158 7696 25366
rect 7760 25362 7788 26726
rect 7852 25378 7880 28478
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7944 25498 7972 25638
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 8036 25430 8064 28562
rect 8128 28082 8156 28750
rect 8392 28688 8444 28694
rect 8392 28630 8444 28636
rect 8404 28558 8432 28630
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 8128 27674 8156 28018
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 8404 27470 8432 27814
rect 8496 27470 8524 29446
rect 8956 28558 8984 30194
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 8852 28484 8904 28490
rect 8852 28426 8904 28432
rect 8668 27668 8720 27674
rect 8668 27610 8720 27616
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 8312 27062 8340 27270
rect 8680 27062 8708 27610
rect 8864 27538 8892 28426
rect 8852 27532 8904 27538
rect 8852 27474 8904 27480
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 8668 27056 8720 27062
rect 8668 26998 8720 27004
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8404 26518 8432 26862
rect 8392 26512 8444 26518
rect 8392 26454 8444 26460
rect 8680 26450 8708 26998
rect 8668 26444 8720 26450
rect 8668 26386 8720 26392
rect 8298 26344 8354 26353
rect 8298 26279 8354 26288
rect 8024 25424 8076 25430
rect 7748 25356 7800 25362
rect 7852 25350 7972 25378
rect 8024 25366 8076 25372
rect 7748 25298 7800 25304
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 7668 24954 7696 25094
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7852 24750 7880 25094
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7576 23730 7604 24006
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7288 23248 7340 23254
rect 7208 23208 7288 23236
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 7012 23044 7064 23050
rect 7012 22986 7064 22992
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 6656 22778 6684 22918
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6748 22642 6776 22918
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6642 22536 6698 22545
rect 6642 22471 6698 22480
rect 6656 22166 6684 22471
rect 6932 22234 6960 22578
rect 7024 22234 7052 22986
rect 7208 22778 7236 23208
rect 7288 23190 7340 23196
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7116 22545 7144 22578
rect 7102 22536 7158 22545
rect 7392 22522 7420 22646
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7102 22471 7158 22480
rect 7208 22494 7420 22522
rect 7208 22438 7236 22494
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7012 22228 7064 22234
rect 7012 22170 7064 22176
rect 6644 22160 6696 22166
rect 6696 22120 6776 22148
rect 6644 22102 6696 22108
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 21622 6684 21830
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6642 20496 6698 20505
rect 6564 20454 6642 20482
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5356 18692 5408 18698
rect 5408 18652 5580 18680
rect 5356 18634 5408 18640
rect 5552 18057 5580 18652
rect 5538 18048 5594 18057
rect 5538 17983 5594 17992
rect 5920 17898 5948 19314
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18630 6040 19110
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 5920 17870 6040 17898
rect 6012 17610 6040 17870
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 17338 5488 17478
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5460 16561 5488 16934
rect 5552 16726 5580 16934
rect 5828 16726 5856 17070
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5816 16720 5868 16726
rect 5816 16662 5868 16668
rect 5446 16552 5502 16561
rect 5446 16487 5502 16496
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 9382 5212 10542
rect 5368 10470 5396 11086
rect 5460 10674 5488 14758
rect 6012 14414 6040 17546
rect 6104 17134 6132 18770
rect 6366 17232 6422 17241
rect 6422 17190 6500 17218
rect 6366 17167 6422 17176
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 16250 6224 16390
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6380 14482 6408 14962
rect 6472 14618 6500 17190
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6380 13802 6408 14418
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6380 13530 6408 13738
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6564 12986 6592 20454
rect 6642 20431 6698 20440
rect 6748 19378 6776 22120
rect 7208 22030 7236 22374
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7104 21956 7156 21962
rect 7104 21898 7156 21904
rect 7116 21842 7144 21898
rect 7300 21842 7328 22374
rect 7484 22234 7512 22578
rect 7576 22438 7604 23666
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7668 23322 7696 23598
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 7838 23080 7894 23089
rect 7838 23015 7894 23024
rect 7656 22772 7708 22778
rect 7656 22714 7708 22720
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7668 22094 7696 22714
rect 7852 22681 7880 23015
rect 7838 22672 7894 22681
rect 7838 22607 7894 22616
rect 7116 21814 7328 21842
rect 7392 22066 7696 22094
rect 7852 22094 7880 22607
rect 7944 22522 7972 25350
rect 8312 24274 8340 26279
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8404 24886 8432 25094
rect 8680 24886 8708 26386
rect 8392 24880 8444 24886
rect 8392 24822 8444 24828
rect 8668 24880 8720 24886
rect 8668 24822 8720 24828
rect 8680 24410 8708 24822
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8116 23316 8168 23322
rect 8116 23258 8168 23264
rect 8128 22710 8156 23258
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8300 23044 8352 23050
rect 8300 22986 8352 22992
rect 8312 22778 8340 22986
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 8496 22545 8524 23054
rect 8482 22536 8538 22545
rect 7944 22494 8248 22522
rect 7852 22066 8156 22094
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 7024 21457 7052 21626
rect 7010 21448 7066 21457
rect 7010 21383 7066 21392
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19514 6960 20198
rect 7024 19938 7052 21383
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 20058 7144 20334
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7024 19910 7144 19938
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 6736 19372 6788 19378
rect 6656 19320 6736 19334
rect 6656 19314 6788 19320
rect 6656 19306 6776 19314
rect 6656 17814 6684 19306
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6840 18290 6868 19178
rect 6932 18834 6960 19450
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7024 18970 7052 19110
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6932 18358 6960 18566
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6656 17066 6684 17750
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6748 16658 6776 18158
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6748 15706 6776 16594
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6840 15162 6868 16118
rect 6932 15502 6960 16594
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6932 15094 6960 15438
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6644 14952 6696 14958
rect 7116 14906 7144 19910
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 7208 18290 7236 19314
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7208 16794 7236 17546
rect 7196 16788 7248 16794
rect 7248 16748 7328 16776
rect 7196 16730 7248 16736
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7208 16250 7236 16458
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 6644 14894 6696 14900
rect 6656 14618 6684 14894
rect 6932 14878 7144 14906
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6840 14006 6868 14486
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6748 13190 6776 13874
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12170 5764 12582
rect 6840 12306 6868 13466
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 6104 11762 6132 12242
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 6104 10606 6132 11698
rect 6196 11354 6224 11698
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 6104 10130 6132 10542
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10266 6408 10406
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 5446 9616 5502 9625
rect 5446 9551 5448 9560
rect 5500 9551 5502 9560
rect 5448 9522 5500 9528
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 9036 5132 9042
rect 4816 8996 5028 9024
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4724 8634 4752 8910
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4908 8514 4936 8842
rect 4632 8492 4936 8514
rect 4632 8486 4712 8492
rect 4764 8486 4936 8492
rect 4712 8434 4764 8440
rect 4264 8350 4660 8378
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7342 4660 8350
rect 4724 7818 4752 8434
rect 5000 8294 5028 8996
rect 5080 8978 5132 8984
rect 5184 8498 5212 9318
rect 5368 9178 5396 9386
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5460 9110 5488 9522
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 8090 5028 8230
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4724 7410 4752 7754
rect 5000 7546 5028 7890
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4724 6662 4752 7346
rect 5184 7342 5212 8434
rect 6104 7954 6132 10066
rect 6380 10010 6408 10066
rect 6288 9994 6408 10010
rect 6276 9988 6408 9994
rect 6328 9982 6408 9988
rect 6276 9930 6328 9936
rect 6564 9722 6592 10610
rect 6932 9926 6960 14878
rect 7300 14822 7328 16748
rect 7392 15162 7420 22066
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7760 21418 7788 21898
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7484 18698 7512 19110
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7576 17882 7604 19314
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7470 17776 7526 17785
rect 8036 17746 8064 19858
rect 7470 17711 7472 17720
rect 7524 17711 7526 17720
rect 8024 17740 8076 17746
rect 7472 17682 7524 17688
rect 8024 17682 8076 17688
rect 8024 17536 8076 17542
rect 8022 17504 8024 17513
rect 8076 17504 8078 17513
rect 8022 17439 8078 17448
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7392 14482 7420 15098
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 13870 7604 14418
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7024 12782 7052 13806
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7012 12776 7064 12782
rect 7064 12736 7144 12764
rect 7012 12718 7064 12724
rect 7116 12084 7144 12736
rect 7208 12238 7236 12922
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7116 12056 7236 12084
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7116 11218 7144 11630
rect 7208 11218 7236 12056
rect 7392 11830 7420 12106
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9722 6960 9862
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 7208 9674 7236 11154
rect 7392 11150 7420 11766
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 9994 7420 11086
rect 7668 10130 7696 14826
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7852 10674 7880 13194
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7932 10056 7984 10062
rect 7852 10004 7932 10010
rect 7852 9998 7984 10004
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7852 9982 7972 9998
rect 7208 9646 7328 9674
rect 7300 9518 7328 9646
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6012 7546 6040 7754
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5092 6934 5120 7278
rect 5276 7002 5304 7346
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 6104 5234 6132 7890
rect 6656 7546 6684 8230
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 7208 6866 7236 8366
rect 7392 7970 7420 9930
rect 7852 9722 7880 9982
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7944 9518 7972 9862
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 8090 7512 8298
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7852 8022 7880 9454
rect 7944 8974 7972 9454
rect 8036 9178 8064 12310
rect 8128 11694 8156 22066
rect 8220 21690 8248 22494
rect 8482 22471 8538 22480
rect 8680 22438 8708 23054
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8300 22160 8352 22166
rect 8298 22128 8300 22137
rect 8352 22128 8354 22137
rect 8298 22063 8354 22072
rect 8404 22030 8432 22374
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 18766 8340 20198
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8312 16590 8340 18702
rect 8496 16726 8524 22374
rect 8576 22160 8628 22166
rect 8576 22102 8628 22108
rect 8588 20602 8616 22102
rect 8864 21622 8892 27474
rect 8956 26246 8984 28494
rect 8944 26240 8996 26246
rect 8944 26182 8996 26188
rect 8944 23044 8996 23050
rect 8944 22986 8996 22992
rect 8956 22710 8984 22986
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 9048 21554 9076 31726
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9416 31278 9444 31622
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9220 31136 9272 31142
rect 9220 31078 9272 31084
rect 9232 30734 9260 31078
rect 9220 30728 9272 30734
rect 9272 30688 9352 30716
rect 9220 30670 9272 30676
rect 9220 30592 9272 30598
rect 9220 30534 9272 30540
rect 9232 30258 9260 30534
rect 9324 30394 9352 30688
rect 9312 30388 9364 30394
rect 9312 30330 9364 30336
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 9128 29776 9180 29782
rect 9128 29718 9180 29724
rect 9140 29578 9168 29718
rect 9128 29572 9180 29578
rect 9128 29514 9180 29520
rect 9140 29238 9168 29514
rect 9128 29232 9180 29238
rect 9128 29174 9180 29180
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9140 28558 9168 28902
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9140 28218 9168 28494
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9128 23044 9180 23050
rect 9128 22986 9180 22992
rect 9140 22030 9168 22986
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9048 20777 9076 21490
rect 9232 21146 9260 30194
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9416 25770 9444 27270
rect 9496 26852 9548 26858
rect 9496 26794 9548 26800
rect 9508 26518 9536 26794
rect 9496 26512 9548 26518
rect 9496 26454 9548 26460
rect 9404 25764 9456 25770
rect 9404 25706 9456 25712
rect 9416 25294 9444 25706
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9416 23254 9444 25230
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9310 22128 9366 22137
rect 9600 22094 9628 31726
rect 9680 31272 9732 31278
rect 9680 31214 9732 31220
rect 9692 30938 9720 31214
rect 9680 30932 9732 30938
rect 9680 30874 9732 30880
rect 9770 30288 9826 30297
rect 9770 30223 9826 30232
rect 9784 30190 9812 30223
rect 9772 30184 9824 30190
rect 9772 30126 9824 30132
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9692 29238 9720 29446
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9680 25424 9732 25430
rect 9680 25366 9732 25372
rect 9692 24954 9720 25366
rect 9680 24948 9732 24954
rect 9680 24890 9732 24896
rect 9784 24750 9812 25434
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9876 22778 9904 33510
rect 9968 32910 9996 34002
rect 10060 33114 10088 37266
rect 10244 35306 10272 38762
rect 10416 38276 10468 38282
rect 10416 38218 10468 38224
rect 10428 38010 10456 38218
rect 10600 38208 10652 38214
rect 10600 38150 10652 38156
rect 10416 38004 10468 38010
rect 10416 37946 10468 37952
rect 10612 37942 10640 38150
rect 10784 38004 10836 38010
rect 10784 37946 10836 37952
rect 10600 37936 10652 37942
rect 10600 37878 10652 37884
rect 10612 36174 10640 37878
rect 10692 36236 10744 36242
rect 10692 36178 10744 36184
rect 10600 36168 10652 36174
rect 10600 36110 10652 36116
rect 10612 35578 10640 36110
rect 10704 35834 10732 36178
rect 10692 35828 10744 35834
rect 10692 35770 10744 35776
rect 10612 35550 10732 35578
rect 10796 35562 10824 37946
rect 11152 37800 11204 37806
rect 11152 37742 11204 37748
rect 11164 37398 11192 37742
rect 11152 37392 11204 37398
rect 11152 37334 11204 37340
rect 10600 35488 10652 35494
rect 10600 35430 10652 35436
rect 10152 35278 10272 35306
rect 10048 33108 10100 33114
rect 10048 33050 10100 33056
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 10048 32904 10100 32910
rect 10048 32846 10100 32852
rect 9968 30258 9996 32846
rect 10060 32502 10088 32846
rect 10048 32496 10100 32502
rect 10048 32438 10100 32444
rect 9956 30252 10008 30258
rect 9956 30194 10008 30200
rect 10152 28994 10180 35278
rect 10612 35154 10640 35430
rect 10600 35148 10652 35154
rect 10600 35090 10652 35096
rect 10704 34950 10732 35550
rect 10784 35556 10836 35562
rect 10784 35498 10836 35504
rect 10232 34944 10284 34950
rect 10232 34886 10284 34892
rect 10692 34944 10744 34950
rect 10692 34886 10744 34892
rect 10244 33998 10272 34886
rect 10704 34610 10732 34886
rect 10692 34604 10744 34610
rect 10692 34546 10744 34552
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 10244 31890 10272 33934
rect 10324 33584 10376 33590
rect 10324 33526 10376 33532
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 10336 29578 10364 33526
rect 10508 33108 10560 33114
rect 10508 33050 10560 33056
rect 10520 30784 10548 33050
rect 10692 32836 10744 32842
rect 10692 32778 10744 32784
rect 10704 32434 10732 32778
rect 10692 32428 10744 32434
rect 10692 32370 10744 32376
rect 10692 32224 10744 32230
rect 10692 32166 10744 32172
rect 10704 31754 10732 32166
rect 10600 31748 10732 31754
rect 10652 31726 10732 31748
rect 10600 31690 10652 31696
rect 10692 30796 10744 30802
rect 10520 30756 10692 30784
rect 10692 30738 10744 30744
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10520 30054 10548 30194
rect 10508 30048 10560 30054
rect 10508 29990 10560 29996
rect 10324 29572 10376 29578
rect 10324 29514 10376 29520
rect 10336 29238 10364 29514
rect 10324 29232 10376 29238
rect 10324 29174 10376 29180
rect 9968 28966 10180 28994
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9310 22063 9312 22072
rect 9364 22063 9366 22072
rect 9508 22066 9628 22094
rect 9312 22034 9364 22040
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9034 20768 9090 20777
rect 9034 20703 9090 20712
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8588 19922 8616 20538
rect 9036 20460 9088 20466
rect 8864 20420 9036 20448
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8666 19816 8722 19825
rect 8666 19751 8722 19760
rect 8680 19378 8708 19751
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 18970 8708 19314
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8312 15094 8340 16526
rect 8496 16250 8524 16662
rect 8588 16250 8616 18226
rect 8680 17746 8708 18906
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8772 18358 8800 18838
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8680 16046 8708 17546
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8312 14414 8340 15030
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 13530 8248 13670
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8220 11354 8248 12786
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8404 10130 8432 12582
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7944 8090 7972 8366
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7840 8016 7892 8022
rect 7392 7942 7512 7970
rect 7840 7958 7892 7964
rect 7484 7818 7512 7942
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 6196 4690 6224 6802
rect 7484 6798 7512 7754
rect 8128 6866 8156 9862
rect 8496 9674 8524 15914
rect 8680 14482 8708 15982
rect 8772 15978 8800 18294
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8772 15162 8800 15438
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8588 10198 8616 13670
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8680 12782 8708 13126
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8772 12238 8800 12854
rect 8864 12442 8892 20420
rect 9036 20402 9088 20408
rect 8944 19304 8996 19310
rect 9140 19292 9168 20878
rect 9324 20584 9352 21490
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 9416 20874 9444 21354
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9508 20602 9536 22066
rect 9968 21842 9996 28966
rect 10232 28960 10284 28966
rect 10232 28902 10284 28908
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10244 28762 10272 28902
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10428 28558 10456 28902
rect 10520 28694 10548 29990
rect 10508 28688 10560 28694
rect 10508 28630 10560 28636
rect 10520 28558 10548 28630
rect 10416 28552 10468 28558
rect 10416 28494 10468 28500
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10324 28484 10376 28490
rect 10324 28426 10376 28432
rect 10140 26988 10192 26994
rect 10140 26930 10192 26936
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10060 25362 10088 25638
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 10048 24948 10100 24954
rect 10048 24890 10100 24896
rect 10060 24614 10088 24890
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 10152 24070 10180 26930
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10244 23746 10272 24686
rect 10336 23866 10364 28426
rect 10600 27600 10652 27606
rect 10600 27542 10652 27548
rect 10612 27062 10640 27542
rect 10704 27538 10732 30738
rect 10796 28642 10824 35498
rect 10876 34944 10928 34950
rect 10876 34886 10928 34892
rect 10888 34746 10916 34886
rect 10876 34740 10928 34746
rect 10876 34682 10928 34688
rect 10876 34604 10928 34610
rect 10876 34546 10928 34552
rect 10888 31754 10916 34546
rect 11060 33312 11112 33318
rect 11060 33254 11112 33260
rect 11072 32502 11100 33254
rect 11060 32496 11112 32502
rect 11060 32438 11112 32444
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 10876 31748 10928 31754
rect 10876 31690 10928 31696
rect 10888 31278 10916 31690
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 11060 31136 11112 31142
rect 11060 31078 11112 31084
rect 11072 30598 11100 31078
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10968 30320 11020 30326
rect 10966 30288 10968 30297
rect 11020 30288 11022 30297
rect 10966 30223 11022 30232
rect 10968 30116 11020 30122
rect 10968 30058 11020 30064
rect 10796 28614 10916 28642
rect 10888 28558 10916 28614
rect 10980 28558 11008 30058
rect 11164 28694 11192 31962
rect 11256 31754 11284 38830
rect 11624 38010 11652 38898
rect 11992 38214 12020 38898
rect 12348 38752 12400 38758
rect 12348 38694 12400 38700
rect 12440 38752 12492 38758
rect 12440 38694 12492 38700
rect 12360 38418 12388 38694
rect 12452 38554 12480 38694
rect 12440 38548 12492 38554
rect 12440 38490 12492 38496
rect 12348 38412 12400 38418
rect 12348 38354 12400 38360
rect 11888 38208 11940 38214
rect 11888 38150 11940 38156
rect 11980 38208 12032 38214
rect 11980 38150 12032 38156
rect 11612 38004 11664 38010
rect 11612 37946 11664 37952
rect 11702 37904 11758 37913
rect 11702 37839 11704 37848
rect 11756 37839 11758 37848
rect 11704 37810 11756 37816
rect 11900 37738 11928 38150
rect 12728 38010 12756 38898
rect 13004 38729 13032 38898
rect 16040 38826 16068 38966
rect 19996 38962 20024 40762
rect 21928 39098 21956 40762
rect 26436 39098 26464 40762
rect 21916 39092 21968 39098
rect 21916 39034 21968 39040
rect 26424 39092 26476 39098
rect 26424 39034 26476 39040
rect 30944 39030 30972 40762
rect 32876 39098 32904 40762
rect 35820 39794 35848 40854
rect 37370 40762 37426 41562
rect 39302 40762 39358 41562
rect 35820 39766 35940 39794
rect 32864 39092 32916 39098
rect 32864 39034 32916 39040
rect 35912 39030 35940 39766
rect 24400 39024 24452 39030
rect 24400 38966 24452 38972
rect 30932 39024 30984 39030
rect 30932 38966 30984 38972
rect 35900 39024 35952 39030
rect 35900 38966 35952 38972
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 16028 38820 16080 38826
rect 16028 38762 16080 38768
rect 22112 38729 22140 38898
rect 12990 38720 13046 38729
rect 12990 38655 13046 38664
rect 22098 38720 22154 38729
rect 22098 38655 22154 38664
rect 24412 38554 24440 38966
rect 37384 38962 37412 40762
rect 24768 38956 24820 38962
rect 24768 38898 24820 38904
rect 25044 38956 25096 38962
rect 25044 38898 25096 38904
rect 27068 38956 27120 38962
rect 27068 38898 27120 38904
rect 33048 38956 33100 38962
rect 33048 38898 33100 38904
rect 35624 38956 35676 38962
rect 35624 38898 35676 38904
rect 37372 38956 37424 38962
rect 37372 38898 37424 38904
rect 17500 38548 17552 38554
rect 17500 38490 17552 38496
rect 22652 38548 22704 38554
rect 22652 38490 22704 38496
rect 24400 38548 24452 38554
rect 24400 38490 24452 38496
rect 14464 38412 14516 38418
rect 14464 38354 14516 38360
rect 14004 38276 14056 38282
rect 14004 38218 14056 38224
rect 13728 38208 13780 38214
rect 13728 38150 13780 38156
rect 13740 38010 13768 38150
rect 12716 38004 12768 38010
rect 12716 37946 12768 37952
rect 13728 38004 13780 38010
rect 13728 37946 13780 37952
rect 13084 37936 13136 37942
rect 13084 37878 13136 37884
rect 11888 37732 11940 37738
rect 11888 37674 11940 37680
rect 12348 37732 12400 37738
rect 12348 37674 12400 37680
rect 11796 37120 11848 37126
rect 11796 37062 11848 37068
rect 11808 36650 11836 37062
rect 11796 36644 11848 36650
rect 11796 36586 11848 36592
rect 11808 35698 11836 36586
rect 12360 36174 12388 37674
rect 12348 36168 12400 36174
rect 12348 36110 12400 36116
rect 12624 36168 12676 36174
rect 12624 36110 12676 36116
rect 12808 36168 12860 36174
rect 12808 36110 12860 36116
rect 12440 36100 12492 36106
rect 12440 36042 12492 36048
rect 11980 35760 12032 35766
rect 11980 35702 12032 35708
rect 11796 35692 11848 35698
rect 11796 35634 11848 35640
rect 11520 32428 11572 32434
rect 11520 32370 11572 32376
rect 11256 31726 11376 31754
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11256 30666 11284 31078
rect 11244 30660 11296 30666
rect 11244 30602 11296 30608
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 10692 27532 10744 27538
rect 10692 27474 10744 27480
rect 10600 27056 10652 27062
rect 10600 26998 10652 27004
rect 10612 26926 10640 26998
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 26586 10640 26726
rect 10600 26580 10652 26586
rect 10600 26522 10652 26528
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10428 25498 10456 25842
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10244 23718 10364 23746
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 23186 10272 23462
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10336 21962 10364 23718
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10796 22574 10824 23666
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10888 22094 10916 28494
rect 10980 27690 11008 28494
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 11072 27946 11100 28358
rect 11348 28234 11376 31726
rect 11532 31482 11560 32370
rect 11702 32056 11758 32065
rect 11702 31991 11704 32000
rect 11756 31991 11758 32000
rect 11704 31962 11756 31968
rect 11520 31476 11572 31482
rect 11520 31418 11572 31424
rect 11520 31136 11572 31142
rect 11520 31078 11572 31084
rect 11532 29102 11560 31078
rect 11808 29322 11836 35634
rect 11992 35290 12020 35702
rect 12256 35624 12308 35630
rect 12256 35566 12308 35572
rect 11888 35284 11940 35290
rect 11888 35226 11940 35232
rect 11980 35284 12032 35290
rect 11980 35226 12032 35232
rect 12072 35284 12124 35290
rect 12072 35226 12124 35232
rect 11900 34610 11928 35226
rect 12084 35034 12112 35226
rect 11992 35006 12112 35034
rect 11992 34950 12020 35006
rect 11980 34944 12032 34950
rect 11980 34886 12032 34892
rect 11888 34604 11940 34610
rect 11888 34546 11940 34552
rect 11980 34196 12032 34202
rect 11980 34138 12032 34144
rect 11992 32881 12020 34138
rect 12268 32994 12296 35566
rect 12452 34610 12480 36042
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 12348 34128 12400 34134
rect 12348 34070 12400 34076
rect 12360 33833 12388 34070
rect 12346 33824 12402 33833
rect 12346 33759 12402 33768
rect 12176 32966 12296 32994
rect 11978 32872 12034 32881
rect 11978 32807 12034 32816
rect 11992 32434 12020 32807
rect 11980 32428 12032 32434
rect 11980 32370 12032 32376
rect 11992 30258 12020 32370
rect 12072 31680 12124 31686
rect 12072 31622 12124 31628
rect 12084 31278 12112 31622
rect 12176 31278 12204 32966
rect 12348 32564 12400 32570
rect 12348 32506 12400 32512
rect 12360 32434 12388 32506
rect 12348 32428 12400 32434
rect 12348 32370 12400 32376
rect 12452 32366 12480 34546
rect 12532 34400 12584 34406
rect 12532 34342 12584 34348
rect 12544 33998 12572 34342
rect 12636 33998 12664 36110
rect 12820 35698 12848 36110
rect 12992 36032 13044 36038
rect 12990 36000 12992 36009
rect 13044 36000 13046 36009
rect 12990 35935 13046 35944
rect 13096 35714 13124 37878
rect 13268 37392 13320 37398
rect 13268 37334 13320 37340
rect 13004 35698 13124 35714
rect 13280 35698 13308 37334
rect 13636 36168 13688 36174
rect 13636 36110 13688 36116
rect 13648 35834 13676 36110
rect 13636 35828 13688 35834
rect 13636 35770 13688 35776
rect 12808 35692 12860 35698
rect 12808 35634 12860 35640
rect 12992 35692 13124 35698
rect 13044 35686 13124 35692
rect 13176 35692 13228 35698
rect 12992 35634 13044 35640
rect 13176 35634 13228 35640
rect 13268 35692 13320 35698
rect 13268 35634 13320 35640
rect 13360 35692 13412 35698
rect 13360 35634 13412 35640
rect 12716 35488 12768 35494
rect 12716 35430 12768 35436
rect 12728 34474 12756 35430
rect 12716 34468 12768 34474
rect 12716 34410 12768 34416
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12624 33992 12676 33998
rect 12624 33934 12676 33940
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 12544 33590 12572 33798
rect 12532 33584 12584 33590
rect 12532 33526 12584 33532
rect 12532 33380 12584 33386
rect 12532 33322 12584 33328
rect 12440 32360 12492 32366
rect 12440 32302 12492 32308
rect 12072 31272 12124 31278
rect 12072 31214 12124 31220
rect 12164 31272 12216 31278
rect 12164 31214 12216 31220
rect 12084 30938 12112 31214
rect 12072 30932 12124 30938
rect 12072 30874 12124 30880
rect 11980 30252 12032 30258
rect 11980 30194 12032 30200
rect 11992 29510 12020 30194
rect 12070 29608 12126 29617
rect 12070 29543 12126 29552
rect 11980 29504 12032 29510
rect 11980 29446 12032 29452
rect 11808 29294 12020 29322
rect 11520 29096 11572 29102
rect 11520 29038 11572 29044
rect 11888 29096 11940 29102
rect 11888 29038 11940 29044
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11164 28206 11376 28234
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 10980 27662 11100 27690
rect 10968 27328 11020 27334
rect 10968 27270 11020 27276
rect 10980 26994 11008 27270
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10968 26784 11020 26790
rect 10968 26726 11020 26732
rect 10980 26314 11008 26726
rect 10968 26308 11020 26314
rect 10968 26250 11020 26256
rect 10980 25922 11008 26250
rect 11072 26042 11100 27662
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 10980 25894 11100 25922
rect 11072 25294 11100 25894
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10796 22066 10916 22094
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 9784 21814 10088 21842
rect 9784 21554 9812 21814
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9876 21434 9904 21490
rect 9784 21406 9904 21434
rect 9784 21350 9812 21406
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9784 20942 9812 21286
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9496 20596 9548 20602
rect 9324 20556 9444 20584
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9324 20058 9352 20402
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9324 19514 9352 19654
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9416 19394 9444 20556
rect 9496 20538 9548 20544
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 8996 19264 9168 19292
rect 9324 19366 9444 19394
rect 9600 19378 9628 19654
rect 9588 19372 9640 19378
rect 8944 19246 8996 19252
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11898 8708 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8772 11558 8800 12174
rect 8864 11762 8892 12378
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8956 11642 8984 19246
rect 9324 19174 9352 19366
rect 9588 19314 9640 19320
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9140 18426 9168 18702
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 9048 16590 9076 18226
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9232 16998 9260 17138
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 16114 9168 16390
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9034 16008 9090 16017
rect 9034 15943 9036 15952
rect 9088 15943 9090 15952
rect 9128 15972 9180 15978
rect 9036 15914 9088 15920
rect 9128 15914 9180 15920
rect 9034 15192 9090 15201
rect 9034 15127 9090 15136
rect 9048 13870 9076 15127
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9048 12714 9076 13806
rect 9140 13258 9168 15914
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9232 12986 9260 16594
rect 9324 16114 9352 19110
rect 9600 18290 9628 19314
rect 9692 18306 9720 20742
rect 9784 20534 9812 20878
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9784 20262 9812 20470
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9876 19786 9904 20810
rect 9968 20806 9996 21490
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9968 19009 9996 20402
rect 9954 19000 10010 19009
rect 9954 18935 10010 18944
rect 9862 18320 9918 18329
rect 9588 18284 9640 18290
rect 9692 18278 9862 18306
rect 9862 18255 9918 18264
rect 9588 18226 9640 18232
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9600 17882 9628 18090
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9692 17746 9720 18090
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9588 17536 9640 17542
rect 9586 17504 9588 17513
rect 9640 17504 9642 17513
rect 9586 17439 9642 17448
rect 9692 17202 9720 17682
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9784 17270 9812 17546
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9600 16612 9812 16640
rect 9496 16584 9548 16590
rect 9600 16572 9628 16612
rect 9548 16544 9628 16572
rect 9496 16526 9548 16532
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9678 16416 9734 16425
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9324 15094 9352 15506
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9324 14006 9352 15030
rect 9416 15026 9444 16390
rect 9600 15706 9628 16390
rect 9678 16351 9734 16360
rect 9692 16114 9720 16351
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9312 13184 9364 13190
rect 9416 13172 9444 14962
rect 9784 14006 9812 16612
rect 9876 14890 9904 18255
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9968 17066 9996 17614
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 10060 16658 10088 21814
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10336 21078 10364 21422
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 10704 20942 10732 21490
rect 10796 21146 10824 22066
rect 10876 21956 10928 21962
rect 10876 21898 10928 21904
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10140 20868 10192 20874
rect 10140 20810 10192 20816
rect 10152 18698 10180 20810
rect 10336 20777 10364 20878
rect 10428 20806 10456 20878
rect 10416 20800 10468 20806
rect 10322 20768 10378 20777
rect 10416 20742 10468 20748
rect 10322 20703 10378 20712
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10152 17882 10180 18226
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9968 15162 9996 15302
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 14006 10180 14214
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9508 13258 9536 13670
rect 9600 13530 9628 13670
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9364 13144 9444 13172
rect 9312 13126 9364 13132
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11830 9260 12174
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 8864 11614 8984 11642
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8680 11150 8708 11494
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8680 10266 8708 10950
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8576 10192 8628 10198
rect 8628 10140 8708 10146
rect 8576 10134 8708 10140
rect 8588 10118 8708 10134
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8208 9648 8260 9654
rect 8206 9616 8208 9625
rect 8312 9646 8524 9674
rect 8588 9654 8616 9862
rect 8260 9616 8262 9625
rect 8312 9586 8340 9646
rect 8206 9551 8262 9560
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9042 8248 9318
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8496 8906 8524 9646
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8680 9586 8708 10118
rect 8772 10062 8800 10406
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8864 9994 8892 11614
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8956 9625 8984 11494
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9048 10130 9076 11222
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9140 10266 9168 10474
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9324 10146 9352 12718
rect 9416 12374 9444 13144
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12782 9628 13126
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9876 12434 9904 13330
rect 9784 12406 9904 12434
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9784 12238 9812 12406
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9416 11558 9444 11834
rect 9508 11626 9536 12038
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 10266 9444 11494
rect 9600 11150 9628 11698
rect 9784 11694 9812 12174
rect 9968 11830 9996 13942
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10060 13394 10088 13874
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 10060 11150 10088 13330
rect 10244 12594 10272 20470
rect 10428 20466 10456 20742
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10336 13530 10364 20402
rect 10428 20262 10456 20402
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10414 19136 10470 19145
rect 10414 19071 10470 19080
rect 10428 18902 10456 19071
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10428 18222 10456 18566
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10414 18048 10470 18057
rect 10414 17983 10470 17992
rect 10428 17542 10456 17983
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10428 12850 10456 13330
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10416 12640 10468 12646
rect 10244 12566 10364 12594
rect 10416 12582 10468 12588
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9140 10118 9352 10146
rect 9140 10062 9168 10118
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8942 9616 8998 9625
rect 8668 9580 8720 9586
rect 8852 9580 8904 9586
rect 8720 9540 8852 9568
rect 8668 9522 8720 9528
rect 8942 9551 8998 9560
rect 8852 9522 8904 9528
rect 9048 9466 9076 9930
rect 8956 9438 9076 9466
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6472 6458 6500 6666
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5370 7328 5510
rect 7484 5370 7512 6734
rect 7944 5914 7972 6734
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6458 8064 6598
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8128 6186 8156 6802
rect 8220 6798 8248 8842
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 8566 8340 8774
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8496 8498 8524 8842
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8588 6866 8616 8910
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8634 8800 8774
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6458 8248 6734
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8312 6458 8340 6666
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6458 8432 6598
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8220 5710 8248 6258
rect 8392 6248 8444 6254
rect 8444 6196 8524 6202
rect 8392 6190 8524 6196
rect 8300 6180 8352 6186
rect 8404 6174 8524 6190
rect 8588 6186 8616 6802
rect 8300 6122 8352 6128
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5370 8248 5646
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 7484 4554 7512 5306
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4826 8248 4966
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8312 4622 8340 6122
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5710 8432 6054
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8496 5234 8524 6174
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8588 5914 8616 6122
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 8312 4146 8340 4558
rect 8588 4282 8616 5170
rect 8680 4826 8708 5170
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 3988 2746 4108 2774
rect 4080 2446 4108 2746
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8220 2446 8248 2790
rect 8956 2774 8984 9438
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9232 7546 9260 7754
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9324 7274 9352 9998
rect 9508 8838 9536 10202
rect 9600 10062 9628 11086
rect 10060 10810 10088 11086
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10138 10704 10194 10713
rect 9772 10668 9824 10674
rect 10138 10639 10194 10648
rect 9772 10610 9824 10616
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9416 7410 9444 8026
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9508 7342 9536 7686
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9048 5710 9076 6394
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5846 9260 6190
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9048 4758 9076 5306
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 9232 4554 9260 5782
rect 9324 5098 9352 6258
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5914 9444 6054
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 5234 9444 5646
rect 9508 5234 9536 7278
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9324 4622 9352 5034
rect 9508 4690 9536 5170
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 8680 2746 8984 2774
rect 8680 2650 8708 2746
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 9600 2446 9628 8774
rect 9784 5710 9812 10610
rect 10152 10606 10180 10639
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10152 10470 10180 10542
rect 10140 10464 10192 10470
rect 10336 10441 10364 12566
rect 10428 12322 10456 12582
rect 10520 12434 10548 20538
rect 10704 20466 10732 20878
rect 10888 20602 10916 21898
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10600 18760 10652 18766
rect 10598 18728 10600 18737
rect 10652 18728 10654 18737
rect 10598 18663 10654 18672
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10612 18426 10640 18566
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10704 18290 10732 18906
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10600 18216 10652 18222
rect 10598 18184 10600 18193
rect 10652 18184 10654 18193
rect 10598 18119 10654 18128
rect 10704 17882 10732 18226
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10796 17746 10824 19246
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10796 17338 10824 17682
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10888 12986 10916 19382
rect 10980 19378 11008 22646
rect 11164 20942 11192 28206
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11348 27674 11376 28018
rect 11336 27668 11388 27674
rect 11336 27610 11388 27616
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11256 20330 11284 24006
rect 11348 23254 11376 25230
rect 11440 24274 11468 28494
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11716 28150 11744 28358
rect 11704 28144 11756 28150
rect 11704 28086 11756 28092
rect 11520 27872 11572 27878
rect 11572 27820 11652 27826
rect 11520 27814 11652 27820
rect 11532 27798 11652 27814
rect 11624 27690 11652 27798
rect 11624 27674 11836 27690
rect 11624 27668 11848 27674
rect 11624 27662 11796 27668
rect 11796 27610 11848 27616
rect 11704 27600 11756 27606
rect 11704 27542 11756 27548
rect 11520 27328 11572 27334
rect 11520 27270 11572 27276
rect 11532 27130 11560 27270
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11716 24818 11744 27542
rect 11796 27328 11848 27334
rect 11796 27270 11848 27276
rect 11808 26926 11836 27270
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11900 25906 11928 29038
rect 11992 27146 12020 29294
rect 12084 29102 12112 29543
rect 12072 29096 12124 29102
rect 12072 29038 12124 29044
rect 12176 28994 12204 31214
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12256 29232 12308 29238
rect 12256 29174 12308 29180
rect 12084 28966 12204 28994
rect 12084 27606 12112 28966
rect 12268 28234 12296 29174
rect 12360 29170 12388 29582
rect 12348 29164 12400 29170
rect 12348 29106 12400 29112
rect 12452 28762 12480 30262
rect 12544 29850 12572 33322
rect 12728 32774 12756 34410
rect 12820 34202 12848 35634
rect 13188 34610 13216 35634
rect 12900 34604 12952 34610
rect 12900 34546 12952 34552
rect 13176 34604 13228 34610
rect 13176 34546 13228 34552
rect 12808 34196 12860 34202
rect 12808 34138 12860 34144
rect 12716 32768 12768 32774
rect 12716 32710 12768 32716
rect 12808 32768 12860 32774
rect 12808 32710 12860 32716
rect 12624 32292 12676 32298
rect 12624 32234 12676 32240
rect 12636 30734 12664 32234
rect 12716 32020 12768 32026
rect 12716 31962 12768 31968
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12440 28756 12492 28762
rect 12440 28698 12492 28704
rect 12176 28206 12296 28234
rect 12072 27600 12124 27606
rect 12072 27542 12124 27548
rect 11992 27118 12112 27146
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 11992 26586 12020 26998
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11900 25786 11928 25842
rect 12084 25786 12112 27118
rect 12176 26586 12204 28206
rect 12256 28144 12308 28150
rect 12256 28086 12308 28092
rect 12268 26790 12296 28086
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12164 26580 12216 26586
rect 12164 26522 12216 26528
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 11808 25758 11928 25786
rect 11992 25758 12112 25786
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11440 23730 11468 24210
rect 11612 23792 11664 23798
rect 11612 23734 11664 23740
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11440 22506 11468 23666
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 11532 22778 11560 23598
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11428 22500 11480 22506
rect 11428 22442 11480 22448
rect 11440 22094 11468 22442
rect 11520 22094 11572 22098
rect 11440 22092 11572 22094
rect 11440 22066 11520 22092
rect 11520 22034 11572 22040
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11164 19514 11192 19722
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 11072 18986 11100 19382
rect 11348 19334 11376 21830
rect 11624 20369 11652 23734
rect 11808 20466 11836 25758
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11900 22778 11928 22986
rect 11992 22778 12020 25758
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 12084 25265 12112 25638
rect 12176 25362 12204 25978
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 12070 25256 12126 25265
rect 12070 25191 12126 25200
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 12084 24410 12112 25094
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11992 22234 12020 22510
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 11886 21312 11942 21321
rect 11886 21247 11942 21256
rect 11900 20602 11928 21247
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11610 20360 11666 20369
rect 11610 20295 11666 20304
rect 11808 19990 11836 20402
rect 11612 19984 11664 19990
rect 11612 19926 11664 19932
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 10980 18958 11100 18986
rect 11256 19306 11376 19334
rect 10980 18902 11008 18958
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10968 18760 11020 18766
rect 10966 18728 10968 18737
rect 11020 18728 11022 18737
rect 10966 18663 11022 18672
rect 10980 18290 11008 18663
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10980 17542 11008 18226
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 17202 11008 17478
rect 11072 17338 11100 18090
rect 11256 17921 11284 19306
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11348 18193 11376 18226
rect 11334 18184 11390 18193
rect 11334 18119 11390 18128
rect 11242 17912 11298 17921
rect 11242 17847 11298 17856
rect 11336 17876 11388 17882
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11164 17338 11192 17682
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11256 17202 11284 17847
rect 11336 17818 11388 17824
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11244 17196 11296 17202
rect 11348 17184 11376 17818
rect 11440 17338 11468 17818
rect 11532 17678 11560 19246
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11428 17196 11480 17202
rect 11348 17156 11428 17184
rect 11244 17138 11296 17144
rect 11428 17138 11480 17144
rect 11440 16998 11468 17138
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 14414 11100 15438
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 11348 15162 11376 15370
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10520 12406 10640 12434
rect 10428 12294 10548 12322
rect 10520 12170 10548 12294
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10416 11552 10468 11558
rect 10612 11540 10640 12406
rect 10468 11512 10640 11540
rect 10416 11494 10468 11500
rect 10428 11150 10456 11494
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10140 10406 10192 10412
rect 10322 10432 10378 10441
rect 10152 9602 10180 10406
rect 10322 10367 10378 10376
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10244 9722 10272 9998
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10152 9586 10272 9602
rect 10152 9580 10284 9586
rect 10152 9574 10232 9580
rect 10232 9522 10284 9528
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8634 10088 8910
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10152 7478 10180 9454
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 5302 10088 5510
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 10244 2514 10272 9522
rect 10336 9042 10364 10367
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10428 6662 10456 11086
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 9586 10640 10406
rect 10888 9654 10916 12922
rect 11072 12306 11100 14350
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11164 13530 11192 14010
rect 11348 13870 11376 14894
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11348 12850 11376 13806
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11624 12442 11652 19926
rect 11900 19922 11928 20538
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11886 19272 11942 19281
rect 11886 19207 11888 19216
rect 11940 19207 11942 19216
rect 11888 19178 11940 19184
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11808 18290 11836 18702
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11702 18048 11758 18057
rect 11702 17983 11758 17992
rect 11716 17762 11744 17983
rect 11808 17882 11836 18226
rect 11900 18086 11928 18702
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18222 12020 18566
rect 12084 18222 12112 24006
rect 12176 22574 12204 25298
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12268 24070 12296 24890
rect 12360 24614 12388 27474
rect 12636 27402 12664 30670
rect 12728 29730 12756 31962
rect 12820 31822 12848 32710
rect 12912 32434 12940 34546
rect 13084 33856 13136 33862
rect 13084 33798 13136 33804
rect 13096 32910 13124 33798
rect 13084 32904 13136 32910
rect 13084 32846 13136 32852
rect 12900 32428 12952 32434
rect 12952 32388 13032 32416
rect 12900 32370 12952 32376
rect 12900 32224 12952 32230
rect 12900 32166 12952 32172
rect 12912 31822 12940 32166
rect 12808 31816 12860 31822
rect 12808 31758 12860 31764
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12900 30320 12952 30326
rect 13004 30308 13032 32388
rect 13096 30734 13124 32846
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13188 32065 13216 32166
rect 13174 32056 13230 32065
rect 13174 31991 13230 32000
rect 13280 31142 13308 35634
rect 13372 35494 13400 35634
rect 13360 35488 13412 35494
rect 13360 35430 13412 35436
rect 13452 32836 13504 32842
rect 13452 32778 13504 32784
rect 13268 31136 13320 31142
rect 13268 31078 13320 31084
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 12952 30280 13032 30308
rect 12900 30262 12952 30268
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12912 29850 12940 29990
rect 12900 29844 12952 29850
rect 12900 29786 12952 29792
rect 12728 29702 13032 29730
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12912 28558 12940 29446
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 12636 25770 12664 27338
rect 12806 27160 12862 27169
rect 12806 27095 12862 27104
rect 12820 27062 12848 27095
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12912 26994 12940 28494
rect 12900 26988 12952 26994
rect 12900 26930 12952 26936
rect 12912 26586 12940 26930
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 12544 24410 12572 24754
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12728 24342 12756 25094
rect 12716 24336 12768 24342
rect 12714 24304 12716 24313
rect 12768 24304 12770 24313
rect 12714 24239 12770 24248
rect 12912 24206 12940 25298
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12728 23866 12756 24142
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12912 23118 12940 24142
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12176 22094 12204 22510
rect 12176 22066 12388 22094
rect 12256 22024 12308 22030
rect 12254 21992 12256 22001
rect 12308 21992 12310 22001
rect 12254 21927 12310 21936
rect 12256 20936 12308 20942
rect 12256 20878 12308 20884
rect 12164 20868 12216 20874
rect 12164 20810 12216 20816
rect 12176 20466 12204 20810
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12162 20360 12218 20369
rect 12162 20295 12218 20304
rect 12176 18970 12204 20295
rect 12268 19922 12296 20878
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11716 17734 11836 17762
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11716 17542 11744 17614
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11716 17202 11744 17478
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11808 15162 11836 17734
rect 11900 17184 11928 18022
rect 12084 17649 12112 18158
rect 12070 17640 12126 17649
rect 12070 17575 12126 17584
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17338 12204 17478
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12360 17270 12388 22066
rect 12452 21146 12480 22578
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 18737 12480 20198
rect 12636 19802 12664 21966
rect 12912 21622 12940 21966
rect 12900 21616 12952 21622
rect 12900 21558 12952 21564
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12728 20466 12756 20878
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12636 19774 12756 19802
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 18970 12572 19246
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12438 18728 12494 18737
rect 12438 18663 12494 18672
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12452 17202 12480 18663
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 18290 12572 18566
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12636 18057 12664 19654
rect 12728 19242 12756 19774
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 19145 12756 19178
rect 12714 19136 12770 19145
rect 12714 19071 12770 19080
rect 12820 18698 12848 19722
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 18426 12756 18566
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12622 18048 12678 18057
rect 12622 17983 12678 17992
rect 12820 17513 12848 18634
rect 12806 17504 12862 17513
rect 12806 17439 12862 17448
rect 11980 17196 12032 17202
rect 11900 17156 11980 17184
rect 11980 17138 12032 17144
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 11992 15366 12020 17138
rect 12176 16182 12204 17138
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11796 15156 11848 15162
rect 11848 15116 11928 15144
rect 11796 15098 11848 15104
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 14074 11744 14214
rect 11808 14074 11836 14282
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11900 13938 11928 15116
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 12084 13734 12112 14894
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11992 12306 12020 12922
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10130 11100 11086
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10980 7410 11008 9862
rect 11164 9518 11192 11698
rect 11532 11150 11560 12038
rect 12084 11762 12112 13670
rect 12268 12986 12296 17002
rect 12912 16946 12940 21422
rect 13004 19378 13032 29702
rect 13096 28966 13124 30670
rect 13464 30258 13492 32778
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13636 30592 13688 30598
rect 13636 30534 13688 30540
rect 13452 30252 13504 30258
rect 13504 30212 13584 30240
rect 13452 30194 13504 30200
rect 13360 29504 13412 29510
rect 13412 29464 13492 29492
rect 13360 29446 13412 29452
rect 13358 29064 13414 29073
rect 13358 28999 13360 29008
rect 13412 28999 13414 29008
rect 13360 28970 13412 28976
rect 13084 28960 13136 28966
rect 13084 28902 13136 28908
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 13096 27062 13124 28698
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 13280 27606 13308 27950
rect 13268 27600 13320 27606
rect 13268 27542 13320 27548
rect 13188 27084 13400 27112
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 13084 26240 13136 26246
rect 13084 26182 13136 26188
rect 13096 25158 13124 26182
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13096 23644 13124 25094
rect 13188 24857 13216 27084
rect 13372 26994 13400 27084
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 13280 26450 13308 26930
rect 13268 26444 13320 26450
rect 13268 26386 13320 26392
rect 13280 25498 13308 26386
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13372 25362 13400 26182
rect 13360 25356 13412 25362
rect 13360 25298 13412 25304
rect 13174 24848 13230 24857
rect 13174 24783 13230 24792
rect 13372 24682 13400 25298
rect 13360 24676 13412 24682
rect 13360 24618 13412 24624
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13280 23798 13308 24550
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13372 23905 13400 24142
rect 13358 23896 13414 23905
rect 13358 23831 13360 23840
rect 13412 23831 13414 23840
rect 13360 23802 13412 23808
rect 13268 23792 13320 23798
rect 13268 23734 13320 23740
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13096 23616 13308 23644
rect 13176 22500 13228 22506
rect 13176 22442 13228 22448
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13188 19258 13216 22442
rect 13280 19666 13308 23616
rect 13372 23526 13400 23666
rect 13464 23644 13492 29464
rect 13556 26994 13584 30212
rect 13648 29646 13676 30534
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 13636 28960 13688 28966
rect 13636 28902 13688 28908
rect 13648 27470 13676 28902
rect 13636 27464 13688 27470
rect 13636 27406 13688 27412
rect 13636 27328 13688 27334
rect 13636 27270 13688 27276
rect 13648 26994 13676 27270
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 13636 26988 13688 26994
rect 13636 26930 13688 26936
rect 13740 25974 13768 31282
rect 14016 30122 14044 38218
rect 14476 38010 14504 38354
rect 16212 38208 16264 38214
rect 16212 38150 16264 38156
rect 14464 38004 14516 38010
rect 14464 37946 14516 37952
rect 14556 38004 14608 38010
rect 14556 37946 14608 37952
rect 14280 37868 14332 37874
rect 14280 37810 14332 37816
rect 14372 37868 14424 37874
rect 14372 37810 14424 37816
rect 14292 37262 14320 37810
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 14188 35692 14240 35698
rect 14188 35634 14240 35640
rect 14096 33584 14148 33590
rect 14096 33526 14148 33532
rect 14108 33425 14136 33526
rect 14094 33416 14150 33425
rect 14094 33351 14150 33360
rect 14004 30116 14056 30122
rect 14004 30058 14056 30064
rect 13910 29880 13966 29889
rect 13910 29815 13966 29824
rect 13924 29646 13952 29815
rect 13912 29640 13964 29646
rect 13912 29582 13964 29588
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13832 26790 13860 27474
rect 13924 27062 13952 29582
rect 14016 29238 14044 30058
rect 14200 29617 14228 35634
rect 14384 35086 14412 37810
rect 14476 37369 14504 37946
rect 14462 37360 14518 37369
rect 14462 37295 14518 37304
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14280 34128 14332 34134
rect 14280 34070 14332 34076
rect 14292 31754 14320 34070
rect 14384 33522 14412 35022
rect 14464 34944 14516 34950
rect 14568 34932 14596 37946
rect 14832 37868 14884 37874
rect 14832 37810 14884 37816
rect 15752 37868 15804 37874
rect 15752 37810 15804 37816
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 14740 36100 14792 36106
rect 14740 36042 14792 36048
rect 14516 34904 14596 34932
rect 14648 34944 14700 34950
rect 14464 34886 14516 34892
rect 14648 34886 14700 34892
rect 14476 33590 14504 34886
rect 14660 34202 14688 34886
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 14752 33998 14780 36042
rect 14844 35086 14872 37810
rect 15200 37664 15252 37670
rect 15200 37606 15252 37612
rect 15108 37188 15160 37194
rect 15108 37130 15160 37136
rect 15120 36825 15148 37130
rect 15106 36816 15162 36825
rect 15106 36751 15162 36760
rect 14832 35080 14884 35086
rect 14832 35022 14884 35028
rect 15120 34610 15148 36751
rect 15212 36174 15240 37606
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15304 36174 15332 36518
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 15292 36168 15344 36174
rect 15292 36110 15344 36116
rect 15568 36168 15620 36174
rect 15568 36110 15620 36116
rect 15580 35834 15608 36110
rect 15568 35828 15620 35834
rect 15568 35770 15620 35776
rect 15384 34944 15436 34950
rect 15384 34886 15436 34892
rect 15108 34604 15160 34610
rect 15108 34546 15160 34552
rect 14740 33992 14792 33998
rect 14924 33992 14976 33998
rect 14792 33952 14872 33980
rect 14740 33934 14792 33940
rect 14464 33584 14516 33590
rect 14464 33526 14516 33532
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14648 33516 14700 33522
rect 14648 33458 14700 33464
rect 14280 31748 14332 31754
rect 14280 31690 14332 31696
rect 14292 31482 14320 31690
rect 14384 31686 14412 33458
rect 14464 32836 14516 32842
rect 14464 32778 14516 32784
rect 14476 32366 14504 32778
rect 14464 32360 14516 32366
rect 14464 32302 14516 32308
rect 14464 31748 14516 31754
rect 14568 31736 14596 33458
rect 14516 31708 14596 31736
rect 14464 31690 14516 31696
rect 14372 31680 14424 31686
rect 14372 31622 14424 31628
rect 14280 31476 14332 31482
rect 14280 31418 14332 31424
rect 14384 30258 14412 31622
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14186 29608 14242 29617
rect 14186 29543 14242 29552
rect 14004 29232 14056 29238
rect 14004 29174 14056 29180
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14200 28626 14228 29106
rect 14188 28620 14240 28626
rect 14188 28562 14240 28568
rect 14384 28082 14412 30194
rect 14476 28234 14504 31690
rect 14660 31686 14688 33458
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 14648 31680 14700 31686
rect 14648 31622 14700 31628
rect 14556 30592 14608 30598
rect 14556 30534 14608 30540
rect 14568 29646 14596 30534
rect 14660 30104 14688 31622
rect 14752 30326 14780 31826
rect 14844 31754 14872 33952
rect 14924 33934 14976 33940
rect 14936 33658 14964 33934
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 15200 32428 15252 32434
rect 15200 32370 15252 32376
rect 14844 31726 15148 31754
rect 14924 31680 14976 31686
rect 14924 31622 14976 31628
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14844 30326 14872 30806
rect 14936 30802 14964 31622
rect 14924 30796 14976 30802
rect 14924 30738 14976 30744
rect 15120 30734 15148 31726
rect 15212 31521 15240 32370
rect 15198 31512 15254 31521
rect 15198 31447 15254 31456
rect 15292 31340 15344 31346
rect 15292 31282 15344 31288
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 14924 30592 14976 30598
rect 14924 30534 14976 30540
rect 14936 30394 14964 30534
rect 15028 30394 15056 30670
rect 14924 30388 14976 30394
rect 14924 30330 14976 30336
rect 15016 30388 15068 30394
rect 15016 30330 15068 30336
rect 14740 30320 14792 30326
rect 14740 30262 14792 30268
rect 14832 30320 14884 30326
rect 14832 30262 14884 30268
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15028 30161 15056 30194
rect 15014 30152 15070 30161
rect 14740 30116 14792 30122
rect 14660 30076 14740 30104
rect 15014 30087 15070 30096
rect 14740 30058 14792 30064
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14476 28206 14596 28234
rect 14568 28150 14596 28206
rect 14556 28144 14608 28150
rect 14556 28086 14608 28092
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14372 28076 14424 28082
rect 14372 28018 14424 28024
rect 14188 27940 14240 27946
rect 14188 27882 14240 27888
rect 14200 27538 14228 27882
rect 14188 27532 14240 27538
rect 14188 27474 14240 27480
rect 14384 27334 14412 28018
rect 14556 27940 14608 27946
rect 14556 27882 14608 27888
rect 14568 27606 14596 27882
rect 14660 27606 14688 28086
rect 14752 28082 14780 30058
rect 14924 29164 14976 29170
rect 14924 29106 14976 29112
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14556 27600 14608 27606
rect 14554 27568 14556 27577
rect 14648 27600 14700 27606
rect 14608 27568 14610 27577
rect 14648 27542 14700 27548
rect 14554 27503 14610 27512
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 14372 27328 14424 27334
rect 14186 27296 14242 27305
rect 14372 27270 14424 27276
rect 14186 27231 14242 27240
rect 13912 27056 13964 27062
rect 13912 26998 13964 27004
rect 14200 26926 14228 27231
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 14200 26518 14228 26862
rect 14188 26512 14240 26518
rect 14188 26454 14240 26460
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 13728 25968 13780 25974
rect 13728 25910 13780 25916
rect 13726 25392 13782 25401
rect 13726 25327 13728 25336
rect 13780 25327 13782 25336
rect 13728 25298 13780 25304
rect 14108 25294 14136 26318
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13556 23798 13584 24754
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 13648 24342 13676 24550
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13832 24206 13860 24754
rect 14108 24750 14136 25230
rect 14200 24750 14228 25230
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14094 24304 14150 24313
rect 14094 24239 14096 24248
rect 14148 24239 14150 24248
rect 14096 24210 14148 24216
rect 14200 24206 14228 24686
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13740 23730 13768 24074
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13464 23616 13584 23644
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 13358 21720 13414 21729
rect 13358 21655 13360 21664
rect 13412 21655 13414 21664
rect 13360 21626 13412 21632
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13372 20942 13400 21490
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13464 19786 13492 23122
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13280 19638 13492 19666
rect 13188 19230 13400 19258
rect 13084 19168 13136 19174
rect 12990 19136 13046 19145
rect 13084 19110 13136 19116
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 12990 19071 13046 19080
rect 13004 18698 13032 19071
rect 13096 18902 13124 19110
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 13084 18760 13136 18766
rect 13082 18728 13084 18737
rect 13136 18728 13138 18737
rect 12992 18692 13044 18698
rect 13082 18663 13138 18672
rect 12992 18634 13044 18640
rect 13004 18154 13032 18634
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18222 13124 18566
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 13096 17377 13124 17546
rect 13082 17368 13138 17377
rect 13082 17303 13138 17312
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12728 16918 12940 16946
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 13938 12480 14214
rect 12544 14074 12572 14894
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12544 13258 12572 13466
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12268 12434 12296 12650
rect 12176 12406 12296 12434
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 10810 11836 11018
rect 11992 10810 12020 11494
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 9926 12112 10610
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12084 9722 12112 9862
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11164 9042 11192 9454
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9178 12112 9318
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 7018 11008 7346
rect 11072 7274 11100 7822
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10888 6990 11008 7018
rect 11072 7002 11100 7210
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11060 6996 11112 7002
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10888 5234 10916 6990
rect 11060 6938 11112 6944
rect 11440 6798 11468 7142
rect 11532 7002 11560 7890
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11624 7410 11652 7822
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11624 6866 11652 7346
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10888 4622 10916 5170
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 11256 2650 11284 6598
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11624 5914 11652 6258
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11716 5574 11744 7278
rect 11900 6662 11928 8434
rect 11992 8430 12020 8910
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12176 8090 12204 12406
rect 12360 11830 12388 12786
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12452 11694 12480 13126
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12268 11354 12296 11494
rect 12452 11354 12480 11630
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 9722 12480 10950
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12636 9586 12664 16390
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12452 8838 12480 9114
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12176 7834 12204 8026
rect 12084 7806 12204 7834
rect 12084 6798 12112 7806
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 12084 6390 12112 6734
rect 12176 6390 12204 7686
rect 12268 7206 12296 7686
rect 12360 7342 12388 8230
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4486 11560 5102
rect 11716 4690 11744 5510
rect 12176 5166 12204 5646
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12268 5234 12296 5510
rect 12544 5370 12572 9386
rect 12636 8838 12664 9522
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12728 5846 12756 16918
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12820 16046 12848 16594
rect 13096 16522 13124 17138
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 12900 16448 12952 16454
rect 12898 16416 12900 16425
rect 12952 16416 12954 16425
rect 12898 16351 12954 16360
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12820 13394 12848 15982
rect 13004 15638 13032 16050
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13096 15745 13124 15982
rect 13082 15736 13138 15745
rect 13082 15671 13138 15680
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 15008 12940 15302
rect 13004 15162 13032 15574
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12992 15020 13044 15026
rect 12912 14980 12992 15008
rect 12992 14962 13044 14968
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12820 12238 12848 12582
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11898 12940 12038
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 11286 12848 11494
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12820 9926 12848 11018
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12912 9058 12940 9454
rect 12820 9042 12940 9058
rect 12808 9036 12940 9042
rect 12860 9030 12940 9036
rect 12808 8978 12860 8984
rect 12820 8090 12848 8978
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12820 6390 12848 8026
rect 13004 7954 13032 14962
rect 13096 14346 13124 15370
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13188 13326 13216 19110
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13280 17610 13308 18634
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 13372 17338 13400 19230
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 15026 13308 15438
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13280 14618 13308 14962
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13372 14074 13400 17274
rect 13464 17270 13492 19638
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13280 11830 13308 12242
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13280 11121 13308 11290
rect 13372 11150 13400 13330
rect 13464 11150 13492 14282
rect 13360 11144 13412 11150
rect 13266 11112 13322 11121
rect 13360 11086 13412 11092
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13266 11047 13322 11056
rect 13556 10742 13584 23616
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13648 19553 13676 23462
rect 13740 23254 13768 23666
rect 13832 23254 13860 24142
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 13910 23896 13966 23905
rect 13910 23831 13912 23840
rect 13964 23831 13966 23840
rect 13912 23802 13964 23808
rect 14016 23730 14044 24074
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 13820 23248 13872 23254
rect 13820 23190 13872 23196
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13740 22506 13768 23054
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13832 20618 13860 20742
rect 13740 20590 13860 20618
rect 13740 20466 13768 20590
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13818 19952 13874 19961
rect 13818 19887 13874 19896
rect 13634 19544 13690 19553
rect 13634 19479 13690 19488
rect 13648 19310 13676 19479
rect 13832 19378 13860 19887
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13634 19136 13690 19145
rect 13634 19071 13690 19080
rect 13648 18834 13676 19071
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13648 18290 13676 18566
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13740 18086 13768 18634
rect 13832 18222 13860 18702
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13726 16824 13782 16833
rect 13726 16759 13782 16768
rect 13740 16658 13768 16759
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13924 16182 13952 23530
rect 14200 23526 14228 24142
rect 14476 23866 14504 27406
rect 14752 27316 14780 28018
rect 14832 27328 14884 27334
rect 14752 27288 14832 27316
rect 14832 27270 14884 27276
rect 14556 26784 14608 26790
rect 14556 26726 14608 26732
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14200 23322 14228 23462
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14200 22420 14228 23054
rect 14292 22642 14320 23666
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 14280 22432 14332 22438
rect 14200 22392 14280 22420
rect 14280 22374 14332 22380
rect 14292 20602 14320 22374
rect 14568 22094 14596 26726
rect 14844 26489 14872 27270
rect 14830 26480 14886 26489
rect 14830 26415 14886 26424
rect 14936 26382 14964 29106
rect 15120 28234 15148 30670
rect 15304 30433 15332 31282
rect 15290 30424 15346 30433
rect 15290 30359 15346 30368
rect 15292 30252 15344 30258
rect 15396 30240 15424 34886
rect 15764 33998 15792 37810
rect 15948 37398 15976 37810
rect 16040 37466 16068 37810
rect 16028 37460 16080 37466
rect 16028 37402 16080 37408
rect 15936 37392 15988 37398
rect 15936 37334 15988 37340
rect 15948 37126 15976 37334
rect 15936 37120 15988 37126
rect 15936 37062 15988 37068
rect 16224 36786 16252 38150
rect 17512 37942 17540 38490
rect 20904 38412 20956 38418
rect 20956 38372 21036 38400
rect 20904 38354 20956 38360
rect 20168 38344 20220 38350
rect 20168 38286 20220 38292
rect 18696 38208 18748 38214
rect 18696 38150 18748 38156
rect 19892 38208 19944 38214
rect 19944 38168 20024 38196
rect 19892 38150 19944 38156
rect 18708 38010 18736 38150
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17868 38004 17920 38010
rect 17868 37946 17920 37952
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18788 38004 18840 38010
rect 18788 37946 18840 37952
rect 17500 37936 17552 37942
rect 17500 37878 17552 37884
rect 15844 36780 15896 36786
rect 15844 36722 15896 36728
rect 16212 36780 16264 36786
rect 16212 36722 16264 36728
rect 16304 36780 16356 36786
rect 16304 36722 16356 36728
rect 15752 33992 15804 33998
rect 15752 33934 15804 33940
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15476 31748 15528 31754
rect 15476 31690 15528 31696
rect 15488 30938 15516 31690
rect 15476 30932 15528 30938
rect 15476 30874 15528 30880
rect 15488 30598 15516 30874
rect 15672 30734 15700 32914
rect 15856 31498 15884 36722
rect 16224 36582 16252 36722
rect 16212 36576 16264 36582
rect 16212 36518 16264 36524
rect 16120 34672 16172 34678
rect 16120 34614 16172 34620
rect 16132 33998 16160 34614
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 16120 33992 16172 33998
rect 16120 33934 16172 33940
rect 15936 33924 15988 33930
rect 15936 33866 15988 33872
rect 15948 33318 15976 33866
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 15764 31470 15884 31498
rect 15660 30728 15712 30734
rect 15660 30670 15712 30676
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 15566 30560 15622 30569
rect 15566 30495 15622 30504
rect 15344 30212 15516 30240
rect 15292 30194 15344 30200
rect 15382 30016 15438 30025
rect 15304 29974 15382 30002
rect 15304 29646 15332 29974
rect 15382 29951 15438 29960
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15488 28529 15516 30212
rect 15580 29714 15608 30495
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 15568 29572 15620 29578
rect 15568 29514 15620 29520
rect 15580 29345 15608 29514
rect 15566 29336 15622 29345
rect 15566 29271 15622 29280
rect 15568 28756 15620 28762
rect 15568 28698 15620 28704
rect 15474 28520 15530 28529
rect 15474 28455 15530 28464
rect 15120 28206 15424 28234
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15212 27130 15240 28018
rect 15396 27985 15424 28206
rect 15382 27976 15438 27985
rect 15382 27911 15384 27920
rect 15436 27911 15438 27920
rect 15384 27882 15436 27888
rect 15488 27470 15516 28455
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15384 27396 15436 27402
rect 15384 27338 15436 27344
rect 15396 27169 15424 27338
rect 15382 27160 15438 27169
rect 15200 27124 15252 27130
rect 15382 27095 15438 27104
rect 15200 27066 15252 27072
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 14660 25906 14688 26318
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 14660 25294 14688 25842
rect 15120 25430 15148 25842
rect 15396 25498 15424 25978
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15108 25424 15160 25430
rect 15108 25366 15160 25372
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14660 24410 14688 25230
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14752 24342 14780 24754
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 15120 24274 15148 25366
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 15120 23186 15148 24210
rect 15396 24206 15424 25434
rect 15580 24936 15608 28698
rect 15672 27538 15700 30670
rect 15764 29646 15792 31470
rect 15948 30716 15976 33254
rect 16040 31754 16068 33934
rect 16132 33590 16160 33934
rect 16120 33584 16172 33590
rect 16120 33526 16172 33532
rect 16316 32978 16344 36722
rect 17224 36712 17276 36718
rect 17224 36654 17276 36660
rect 17132 36236 17184 36242
rect 17132 36178 17184 36184
rect 17144 35834 17172 36178
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 17236 34678 17264 36654
rect 17500 36372 17552 36378
rect 17500 36314 17552 36320
rect 17408 36032 17460 36038
rect 17408 35974 17460 35980
rect 17420 35154 17448 35974
rect 17512 35222 17540 36314
rect 17696 36174 17724 37946
rect 17880 37466 17908 37946
rect 18144 37868 18196 37874
rect 18144 37810 18196 37816
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 17868 37460 17920 37466
rect 17868 37402 17920 37408
rect 18052 37324 18104 37330
rect 18052 37266 18104 37272
rect 17776 36304 17828 36310
rect 17774 36272 17776 36281
rect 17828 36272 17830 36281
rect 17774 36207 17830 36216
rect 17684 36168 17736 36174
rect 17684 36110 17736 36116
rect 17776 36168 17828 36174
rect 17776 36110 17828 36116
rect 17500 35216 17552 35222
rect 17500 35158 17552 35164
rect 17408 35148 17460 35154
rect 17408 35090 17460 35096
rect 16764 34672 16816 34678
rect 16764 34614 16816 34620
rect 17224 34672 17276 34678
rect 17224 34614 17276 34620
rect 16672 34468 16724 34474
rect 16672 34410 16724 34416
rect 16396 34400 16448 34406
rect 16396 34342 16448 34348
rect 16408 33402 16436 34342
rect 16684 33998 16712 34410
rect 16488 33992 16540 33998
rect 16672 33992 16724 33998
rect 16540 33952 16620 33980
rect 16488 33934 16540 33940
rect 16486 33416 16542 33425
rect 16408 33374 16486 33402
rect 16486 33351 16542 33360
rect 16304 32972 16356 32978
rect 16304 32914 16356 32920
rect 16304 32836 16356 32842
rect 16304 32778 16356 32784
rect 16316 31754 16344 32778
rect 16592 32201 16620 33952
rect 16672 33934 16724 33940
rect 16578 32192 16634 32201
rect 16578 32127 16634 32136
rect 16486 31920 16542 31929
rect 16486 31855 16542 31864
rect 16040 31726 16160 31754
rect 16028 30728 16080 30734
rect 15948 30688 16028 30716
rect 16028 30670 16080 30676
rect 15842 30016 15898 30025
rect 15842 29951 15898 29960
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15660 27532 15712 27538
rect 15660 27474 15712 27480
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 15672 26994 15700 27270
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15660 26512 15712 26518
rect 15660 26454 15712 26460
rect 15488 24908 15608 24936
rect 15488 24342 15516 24908
rect 15566 24848 15622 24857
rect 15566 24783 15622 24792
rect 15476 24336 15528 24342
rect 15476 24278 15528 24284
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 15304 23798 15332 24142
rect 15292 23792 15344 23798
rect 15580 23769 15608 24783
rect 15672 24188 15700 26454
rect 15764 26314 15792 27406
rect 15856 26994 15884 29951
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15948 27402 15976 29446
rect 16040 28966 16068 30670
rect 16132 29646 16160 31726
rect 16304 31748 16356 31754
rect 16304 31690 16356 31696
rect 16212 31136 16264 31142
rect 16212 31078 16264 31084
rect 16120 29640 16172 29646
rect 16120 29582 16172 29588
rect 16028 28960 16080 28966
rect 16028 28902 16080 28908
rect 16132 28121 16160 29582
rect 16224 29578 16252 31078
rect 16212 29572 16264 29578
rect 16212 29514 16264 29520
rect 16316 29492 16344 31690
rect 16396 29504 16448 29510
rect 16316 29464 16396 29492
rect 16396 29446 16448 29452
rect 16304 29300 16356 29306
rect 16304 29242 16356 29248
rect 16212 29232 16264 29238
rect 16210 29200 16212 29209
rect 16264 29200 16266 29209
rect 16210 29135 16266 29144
rect 16212 29028 16264 29034
rect 16212 28970 16264 28976
rect 16118 28112 16174 28121
rect 16118 28047 16120 28056
rect 16172 28047 16174 28056
rect 16120 28018 16172 28024
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15948 26874 15976 27338
rect 16040 26994 16068 27406
rect 16120 27056 16172 27062
rect 16120 26998 16172 27004
rect 16028 26988 16080 26994
rect 16028 26930 16080 26936
rect 15856 26846 15976 26874
rect 15752 26308 15804 26314
rect 15752 26250 15804 26256
rect 15752 24200 15804 24206
rect 15672 24160 15752 24188
rect 15856 24177 15884 26846
rect 16132 25906 16160 26998
rect 16224 26228 16252 28970
rect 16316 27946 16344 29242
rect 16304 27940 16356 27946
rect 16304 27882 16356 27888
rect 16408 26382 16436 29446
rect 16500 28150 16528 31855
rect 16592 31414 16620 32127
rect 16776 31736 16804 34614
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 16948 34536 17000 34542
rect 17328 34490 17356 34546
rect 16948 34478 17000 34484
rect 16856 34400 16908 34406
rect 16856 34342 16908 34348
rect 16868 34202 16896 34342
rect 16960 34202 16988 34478
rect 17236 34462 17356 34490
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16948 34196 17000 34202
rect 16948 34138 17000 34144
rect 16854 34096 16910 34105
rect 16854 34031 16910 34040
rect 16868 33522 16896 34031
rect 16948 33992 17000 33998
rect 16948 33934 17000 33940
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16868 31822 16896 33458
rect 16960 32774 16988 33934
rect 17236 33862 17264 34462
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 17224 33856 17276 33862
rect 17224 33798 17276 33804
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 17144 33114 17172 33798
rect 17132 33108 17184 33114
rect 17132 33050 17184 33056
rect 17236 32842 17264 33798
rect 17328 33454 17356 33798
rect 17420 33590 17448 35090
rect 17512 33590 17540 35158
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17408 33584 17460 33590
rect 17408 33526 17460 33532
rect 17500 33584 17552 33590
rect 17500 33526 17552 33532
rect 17316 33448 17368 33454
rect 17408 33448 17460 33454
rect 17316 33390 17368 33396
rect 17406 33416 17408 33425
rect 17460 33416 17462 33425
rect 17406 33351 17462 33360
rect 17696 33114 17724 34546
rect 17788 33522 17816 36110
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 17880 34105 17908 34546
rect 17866 34096 17922 34105
rect 17866 34031 17922 34040
rect 18064 33998 18092 37266
rect 18156 36174 18184 37810
rect 18236 37392 18288 37398
rect 18236 37334 18288 37340
rect 18248 36922 18276 37334
rect 18236 36916 18288 36922
rect 18236 36858 18288 36864
rect 18524 36582 18552 37810
rect 18800 37126 18828 37946
rect 19996 37942 20024 38168
rect 20180 38010 20208 38286
rect 20168 38004 20220 38010
rect 20168 37946 20220 37952
rect 19984 37936 20036 37942
rect 19984 37878 20036 37884
rect 18880 37868 18932 37874
rect 18880 37810 18932 37816
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 19156 37868 19208 37874
rect 19156 37810 19208 37816
rect 18788 37120 18840 37126
rect 18788 37062 18840 37068
rect 18512 36576 18564 36582
rect 18512 36518 18564 36524
rect 18328 36372 18380 36378
rect 18328 36314 18380 36320
rect 18420 36372 18472 36378
rect 18420 36314 18472 36320
rect 18340 36242 18368 36314
rect 18328 36236 18380 36242
rect 18328 36178 18380 36184
rect 18144 36168 18196 36174
rect 18196 36116 18368 36122
rect 18144 36110 18368 36116
rect 18156 36094 18368 36110
rect 18340 35737 18368 36094
rect 18326 35728 18382 35737
rect 18326 35663 18382 35672
rect 18236 34944 18288 34950
rect 18236 34886 18288 34892
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 17868 33924 17920 33930
rect 17868 33866 17920 33872
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17224 32836 17276 32842
rect 17224 32778 17276 32784
rect 16948 32768 17000 32774
rect 16948 32710 17000 32716
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 16684 31708 16804 31736
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 16592 30802 16620 31214
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16592 30190 16620 30534
rect 16684 30326 16712 31708
rect 16960 31668 16988 32710
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 16776 31640 16988 31668
rect 16776 30938 16804 31640
rect 16948 31408 17000 31414
rect 16868 31356 16948 31362
rect 16868 31350 17000 31356
rect 16868 31334 16988 31350
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16488 28144 16540 28150
rect 16488 28086 16540 28092
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16500 26790 16528 27406
rect 16488 26784 16540 26790
rect 16488 26726 16540 26732
rect 16592 26382 16620 29582
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16684 29034 16712 29446
rect 16672 29028 16724 29034
rect 16672 28970 16724 28976
rect 16776 28540 16804 30874
rect 16868 29730 16896 31334
rect 16948 31272 17000 31278
rect 16948 31214 17000 31220
rect 16960 30938 16988 31214
rect 17040 31136 17092 31142
rect 17040 31078 17092 31084
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 17052 30870 17080 31078
rect 17040 30864 17092 30870
rect 17040 30806 17092 30812
rect 16948 30660 17000 30666
rect 16948 30602 17000 30608
rect 16960 30410 16988 30602
rect 16960 30382 17080 30410
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16960 29850 16988 30194
rect 16948 29844 17000 29850
rect 16948 29786 17000 29792
rect 16868 29702 16988 29730
rect 16856 28552 16908 28558
rect 16776 28512 16856 28540
rect 16856 28494 16908 28500
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16684 27130 16712 27406
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16776 26994 16804 27814
rect 16868 27130 16896 28494
rect 16960 27130 16988 29702
rect 17052 27538 17080 30382
rect 17144 29646 17172 31758
rect 17420 31210 17448 33050
rect 17592 32768 17644 32774
rect 17592 32710 17644 32716
rect 17604 31929 17632 32710
rect 17590 31920 17646 31929
rect 17590 31855 17646 31864
rect 17604 31414 17632 31855
rect 17592 31408 17644 31414
rect 17788 31385 17816 33458
rect 17880 32978 17908 33866
rect 17972 33386 18000 33866
rect 17960 33380 18012 33386
rect 17960 33322 18012 33328
rect 17868 32972 17920 32978
rect 17868 32914 17920 32920
rect 17972 32910 18000 33322
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 17960 32768 18012 32774
rect 17960 32710 18012 32716
rect 17972 31668 18000 32710
rect 18064 31754 18092 33934
rect 18248 32994 18276 34886
rect 18328 33312 18380 33318
rect 18328 33254 18380 33260
rect 18340 33114 18368 33254
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 18248 32966 18368 32994
rect 18236 32904 18288 32910
rect 18156 32881 18236 32892
rect 18142 32872 18236 32881
rect 18198 32864 18236 32872
rect 18236 32846 18288 32852
rect 18142 32807 18198 32816
rect 18248 32434 18276 32846
rect 18340 32434 18368 32966
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18236 32224 18288 32230
rect 18236 32166 18288 32172
rect 18248 32065 18276 32166
rect 18234 32056 18290 32065
rect 18234 31991 18290 32000
rect 18064 31726 18368 31754
rect 17972 31640 18092 31668
rect 17592 31350 17644 31356
rect 17774 31376 17830 31385
rect 17500 31340 17552 31346
rect 17774 31311 17830 31320
rect 17500 31282 17552 31288
rect 17408 31204 17460 31210
rect 17408 31146 17460 31152
rect 17224 30864 17276 30870
rect 17224 30806 17276 30812
rect 17236 30734 17264 30806
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17328 30394 17356 30534
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 17224 30252 17276 30258
rect 17276 30212 17356 30240
rect 17224 30194 17276 30200
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 17224 28960 17276 28966
rect 17224 28902 17276 28908
rect 17236 28558 17264 28902
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17236 27878 17264 28494
rect 17224 27872 17276 27878
rect 17224 27814 17276 27820
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16304 26240 16356 26246
rect 16224 26200 16304 26228
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 16028 25764 16080 25770
rect 16028 25706 16080 25712
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 15948 24857 15976 24890
rect 15934 24848 15990 24857
rect 15934 24783 15990 24792
rect 15752 24142 15804 24148
rect 15842 24168 15898 24177
rect 15292 23734 15344 23740
rect 15566 23760 15622 23769
rect 15200 23724 15252 23730
rect 15566 23695 15622 23704
rect 15200 23666 15252 23672
rect 15108 23180 15160 23186
rect 15108 23122 15160 23128
rect 15212 23066 15240 23666
rect 15580 23662 15608 23695
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15028 23038 15240 23066
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15028 22982 15056 23038
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 15016 22772 15068 22778
rect 15120 22760 15148 22918
rect 15068 22732 15148 22760
rect 15016 22714 15068 22720
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 14568 22066 14688 22094
rect 14464 21004 14516 21010
rect 14516 20964 14596 20992
rect 14464 20946 14516 20952
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14108 20058 14136 20402
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14016 19145 14044 19994
rect 14002 19136 14058 19145
rect 14002 19071 14058 19080
rect 14200 17542 14228 20538
rect 14384 20466 14412 20742
rect 14568 20466 14596 20964
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14278 20088 14334 20097
rect 14278 20023 14334 20032
rect 14292 19854 14320 20023
rect 14384 19990 14412 20402
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14280 19848 14332 19854
rect 14476 19802 14504 20334
rect 14568 20262 14596 20402
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14280 19790 14332 19796
rect 14384 19774 14504 19802
rect 14384 18698 14412 19774
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13004 7342 13032 7890
rect 13096 7886 13124 9522
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13280 8294 13308 8978
rect 13556 8906 13584 9862
rect 13648 9110 13676 12718
rect 13924 12434 13952 14554
rect 13832 12406 13952 12434
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13740 10606 13768 11018
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13832 9518 13860 12406
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13924 10606 13952 11630
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13832 8634 13860 9318
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13280 7954 13308 8230
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7546 13308 7686
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 6458 13216 6734
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 13188 5914 13216 6394
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 12452 4282 12480 4490
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12820 4146 12848 5510
rect 13096 5302 13124 5850
rect 13556 5778 13584 6054
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13648 5370 13676 6190
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 13096 4214 13124 5238
rect 13648 5148 13676 5306
rect 13740 5234 13768 6258
rect 14016 6118 14044 17478
rect 14384 17338 14412 18634
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14108 11014 14136 12854
rect 14200 11354 14228 16934
rect 14384 16658 14412 16934
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14568 16454 14596 17614
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14476 15570 14504 16390
rect 14568 15706 14596 16390
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 14618 14412 15302
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14568 13326 14596 13466
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14660 12434 14688 22066
rect 14752 21146 14780 22578
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14936 21554 14964 21830
rect 15028 21554 15056 22578
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14752 20602 14780 20810
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14752 20330 14780 20538
rect 14936 20346 14964 21490
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15028 20482 15056 20878
rect 15120 20602 15148 22732
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15212 22030 15240 22442
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15212 21622 15240 21966
rect 15200 21616 15252 21622
rect 15200 21558 15252 21564
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15028 20466 15148 20482
rect 15028 20460 15160 20466
rect 15028 20454 15108 20460
rect 15108 20402 15160 20408
rect 14740 20324 14792 20330
rect 14936 20318 15056 20346
rect 14740 20266 14792 20272
rect 14752 19922 14780 20266
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14936 19281 14964 19314
rect 14922 19272 14978 19281
rect 14922 19207 14978 19216
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 14936 18698 14964 19110
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14936 18057 14964 18634
rect 14922 18048 14978 18057
rect 14922 17983 14978 17992
rect 15028 17678 15056 20318
rect 15120 20058 15148 20402
rect 15212 20330 15240 20742
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15212 19514 15240 19858
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15120 19310 15148 19450
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15304 17814 15332 23054
rect 15764 22710 15792 24142
rect 15842 24103 15898 24112
rect 15844 24064 15896 24070
rect 15842 24032 15844 24041
rect 15896 24032 15898 24041
rect 15842 23967 15898 23976
rect 15948 23798 15976 24783
rect 16040 24682 16068 25706
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16028 24676 16080 24682
rect 16028 24618 16080 24624
rect 16040 24206 16068 24618
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15856 23633 15884 23666
rect 15842 23624 15898 23633
rect 15842 23559 15898 23568
rect 16040 23254 16068 24142
rect 16132 23594 16160 24754
rect 16224 24290 16252 26200
rect 16304 26182 16356 26188
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16316 24410 16344 24754
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16224 24274 16344 24290
rect 16224 24268 16356 24274
rect 16224 24262 16304 24268
rect 16304 24210 16356 24216
rect 16120 23588 16172 23594
rect 16120 23530 16172 23536
rect 16212 23588 16264 23594
rect 16212 23530 16264 23536
rect 16028 23248 16080 23254
rect 16028 23190 16080 23196
rect 16224 23118 16252 23530
rect 16316 23254 16344 24210
rect 16408 24206 16436 26318
rect 16592 25786 16620 26318
rect 16592 25758 16712 25786
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16592 25265 16620 25638
rect 16684 25294 16712 25758
rect 16672 25288 16724 25294
rect 16578 25256 16634 25265
rect 16672 25230 16724 25236
rect 16578 25191 16634 25200
rect 16684 24818 16712 25230
rect 16776 25226 16804 26930
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16672 24812 16724 24818
rect 16724 24772 16804 24800
rect 16672 24754 16724 24760
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16500 23497 16528 24550
rect 16486 23488 16542 23497
rect 16486 23423 16542 23432
rect 16304 23248 16356 23254
rect 16304 23190 16356 23196
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16212 23112 16264 23118
rect 16212 23054 16264 23060
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15396 22166 15424 22578
rect 15384 22160 15436 22166
rect 15384 22102 15436 22108
rect 15488 21690 15516 22578
rect 15856 22098 15884 22578
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 16408 21622 16436 23054
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15672 20466 15700 20742
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15488 19786 15516 20402
rect 15672 19990 15700 20402
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15660 19848 15712 19854
rect 15764 19836 15792 20810
rect 16040 20806 16068 21490
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15856 19990 15884 20266
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15712 19808 15792 19836
rect 15660 19790 15712 19796
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15488 19378 15516 19722
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15476 19372 15528 19378
rect 15396 19320 15476 19334
rect 15396 19314 15528 19320
rect 15396 19306 15516 19314
rect 15396 18766 15424 19306
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15396 17882 15424 18702
rect 15580 18426 15608 19450
rect 15672 18766 15700 19790
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15568 18420 15620 18426
rect 15856 18408 15884 19926
rect 16040 19854 16068 20742
rect 16224 20262 16252 21490
rect 16500 20942 16528 22442
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19334 16068 19790
rect 16040 19306 16160 19334
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 16040 18426 16068 18634
rect 15568 18362 15620 18368
rect 15672 18380 15884 18408
rect 16028 18420 16080 18426
rect 15568 18148 15620 18154
rect 15568 18090 15620 18096
rect 15580 17921 15608 18090
rect 15566 17912 15622 17921
rect 15384 17876 15436 17882
rect 15566 17847 15622 17856
rect 15384 17818 15436 17824
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14752 15570 14780 15642
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14752 13938 14780 15506
rect 14844 15026 14872 16458
rect 15028 15570 15056 17614
rect 15212 17134 15240 17614
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15304 16590 15332 17206
rect 15396 17202 15424 17478
rect 15384 17196 15436 17202
rect 15580 17184 15608 17750
rect 15672 17678 15700 18380
rect 16028 18362 16080 18368
rect 16132 18290 16160 19306
rect 15752 18284 15804 18290
rect 15936 18284 15988 18290
rect 15804 18244 15884 18272
rect 15752 18226 15804 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 17678 15792 18022
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15856 17270 15884 18244
rect 16120 18284 16172 18290
rect 15988 18244 16068 18272
rect 15936 18226 15988 18232
rect 16040 17542 16068 18244
rect 16120 18226 16172 18232
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15752 17196 15804 17202
rect 15580 17156 15752 17184
rect 15384 17138 15436 17144
rect 15752 17138 15804 17144
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 15396 14890 15424 16730
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 15570 15516 16594
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 15586 15700 16458
rect 15764 15858 15792 17138
rect 15842 15872 15898 15881
rect 15764 15830 15842 15858
rect 15842 15807 15898 15816
rect 15842 15600 15898 15609
rect 15476 15564 15528 15570
rect 15672 15558 15842 15586
rect 15842 15535 15898 15544
rect 15476 15506 15528 15512
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15028 14414 15056 14758
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 14074 14872 14214
rect 14936 14074 14964 14350
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15028 13530 15056 13874
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15212 13326 15240 14758
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15304 14074 15332 14350
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15200 13320 15252 13326
rect 15396 13308 15424 14826
rect 15488 14618 15516 15506
rect 15856 15502 15884 15535
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15672 15094 15700 15302
rect 15856 15201 15884 15302
rect 15842 15192 15898 15201
rect 15842 15127 15898 15136
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15750 15056 15806 15065
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13462 15516 13874
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15672 13326 15700 15030
rect 15750 14991 15752 15000
rect 15804 14991 15806 15000
rect 15752 14962 15804 14968
rect 15764 14550 15792 14962
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15948 14414 15976 17478
rect 16040 17202 16068 17478
rect 16132 17338 16160 18226
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16224 16046 16252 20198
rect 16316 18426 16344 20878
rect 16592 20874 16620 21082
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16592 20534 16620 20810
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16500 18766 16528 19790
rect 16578 19544 16634 19553
rect 16578 19479 16580 19488
rect 16632 19479 16634 19488
rect 16580 19450 16632 19456
rect 16684 19334 16712 23122
rect 16776 22166 16804 24772
rect 16868 24070 16896 27066
rect 16960 24274 16988 27066
rect 17052 25430 17080 27474
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17144 26382 17172 27270
rect 17328 26382 17356 30212
rect 17420 29510 17448 31146
rect 17512 29850 17540 31282
rect 17684 31136 17736 31142
rect 17684 31078 17736 31084
rect 17696 30977 17724 31078
rect 17682 30968 17738 30977
rect 17682 30903 17738 30912
rect 17592 30864 17644 30870
rect 17788 30818 17816 31311
rect 17960 31204 18012 31210
rect 17960 31146 18012 31152
rect 17644 30812 17816 30818
rect 17592 30806 17816 30812
rect 17868 30864 17920 30870
rect 17868 30806 17920 30812
rect 17604 30790 17816 30806
rect 17788 30376 17816 30790
rect 17880 30569 17908 30806
rect 17866 30560 17922 30569
rect 17866 30495 17922 30504
rect 17788 30348 17908 30376
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 17512 28082 17540 29786
rect 17408 28076 17460 28082
rect 17408 28018 17460 28024
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 17420 27577 17448 28018
rect 17406 27568 17462 27577
rect 17406 27503 17462 27512
rect 17420 27470 17448 27503
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17696 26382 17724 30194
rect 17880 28422 17908 30348
rect 17972 30326 18000 31146
rect 18064 30598 18092 31640
rect 18144 31272 18196 31278
rect 18144 31214 18196 31220
rect 18156 30734 18184 31214
rect 18236 31136 18288 31142
rect 18236 31078 18288 31084
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18052 30592 18104 30598
rect 18052 30534 18104 30540
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 18248 30258 18276 31078
rect 18340 30841 18368 31726
rect 18432 31226 18460 36314
rect 18524 36174 18552 36518
rect 18604 36304 18656 36310
rect 18602 36272 18604 36281
rect 18656 36272 18658 36281
rect 18602 36207 18658 36216
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18604 36100 18656 36106
rect 18604 36042 18656 36048
rect 18616 35698 18644 36042
rect 18708 35834 18736 36178
rect 18800 36174 18828 37062
rect 18892 36854 18920 37810
rect 19076 37398 19104 37810
rect 19064 37392 19116 37398
rect 19064 37334 19116 37340
rect 19168 37126 19196 37810
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 19800 37664 19852 37670
rect 19800 37606 19852 37612
rect 19352 37330 19380 37606
rect 19340 37324 19392 37330
rect 19340 37266 19392 37272
rect 19812 37262 19840 37606
rect 19800 37256 19852 37262
rect 19800 37198 19852 37204
rect 19432 37188 19484 37194
rect 19432 37130 19484 37136
rect 19156 37120 19208 37126
rect 19076 37080 19156 37108
rect 18880 36848 18932 36854
rect 18880 36790 18932 36796
rect 18892 36174 18920 36790
rect 18788 36168 18840 36174
rect 18788 36110 18840 36116
rect 18880 36168 18932 36174
rect 18880 36110 18932 36116
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18604 35692 18656 35698
rect 18604 35634 18656 35640
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18524 33658 18552 33798
rect 18512 33652 18564 33658
rect 18512 33594 18564 33600
rect 18616 32314 18644 35634
rect 18786 33824 18842 33833
rect 18786 33759 18842 33768
rect 18800 33522 18828 33759
rect 18788 33516 18840 33522
rect 18788 33458 18840 33464
rect 18880 33448 18932 33454
rect 18880 33390 18932 33396
rect 18892 32978 18920 33390
rect 18880 32972 18932 32978
rect 18880 32914 18932 32920
rect 18972 32972 19024 32978
rect 18972 32914 19024 32920
rect 18696 32836 18748 32842
rect 18696 32778 18748 32784
rect 18708 32434 18736 32778
rect 18696 32428 18748 32434
rect 18696 32370 18748 32376
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 18616 32286 18736 32314
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18616 31346 18644 31962
rect 18708 31346 18736 32286
rect 18788 31680 18840 31686
rect 18788 31622 18840 31628
rect 18604 31340 18656 31346
rect 18604 31282 18656 31288
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18432 31198 18644 31226
rect 18420 31136 18472 31142
rect 18420 31078 18472 31084
rect 18326 30832 18382 30841
rect 18326 30767 18382 30776
rect 18328 30660 18380 30666
rect 18432 30648 18460 31078
rect 18380 30620 18460 30648
rect 18512 30660 18564 30666
rect 18328 30602 18380 30608
rect 18512 30602 18564 30608
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17972 29646 18000 29990
rect 17960 29640 18012 29646
rect 18340 29628 18368 30602
rect 18420 30388 18472 30394
rect 18420 30330 18472 30336
rect 18432 29696 18460 30330
rect 18524 30054 18552 30602
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 18512 29708 18564 29714
rect 18432 29668 18512 29696
rect 18512 29650 18564 29656
rect 18340 29600 18460 29628
rect 17960 29582 18012 29588
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 17972 29306 18000 29446
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 18050 29064 18106 29073
rect 18050 28999 18052 29008
rect 18104 28999 18106 29008
rect 18052 28970 18104 28976
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17868 28416 17920 28422
rect 17868 28358 17920 28364
rect 17776 28144 17828 28150
rect 17776 28086 17828 28092
rect 17788 26382 17816 28086
rect 17880 27538 17908 28358
rect 17972 28218 18000 28494
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17040 25424 17092 25430
rect 17040 25366 17092 25372
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 17144 24449 17172 24686
rect 17130 24440 17186 24449
rect 17130 24375 17186 24384
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 22574 16896 24006
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16960 23050 16988 23258
rect 17052 23186 17080 23598
rect 17236 23594 17264 25094
rect 17696 24698 17724 26318
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 17972 24818 18000 25774
rect 18064 24818 18092 27270
rect 18156 27130 18184 28018
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18156 25294 18184 26182
rect 18248 25906 18276 29446
rect 18432 28801 18460 29600
rect 18512 29504 18564 29510
rect 18512 29446 18564 29452
rect 18524 29170 18552 29446
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18418 28792 18474 28801
rect 18418 28727 18474 28736
rect 18432 27614 18460 28727
rect 18340 27586 18460 27614
rect 18340 26994 18368 27586
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 18432 26382 18460 26930
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17866 24712 17922 24721
rect 17696 24670 17866 24698
rect 17866 24647 17922 24656
rect 17880 24410 17908 24647
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 17316 24132 17368 24138
rect 17316 24074 17368 24080
rect 17224 23588 17276 23594
rect 17224 23530 17276 23536
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 17328 22964 17356 24074
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17420 23118 17448 23666
rect 17592 23248 17644 23254
rect 17776 23248 17828 23254
rect 17644 23208 17776 23236
rect 17592 23190 17644 23196
rect 17776 23190 17828 23196
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17328 22936 17448 22964
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 16856 22568 16908 22574
rect 17132 22568 17184 22574
rect 16856 22510 16908 22516
rect 16960 22528 17132 22556
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16856 22024 16908 22030
rect 16960 22012 16988 22528
rect 17132 22510 17184 22516
rect 17328 22094 17356 22578
rect 17144 22066 17356 22094
rect 17144 22030 17172 22066
rect 16908 21984 16988 22012
rect 16856 21966 16908 21972
rect 16776 21690 16804 21966
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16776 20602 16804 21354
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16868 19689 16896 19790
rect 16854 19680 16910 19689
rect 16854 19615 16910 19624
rect 16684 19306 16804 19334
rect 16776 18834 16804 19306
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16316 18086 16344 18362
rect 16500 18222 16528 18362
rect 16592 18222 16620 18770
rect 16868 18766 16896 19615
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16316 17082 16344 18022
rect 16500 17678 16528 18158
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16408 17270 16436 17614
rect 16592 17610 16620 18158
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16500 17202 16528 17274
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16316 17054 16436 17082
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15856 14074 15884 14282
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 14074 15976 14214
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16040 13734 16068 15982
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15570 16252 15846
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16132 15162 16160 15370
rect 16224 15162 16252 15506
rect 16316 15434 16344 16934
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16302 15328 16358 15337
rect 16302 15263 16358 15272
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16224 14414 16252 15098
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 13938 16160 14214
rect 16316 13938 16344 15263
rect 16408 15162 16436 17054
rect 16500 16794 16528 17138
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16500 15570 16528 16526
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16592 15450 16620 17546
rect 16684 17338 16712 17682
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16500 15422 16620 15450
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16500 14822 16528 15422
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16592 14482 16620 15302
rect 16684 14890 16712 17070
rect 16776 16590 16804 18158
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16868 15978 16896 18702
rect 16960 17882 16988 21984
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 17052 19922 17080 20334
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16960 17202 16988 17546
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16854 15872 16910 15881
rect 16854 15807 16910 15816
rect 16868 15502 16896 15807
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15476 13320 15528 13326
rect 15396 13280 15476 13308
rect 15200 13262 15252 13268
rect 15476 13262 15528 13268
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15028 12986 15056 13262
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14660 12406 14872 12434
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10810 14136 10950
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14200 10266 14228 11290
rect 14660 10674 14688 11494
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14464 10600 14516 10606
rect 14660 10554 14688 10610
rect 14464 10542 14516 10548
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14384 10062 14412 10542
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14292 8974 14320 9658
rect 14476 9058 14504 10542
rect 14384 9030 14504 9058
rect 14568 10526 14780 10554
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14292 8090 14320 8434
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14384 8022 14412 9030
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14476 7886 14504 8910
rect 14568 8634 14596 10526
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14660 10062 14688 10406
rect 14752 10130 14780 10526
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9722 14780 9862
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14660 8566 14688 8774
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14752 8294 14780 9522
rect 14844 9450 14872 12406
rect 14936 11830 14964 12786
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15028 11558 15056 11834
rect 15120 11778 15148 12378
rect 15212 12306 15240 13262
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15212 11898 15240 12038
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15120 11750 15240 11778
rect 15016 11552 15068 11558
rect 15068 11512 15148 11540
rect 15016 11494 15068 11500
rect 14924 11144 14976 11150
rect 14976 11104 15056 11132
rect 14924 11086 14976 11092
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14936 10266 14964 10678
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15028 9761 15056 11104
rect 15014 9752 15070 9761
rect 15014 9687 15070 9696
rect 15028 9518 15056 9687
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15028 8906 15056 9114
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 7954 14780 8230
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14292 7274 14320 7414
rect 14844 7342 14872 7890
rect 15120 7478 15148 11512
rect 15212 9586 15240 11750
rect 15304 11354 15332 12038
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15212 8430 15240 8774
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15304 7546 15332 11290
rect 15396 11218 15424 12718
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15488 11150 15516 13262
rect 16040 12918 16068 13670
rect 16132 12986 16160 13874
rect 16592 13870 16620 14418
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16684 13462 16712 14826
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16776 14113 16804 14554
rect 16762 14104 16818 14113
rect 16762 14039 16818 14048
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16776 13326 16804 14039
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16868 12850 16896 15438
rect 16960 15026 16988 16118
rect 17052 15094 17080 19858
rect 17144 19242 17172 21966
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17236 20466 17264 21354
rect 17328 21146 17356 21422
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 17328 20534 17356 21082
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17420 20058 17448 22936
rect 17512 21146 17540 22986
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17604 22098 17632 22510
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 17604 21554 17632 22034
rect 17696 21690 17724 22578
rect 18064 22556 18092 24142
rect 18156 23526 18184 24754
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18156 22710 18184 23462
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 18064 22528 18184 22556
rect 18156 22030 18184 22528
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17604 21010 17632 21286
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17696 20924 17724 21286
rect 17788 21146 17816 21490
rect 17972 21418 18000 21490
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17880 21078 17908 21286
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17972 20942 18000 21354
rect 17776 20936 17828 20942
rect 17696 20896 17776 20924
rect 17776 20878 17828 20884
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17696 20534 17724 20742
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17592 19848 17644 19854
rect 17696 19836 17724 20334
rect 17644 19808 17724 19836
rect 17592 19790 17644 19796
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17132 19236 17184 19242
rect 17184 19196 17264 19224
rect 17132 19178 17184 19184
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17144 18426 17172 18702
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17144 16998 17172 18022
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17236 15722 17264 19196
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17512 18766 17540 19110
rect 17604 18970 17632 19382
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17604 18290 17632 18702
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17512 17338 17540 18158
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17144 15706 17264 15722
rect 17132 15700 17264 15706
rect 17184 15694 17264 15700
rect 17132 15642 17184 15648
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 17236 14958 17264 15694
rect 17328 15366 17356 16390
rect 17512 16114 17540 16934
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17408 15700 17460 15706
rect 17512 15688 17540 16050
rect 17460 15660 17540 15688
rect 17408 15642 17460 15648
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17236 14414 17264 14894
rect 17512 14482 17540 15030
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17512 12850 17540 13262
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 12306 15608 12718
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11558 15608 12038
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15580 10742 15608 11494
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15672 10810 15700 10950
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15580 10130 15608 10678
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15580 9994 15608 10066
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15108 7472 15160 7478
rect 15028 7420 15108 7426
rect 15028 7414 15160 7420
rect 15028 7398 15148 7414
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5710 14044 6054
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14476 5370 14504 5578
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13556 5120 13676 5148
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4282 13308 4966
rect 13464 4622 13492 5034
rect 13556 4826 13584 5120
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13648 4622 13676 4966
rect 13740 4842 13768 5170
rect 13740 4826 13860 4842
rect 13740 4820 13872 4826
rect 13740 4814 13820 4820
rect 13820 4762 13872 4768
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 15028 4554 15056 7398
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6798 15240 7142
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15120 5778 15148 6054
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15212 5250 15240 6122
rect 15304 5370 15332 6734
rect 15764 6186 15792 12650
rect 17604 12434 17632 16390
rect 17696 16232 17724 19808
rect 17788 19242 17816 20878
rect 17866 20088 17922 20097
rect 17866 20023 17922 20032
rect 17880 19922 17908 20023
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17880 19689 17908 19722
rect 17866 19680 17922 19689
rect 17866 19615 17922 19624
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17788 17377 17816 18906
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17880 18086 17908 18634
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17774 17368 17830 17377
rect 17774 17303 17830 17312
rect 17788 16980 17816 17303
rect 17972 17134 18000 20878
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 18064 18698 18092 20334
rect 18156 18970 18184 21966
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18156 18408 18184 18770
rect 18064 18380 18184 18408
rect 18064 18222 18092 18380
rect 18052 18216 18104 18222
rect 18104 18176 18184 18204
rect 18052 18158 18104 18164
rect 18156 17678 18184 18176
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17788 16952 18092 16980
rect 17958 16552 18014 16561
rect 17958 16487 17960 16496
rect 18012 16487 18014 16496
rect 17960 16458 18012 16464
rect 17696 16204 17908 16232
rect 17880 16114 17908 16204
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17696 15416 17724 16050
rect 17788 15706 17816 16050
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17880 15609 17908 16050
rect 18064 15706 18092 16952
rect 18156 16794 18184 17614
rect 18248 17270 18276 25094
rect 18432 24954 18460 26318
rect 18524 25702 18552 28902
rect 18616 26217 18644 31198
rect 18694 30832 18750 30841
rect 18694 30767 18750 30776
rect 18708 30734 18736 30767
rect 18696 30728 18748 30734
rect 18696 30670 18748 30676
rect 18708 30297 18736 30670
rect 18800 30326 18828 31622
rect 18892 31498 18920 32370
rect 18984 31754 19012 32914
rect 19076 31822 19104 37080
rect 19156 37062 19208 37068
rect 19444 36378 19472 37130
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19892 36576 19944 36582
rect 19892 36518 19944 36524
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19904 36174 19932 36518
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 19340 36100 19392 36106
rect 19340 36042 19392 36048
rect 19352 35086 19380 36042
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35086 20024 37878
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 20076 37120 20128 37126
rect 20076 37062 20128 37068
rect 19340 35080 19392 35086
rect 19432 35080 19484 35086
rect 19340 35022 19392 35028
rect 19430 35048 19432 35057
rect 19984 35080 20036 35086
rect 19484 35048 19486 35057
rect 19984 35022 20036 35028
rect 19430 34983 19486 34992
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19430 34776 19486 34785
rect 19574 34779 19882 34788
rect 19430 34711 19432 34720
rect 19484 34711 19486 34720
rect 19432 34682 19484 34688
rect 19800 34672 19852 34678
rect 19800 34614 19852 34620
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19340 33924 19392 33930
rect 19340 33866 19392 33872
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 18972 31748 19024 31754
rect 18972 31690 19024 31696
rect 18892 31470 19104 31498
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 18788 30320 18840 30326
rect 18694 30288 18750 30297
rect 18788 30262 18840 30268
rect 18694 30223 18750 30232
rect 18708 26994 18736 30223
rect 18788 30184 18840 30190
rect 18788 30126 18840 30132
rect 18800 29714 18828 30126
rect 18892 30025 18920 31350
rect 18970 30968 19026 30977
rect 18970 30903 19026 30912
rect 18984 30870 19012 30903
rect 18972 30864 19024 30870
rect 18972 30806 19024 30812
rect 18970 30424 19026 30433
rect 18970 30359 18972 30368
rect 19024 30359 19026 30368
rect 18972 30330 19024 30336
rect 18878 30016 18934 30025
rect 18878 29951 18934 29960
rect 18788 29708 18840 29714
rect 18788 29650 18840 29656
rect 19076 29458 19104 31470
rect 19168 31346 19196 32370
rect 19156 31340 19208 31346
rect 19156 31282 19208 31288
rect 19168 30841 19196 31282
rect 19352 31142 19380 33866
rect 19444 33454 19472 34546
rect 19812 33998 19840 34614
rect 19996 34542 20024 34886
rect 19984 34536 20036 34542
rect 19984 34478 20036 34484
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19616 33448 19668 33454
rect 19616 33390 19668 33396
rect 19628 33289 19656 33390
rect 19614 33280 19670 33289
rect 19614 33215 19670 33224
rect 19432 32836 19484 32842
rect 19432 32778 19484 32784
rect 19340 31136 19392 31142
rect 19340 31078 19392 31084
rect 19154 30832 19210 30841
rect 19154 30767 19210 30776
rect 19340 30728 19392 30734
rect 19260 30676 19340 30682
rect 19260 30670 19392 30676
rect 19260 30654 19380 30670
rect 19156 30116 19208 30122
rect 19260 30104 19288 30654
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19208 30076 19288 30104
rect 19156 30058 19208 30064
rect 19154 30016 19210 30025
rect 19154 29951 19210 29960
rect 19168 29646 19196 29951
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 19248 29572 19300 29578
rect 19248 29514 19300 29520
rect 18800 29430 19196 29458
rect 18800 29306 18828 29430
rect 18878 29336 18934 29345
rect 18788 29300 18840 29306
rect 18878 29271 18934 29280
rect 19064 29300 19116 29306
rect 18788 29242 18840 29248
rect 18892 29084 18920 29271
rect 19064 29242 19116 29248
rect 19076 29209 19104 29242
rect 19062 29200 19118 29209
rect 19062 29135 19118 29144
rect 19064 29096 19116 29102
rect 18786 29064 18842 29073
rect 18892 29056 19064 29084
rect 19064 29038 19116 29044
rect 18786 28999 18842 29008
rect 18800 28218 18828 28999
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 19064 27056 19116 27062
rect 18984 27016 19064 27044
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 18800 26450 18828 26930
rect 18984 26858 19012 27016
rect 19064 26998 19116 27004
rect 18880 26852 18932 26858
rect 18880 26794 18932 26800
rect 18972 26852 19024 26858
rect 18972 26794 19024 26800
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 18892 26314 18920 26794
rect 18880 26308 18932 26314
rect 18880 26250 18932 26256
rect 18602 26208 18658 26217
rect 18602 26143 18658 26152
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18328 24676 18380 24682
rect 18328 24618 18380 24624
rect 18340 24410 18368 24618
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 18432 24290 18460 24754
rect 18340 24262 18460 24290
rect 18340 23866 18368 24262
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18340 22642 18368 23802
rect 18432 23730 18460 24006
rect 18524 23866 18552 25638
rect 18616 25362 18644 25638
rect 18604 25356 18656 25362
rect 18604 25298 18656 25304
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18708 24750 18736 25230
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 19076 24682 19104 26794
rect 19168 25226 19196 29430
rect 19260 29238 19288 29514
rect 19352 29510 19380 30534
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19248 29232 19300 29238
rect 19248 29174 19300 29180
rect 19444 28694 19472 32778
rect 19904 32774 19932 33458
rect 20088 32858 20116 37062
rect 20180 36786 20208 37810
rect 21008 37806 21036 38372
rect 22560 38344 22612 38350
rect 22558 38312 22560 38321
rect 22612 38312 22614 38321
rect 22558 38247 22614 38256
rect 22284 38208 22336 38214
rect 22284 38150 22336 38156
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 22008 37868 22060 37874
rect 22008 37810 22060 37816
rect 20904 37800 20956 37806
rect 20904 37742 20956 37748
rect 20996 37800 21048 37806
rect 20996 37742 21048 37748
rect 20168 36780 20220 36786
rect 20168 36722 20220 36728
rect 20180 34746 20208 36722
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20352 36576 20404 36582
rect 20352 36518 20404 36524
rect 20364 36174 20392 36518
rect 20456 36174 20484 36654
rect 20916 36582 20944 37742
rect 21548 37732 21600 37738
rect 21548 37674 21600 37680
rect 21560 37262 21588 37674
rect 21548 37256 21600 37262
rect 21548 37198 21600 37204
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21456 36848 21508 36854
rect 21456 36790 21508 36796
rect 20904 36576 20956 36582
rect 20904 36518 20956 36524
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20444 36168 20496 36174
rect 20720 36168 20772 36174
rect 20444 36110 20496 36116
rect 20548 36128 20720 36156
rect 20352 36032 20404 36038
rect 20352 35974 20404 35980
rect 20168 34740 20220 34746
rect 20168 34682 20220 34688
rect 20180 34202 20208 34682
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 20168 33108 20220 33114
rect 20168 33050 20220 33056
rect 19996 32830 20116 32858
rect 19892 32768 19944 32774
rect 19892 32710 19944 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19524 32428 19576 32434
rect 19524 32370 19576 32376
rect 19536 31754 19564 32370
rect 19892 32224 19944 32230
rect 19892 32166 19944 32172
rect 19536 31726 19840 31754
rect 19812 31686 19840 31726
rect 19800 31680 19852 31686
rect 19904 31668 19932 32166
rect 19996 31906 20024 32830
rect 20076 32768 20128 32774
rect 20076 32710 20128 32716
rect 20088 32434 20116 32710
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 20180 32366 20208 33050
rect 20168 32360 20220 32366
rect 20168 32302 20220 32308
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 19996 31878 20116 31906
rect 19984 31816 20036 31822
rect 19982 31784 19984 31793
rect 20036 31784 20038 31793
rect 19982 31719 20038 31728
rect 19904 31640 20024 31668
rect 19800 31622 19852 31628
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19892 31340 19944 31346
rect 19892 31282 19944 31288
rect 19904 30938 19932 31282
rect 19892 30932 19944 30938
rect 19892 30874 19944 30880
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19892 30252 19944 30258
rect 19892 30194 19944 30200
rect 19708 30116 19760 30122
rect 19708 30058 19760 30064
rect 19720 29850 19748 30058
rect 19800 30048 19852 30054
rect 19904 30025 19932 30194
rect 19800 29990 19852 29996
rect 19890 30016 19946 30025
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 19616 29708 19668 29714
rect 19616 29650 19668 29656
rect 19628 29510 19656 29650
rect 19812 29617 19840 29990
rect 19890 29951 19946 29960
rect 19996 29646 20024 31640
rect 20088 31124 20116 31878
rect 20180 31385 20208 32166
rect 20166 31376 20222 31385
rect 20166 31311 20222 31320
rect 20272 31278 20300 34546
rect 20364 34524 20392 35974
rect 20548 34678 20576 36128
rect 20720 36110 20772 36116
rect 20904 35760 20956 35766
rect 20904 35702 20956 35708
rect 20916 35222 20944 35702
rect 20720 35216 20772 35222
rect 20720 35158 20772 35164
rect 20904 35216 20956 35222
rect 20904 35158 20956 35164
rect 20732 34950 20760 35158
rect 21468 35086 21496 36790
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20996 35080 21048 35086
rect 21456 35080 21508 35086
rect 20996 35022 21048 35028
rect 21270 35048 21326 35057
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20444 34672 20496 34678
rect 20442 34640 20444 34649
rect 20536 34672 20588 34678
rect 20496 34640 20498 34649
rect 20536 34614 20588 34620
rect 20628 34672 20680 34678
rect 20628 34614 20680 34620
rect 20442 34575 20498 34584
rect 20364 34496 20576 34524
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 20364 32026 20392 34342
rect 20442 34232 20498 34241
rect 20442 34167 20498 34176
rect 20456 33998 20484 34167
rect 20444 33992 20496 33998
rect 20444 33934 20496 33940
rect 20548 33930 20576 34496
rect 20536 33924 20588 33930
rect 20536 33866 20588 33872
rect 20536 33516 20588 33522
rect 20536 33458 20588 33464
rect 20444 33040 20496 33046
rect 20444 32982 20496 32988
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20364 31890 20392 31962
rect 20352 31884 20404 31890
rect 20352 31826 20404 31832
rect 20352 31680 20404 31686
rect 20456 31657 20484 32982
rect 20548 31890 20576 33458
rect 20640 32910 20668 34614
rect 20628 32904 20680 32910
rect 20628 32846 20680 32852
rect 20628 32768 20680 32774
rect 20628 32710 20680 32716
rect 20640 31958 20668 32710
rect 20732 32502 20760 34886
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20824 34241 20852 34546
rect 20810 34232 20866 34241
rect 20810 34167 20866 34176
rect 20720 32496 20772 32502
rect 20720 32438 20772 32444
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20732 31958 20760 32234
rect 20916 32201 20944 35022
rect 21008 34746 21036 35022
rect 21180 35012 21232 35018
rect 21456 35022 21508 35028
rect 21270 34983 21272 34992
rect 21180 34954 21232 34960
rect 21324 34983 21326 34992
rect 21272 34954 21324 34960
rect 20996 34740 21048 34746
rect 20996 34682 21048 34688
rect 21192 34066 21220 34954
rect 21180 34060 21232 34066
rect 21180 34002 21232 34008
rect 21088 33584 21140 33590
rect 21088 33526 21140 33532
rect 20996 32904 21048 32910
rect 20996 32846 21048 32852
rect 20902 32192 20958 32201
rect 20902 32127 20958 32136
rect 20916 31958 20944 32127
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 20904 31952 20956 31958
rect 20904 31894 20956 31900
rect 20536 31884 20588 31890
rect 20536 31826 20588 31832
rect 20352 31622 20404 31628
rect 20442 31648 20498 31657
rect 20260 31272 20312 31278
rect 20260 31214 20312 31220
rect 20088 31096 20300 31124
rect 20076 30320 20128 30326
rect 20076 30262 20128 30268
rect 20088 29850 20116 30262
rect 20272 30258 20300 31096
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20180 29850 20208 30194
rect 20364 30054 20392 31622
rect 20442 31583 20498 31592
rect 20352 30048 20404 30054
rect 20352 29990 20404 29996
rect 20364 29850 20392 29990
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 20168 29844 20220 29850
rect 20168 29786 20220 29792
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 19984 29640 20036 29646
rect 19798 29608 19854 29617
rect 19984 29582 20036 29588
rect 19798 29543 19854 29552
rect 19616 29504 19668 29510
rect 19996 29481 20024 29582
rect 19616 29446 19668 29452
rect 19982 29472 20038 29481
rect 19574 29404 19882 29413
rect 19982 29407 20038 29416
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 20088 28966 20116 29786
rect 20166 29744 20222 29753
rect 20166 29679 20168 29688
rect 20220 29679 20222 29688
rect 20168 29650 20220 29656
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20076 28960 20128 28966
rect 20076 28902 20128 28908
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 20272 28558 20300 29582
rect 20364 28626 20392 29786
rect 20456 28994 20484 31583
rect 20536 31408 20588 31414
rect 20536 31350 20588 31356
rect 20548 31113 20576 31350
rect 20640 31278 20668 31894
rect 20812 31884 20864 31890
rect 20812 31826 20864 31832
rect 20824 31482 20852 31826
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20628 31272 20680 31278
rect 20628 31214 20680 31220
rect 20628 31136 20680 31142
rect 20534 31104 20590 31113
rect 20628 31078 20680 31084
rect 20534 31039 20590 31048
rect 20640 30326 20668 31078
rect 20732 30977 20760 31282
rect 20718 30968 20774 30977
rect 20718 30903 20774 30912
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20548 29832 20576 30262
rect 20640 30002 20668 30262
rect 20732 30258 20760 30903
rect 20824 30870 20852 31418
rect 20916 31346 20944 31894
rect 21008 31754 21036 32846
rect 20996 31748 21048 31754
rect 20996 31690 21048 31696
rect 20904 31340 20956 31346
rect 20904 31282 20956 31288
rect 21008 31142 21036 31690
rect 20996 31136 21048 31142
rect 20996 31078 21048 31084
rect 20812 30864 20864 30870
rect 20812 30806 20864 30812
rect 21100 30326 21128 33526
rect 21468 33522 21496 35022
rect 21560 34649 21588 37198
rect 21640 36032 21692 36038
rect 21640 35974 21692 35980
rect 21652 35766 21680 35974
rect 21640 35760 21692 35766
rect 21640 35702 21692 35708
rect 21836 35698 21864 37198
rect 21928 36854 21956 37198
rect 21916 36848 21968 36854
rect 21916 36790 21968 36796
rect 21928 36582 21956 36790
rect 21916 36576 21968 36582
rect 21916 36518 21968 36524
rect 21916 35760 21968 35766
rect 21916 35702 21968 35708
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21546 34640 21602 34649
rect 21546 34575 21602 34584
rect 21652 34542 21680 35022
rect 21744 34678 21772 35634
rect 21824 35488 21876 35494
rect 21824 35430 21876 35436
rect 21732 34672 21784 34678
rect 21732 34614 21784 34620
rect 21640 34536 21692 34542
rect 21836 34524 21864 35430
rect 21640 34478 21692 34484
rect 21744 34496 21864 34524
rect 21548 33856 21600 33862
rect 21548 33798 21600 33804
rect 21456 33516 21508 33522
rect 21456 33458 21508 33464
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21180 32768 21232 32774
rect 21180 32710 21232 32716
rect 21192 31890 21220 32710
rect 21180 31884 21232 31890
rect 21180 31826 21232 31832
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 21272 31680 21324 31686
rect 21272 31622 21324 31628
rect 21192 30870 21220 31622
rect 21180 30864 21232 30870
rect 21180 30806 21232 30812
rect 21284 30734 21312 31622
rect 21376 31521 21404 33254
rect 21456 32768 21508 32774
rect 21456 32710 21508 32716
rect 21468 31958 21496 32710
rect 21456 31952 21508 31958
rect 21456 31894 21508 31900
rect 21362 31512 21418 31521
rect 21362 31447 21418 31456
rect 21560 31464 21588 33798
rect 21652 31686 21680 34478
rect 21744 33998 21772 34496
rect 21824 34400 21876 34406
rect 21824 34342 21876 34348
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21732 33380 21784 33386
rect 21732 33322 21784 33328
rect 21744 32366 21772 33322
rect 21836 33289 21864 34342
rect 21928 33862 21956 35702
rect 21916 33856 21968 33862
rect 21916 33798 21968 33804
rect 22020 33590 22048 37810
rect 22100 37664 22152 37670
rect 22100 37606 22152 37612
rect 22112 37262 22140 37606
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22100 36236 22152 36242
rect 22100 36178 22152 36184
rect 22112 36145 22140 36178
rect 22098 36136 22154 36145
rect 22098 36071 22154 36080
rect 22204 35816 22232 37946
rect 22296 37942 22324 38150
rect 22664 38010 22692 38490
rect 24400 38412 24452 38418
rect 24400 38354 24452 38360
rect 22652 38004 22704 38010
rect 22652 37946 22704 37952
rect 23940 38004 23992 38010
rect 23940 37946 23992 37952
rect 22284 37936 22336 37942
rect 22284 37878 22336 37884
rect 22296 36122 22324 37878
rect 22468 37868 22520 37874
rect 22468 37810 22520 37816
rect 22652 37868 22704 37874
rect 22652 37810 22704 37816
rect 22836 37868 22888 37874
rect 22836 37810 22888 37816
rect 22928 37868 22980 37874
rect 22980 37828 23060 37856
rect 22928 37810 22980 37816
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 22388 37262 22416 37606
rect 22376 37256 22428 37262
rect 22376 37198 22428 37204
rect 22480 36378 22508 37810
rect 22664 37262 22692 37810
rect 22848 37738 22876 37810
rect 22836 37732 22888 37738
rect 22836 37674 22888 37680
rect 22652 37256 22704 37262
rect 22652 37198 22704 37204
rect 22664 36922 22692 37198
rect 22836 37188 22888 37194
rect 22836 37130 22888 37136
rect 22928 37188 22980 37194
rect 22928 37130 22980 37136
rect 22652 36916 22704 36922
rect 22652 36858 22704 36864
rect 22468 36372 22520 36378
rect 22468 36314 22520 36320
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22468 36168 22520 36174
rect 22296 36094 22416 36122
rect 22468 36110 22520 36116
rect 22112 35788 22232 35816
rect 22112 33590 22140 35788
rect 22388 35698 22416 36094
rect 22192 35692 22244 35698
rect 22376 35692 22428 35698
rect 22192 35634 22244 35640
rect 22296 35652 22376 35680
rect 22204 35601 22232 35634
rect 22190 35592 22246 35601
rect 22190 35527 22246 35536
rect 22190 35456 22246 35465
rect 22190 35391 22246 35400
rect 22204 35290 22232 35391
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 22296 35086 22324 35652
rect 22376 35634 22428 35640
rect 22376 35488 22428 35494
rect 22480 35476 22508 36110
rect 22560 35692 22612 35698
rect 22664 35680 22692 36178
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22756 35834 22784 36110
rect 22848 36009 22876 37130
rect 22940 36650 22968 37130
rect 22928 36644 22980 36650
rect 22928 36586 22980 36592
rect 22834 36000 22890 36009
rect 22834 35935 22890 35944
rect 22744 35828 22796 35834
rect 22744 35770 22796 35776
rect 22836 35692 22888 35698
rect 22664 35652 22836 35680
rect 22560 35634 22612 35640
rect 22836 35634 22888 35640
rect 22428 35448 22508 35476
rect 22376 35430 22428 35436
rect 22284 35080 22336 35086
rect 22204 35040 22284 35068
rect 22204 34610 22232 35040
rect 22284 35022 22336 35028
rect 22284 34944 22336 34950
rect 22284 34886 22336 34892
rect 22296 34610 22324 34886
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22388 34490 22416 35430
rect 22204 34462 22416 34490
rect 22466 34504 22522 34513
rect 22008 33584 22060 33590
rect 22008 33526 22060 33532
rect 22100 33584 22152 33590
rect 22100 33526 22152 33532
rect 21822 33280 21878 33289
rect 21822 33215 21878 33224
rect 21916 33040 21968 33046
rect 21916 32982 21968 32988
rect 21824 32768 21876 32774
rect 21824 32710 21876 32716
rect 21836 32570 21864 32710
rect 21824 32564 21876 32570
rect 21824 32506 21876 32512
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21732 32224 21784 32230
rect 21732 32166 21784 32172
rect 21640 31680 21692 31686
rect 21638 31648 21640 31657
rect 21692 31648 21694 31657
rect 21638 31583 21694 31592
rect 21376 30734 21404 31447
rect 21560 31436 21680 31464
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 21456 31136 21508 31142
rect 21456 31078 21508 31084
rect 21468 30870 21496 31078
rect 21456 30864 21508 30870
rect 21456 30806 21508 30812
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21468 30326 21496 30670
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 21088 30320 21140 30326
rect 21088 30262 21140 30268
rect 21272 30320 21324 30326
rect 21272 30262 21324 30268
rect 21456 30320 21508 30326
rect 21456 30262 21508 30268
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20718 30152 20774 30161
rect 20824 30138 20852 30262
rect 20774 30110 20852 30138
rect 20718 30087 20774 30096
rect 20640 29974 20852 30002
rect 20720 29844 20772 29850
rect 20548 29804 20720 29832
rect 20720 29786 20772 29792
rect 20824 29714 20852 29974
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20548 29578 20760 29594
rect 20536 29572 20760 29578
rect 20588 29566 20760 29572
rect 20536 29514 20588 29520
rect 20732 29170 20760 29566
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20456 28966 20576 28994
rect 20352 28620 20404 28626
rect 20352 28562 20404 28568
rect 20548 28558 20576 28966
rect 20628 28960 20680 28966
rect 20628 28902 20680 28908
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 20260 28552 20312 28558
rect 20260 28494 20312 28500
rect 20536 28552 20588 28558
rect 20536 28494 20588 28500
rect 19352 27878 19380 28494
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 27946 20024 28358
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 19800 27940 19852 27946
rect 19800 27882 19852 27888
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 19444 27577 19472 27882
rect 19524 27872 19576 27878
rect 19522 27840 19524 27849
rect 19576 27840 19578 27849
rect 19522 27775 19578 27784
rect 19812 27674 19840 27882
rect 20088 27674 20116 28018
rect 19800 27668 19852 27674
rect 19800 27610 19852 27616
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 19430 27568 19486 27577
rect 19430 27503 19486 27512
rect 19444 27470 19472 27503
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 19536 27316 19564 27406
rect 19984 27396 20036 27402
rect 19984 27338 20036 27344
rect 19444 27288 19564 27316
rect 19340 26784 19392 26790
rect 19340 26726 19392 26732
rect 19352 26586 19380 26726
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19338 26480 19394 26489
rect 19338 26415 19394 26424
rect 19156 25220 19208 25226
rect 19156 25162 19208 25168
rect 19064 24676 19116 24682
rect 19064 24618 19116 24624
rect 18604 24336 18656 24342
rect 18604 24278 18656 24284
rect 18616 24041 18644 24278
rect 19076 24274 19104 24618
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 18602 24032 18658 24041
rect 18602 23967 18658 23976
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18510 23760 18566 23769
rect 18420 23724 18472 23730
rect 18510 23695 18512 23704
rect 18420 23666 18472 23672
rect 18564 23695 18566 23704
rect 18604 23724 18656 23730
rect 18512 23666 18564 23672
rect 18604 23666 18656 23672
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18340 20534 18368 20878
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18432 20058 18460 23666
rect 18616 23322 18644 23666
rect 18972 23520 19024 23526
rect 18972 23462 19024 23468
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18880 23180 18932 23186
rect 18708 23140 18880 23168
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18524 22794 18552 23054
rect 18616 22982 18644 23054
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18708 22794 18736 23140
rect 18880 23122 18932 23128
rect 18984 23050 19012 23462
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 18880 22976 18932 22982
rect 18932 22924 19012 22930
rect 18880 22918 19012 22924
rect 18892 22902 19012 22918
rect 18524 22766 18736 22794
rect 18984 22642 19012 22902
rect 19076 22642 19104 23054
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18604 20868 18656 20874
rect 18604 20810 18656 20816
rect 18616 20534 18644 20810
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18432 19666 18460 19722
rect 18432 19638 18552 19666
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18340 17202 18368 18634
rect 18524 18290 18552 19638
rect 18616 19310 18644 20470
rect 18708 20398 18736 22102
rect 18892 21622 18920 22510
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 18880 21412 18932 21418
rect 18880 21354 18932 21360
rect 18892 21078 18920 21354
rect 18880 21072 18932 21078
rect 18880 21014 18932 21020
rect 18892 20942 18920 21014
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18708 19854 18736 20334
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18708 18426 18736 19314
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18432 17678 18460 18158
rect 18524 17882 18552 18226
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18420 17536 18472 17542
rect 18418 17504 18420 17513
rect 18472 17504 18474 17513
rect 18418 17439 18474 17448
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17866 15600 17922 15609
rect 17866 15535 17922 15544
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17776 15428 17828 15434
rect 17696 15388 17776 15416
rect 17776 15370 17828 15376
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17696 13938 17724 14418
rect 17788 13938 17816 15370
rect 17958 15056 18014 15065
rect 17868 15020 17920 15026
rect 18064 15042 18092 15438
rect 18014 15026 18092 15042
rect 18014 15020 18104 15026
rect 18014 15014 18052 15020
rect 17958 14991 18014 15000
rect 17868 14962 17920 14968
rect 18052 14962 18104 14968
rect 17880 14414 17908 14962
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17972 14074 18000 14282
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17866 13968 17922 13977
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17776 13932 17828 13938
rect 17866 13903 17922 13912
rect 17776 13874 17828 13880
rect 17512 12406 17632 12434
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16224 11898 16252 12106
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10470 17356 11086
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 10266 17356 10406
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 8430 16160 9862
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15488 5370 15516 5578
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15120 5234 15240 5250
rect 15108 5228 15240 5234
rect 15160 5222 15240 5228
rect 15108 5170 15160 5176
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 15304 4486 15332 5306
rect 15580 4826 15608 5850
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16408 5234 16436 5510
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 11794 4040 11850 4049
rect 11794 3975 11850 3984
rect 13174 4040 13230 4049
rect 13174 3975 13230 3984
rect 11808 3058 11836 3975
rect 13188 3058 13216 3975
rect 16500 3194 16528 8842
rect 16684 8634 16712 10066
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 9110 17264 9318
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17512 8974 17540 12406
rect 17696 11830 17724 13874
rect 17788 12782 17816 13874
rect 17880 13802 17908 13903
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 18156 12986 18184 16730
rect 18248 15162 18276 17070
rect 18326 15192 18382 15201
rect 18236 15156 18288 15162
rect 18326 15127 18382 15136
rect 18236 15098 18288 15104
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18248 14278 18276 14894
rect 18340 14822 18368 15127
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 18156 12238 18184 12922
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17696 11150 17724 11766
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17604 10742 17632 11018
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 10130 17908 10406
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17972 10062 18000 11494
rect 18248 11150 18276 14214
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18340 13530 18368 13874
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18064 10674 18092 11086
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18248 9926 18276 9998
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18142 9752 18198 9761
rect 18142 9687 18198 9696
rect 17866 9616 17922 9625
rect 17866 9551 17922 9560
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7410 17632 7822
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17052 6934 17080 7346
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 7002 17264 7142
rect 17420 7002 17448 7346
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17604 6798 17632 6870
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16592 5302 16620 6666
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 17696 3194 17724 9114
rect 17880 9042 17908 9551
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17972 8974 18000 9454
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 8974 18092 9318
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18156 7886 18184 9687
rect 18340 8906 18368 12786
rect 18432 10470 18460 17206
rect 18524 16658 18552 17682
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18524 11150 18552 14282
rect 18616 13938 18644 18226
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18708 17338 18736 17750
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18800 16590 18828 18022
rect 18892 17338 18920 20878
rect 18984 20806 19012 22578
rect 19076 22098 19104 22578
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19076 20942 19104 21490
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 19076 20534 19104 20878
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18984 20058 19012 20198
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 19076 19378 19104 19654
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18984 19174 19012 19246
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18984 18290 19012 19110
rect 19076 18698 19104 19314
rect 19064 18692 19116 18698
rect 19064 18634 19116 18640
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18970 18184 19026 18193
rect 18970 18119 19026 18128
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18892 16454 18920 17070
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 16250 18920 16390
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18984 16114 19012 18119
rect 19076 18086 19104 18634
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18616 12918 18644 13874
rect 18708 13394 18736 15846
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18800 14482 18828 14962
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18786 14104 18842 14113
rect 18786 14039 18788 14048
rect 18840 14039 18842 14048
rect 18788 14010 18840 14016
rect 18788 13864 18840 13870
rect 18892 13852 18920 15506
rect 18984 15502 19012 16050
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 19076 14482 19104 16526
rect 19168 14618 19196 25162
rect 19352 24138 19380 26415
rect 19444 24886 19472 27288
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19706 25800 19762 25809
rect 19996 25770 20024 27338
rect 20088 26314 20116 27406
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 19706 25735 19708 25744
rect 19760 25735 19762 25744
rect 19984 25764 20036 25770
rect 19708 25706 19760 25712
rect 19984 25706 20036 25712
rect 19706 25528 19762 25537
rect 19706 25463 19762 25472
rect 19720 25294 19748 25463
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19432 24880 19484 24886
rect 19432 24822 19484 24828
rect 19996 24410 20024 25094
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 23526 19288 24006
rect 19444 23798 19472 24142
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19260 22642 19288 23462
rect 19892 23044 19944 23050
rect 19996 23032 20024 24142
rect 20088 23050 20116 26250
rect 20180 25498 20208 28018
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 20180 24818 20208 25434
rect 20272 25378 20300 28494
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 20364 28150 20392 28426
rect 20548 28218 20576 28494
rect 20536 28212 20588 28218
rect 20536 28154 20588 28160
rect 20352 28144 20404 28150
rect 20640 28098 20668 28902
rect 20720 28756 20772 28762
rect 20720 28698 20772 28704
rect 20732 28150 20760 28698
rect 21100 28218 21128 30262
rect 21284 30138 21312 30262
rect 21284 30110 21404 30138
rect 21272 30048 21324 30054
rect 21272 29990 21324 29996
rect 21284 29889 21312 29990
rect 21270 29880 21326 29889
rect 21270 29815 21326 29824
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21088 28212 21140 28218
rect 21088 28154 21140 28160
rect 20352 28086 20404 28092
rect 20456 28070 20668 28098
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20456 27470 20484 28070
rect 20628 27668 20680 27674
rect 20628 27610 20680 27616
rect 20444 27464 20496 27470
rect 20444 27406 20496 27412
rect 20534 27432 20590 27441
rect 20534 27367 20590 27376
rect 20548 26489 20576 27367
rect 20534 26480 20590 26489
rect 20534 26415 20590 26424
rect 20536 26308 20588 26314
rect 20536 26250 20588 26256
rect 20352 25968 20404 25974
rect 20352 25910 20404 25916
rect 20364 25498 20392 25910
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20352 25492 20404 25498
rect 20352 25434 20404 25440
rect 20272 25350 20392 25378
rect 20456 25362 20484 25638
rect 20258 25120 20314 25129
rect 20258 25055 20314 25064
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20272 24342 20300 25055
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 19944 23004 20024 23032
rect 20076 23044 20128 23050
rect 19892 22986 19944 22992
rect 20076 22986 20128 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19260 18766 19288 19790
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 18193 19288 18226
rect 19246 18184 19302 18193
rect 19246 18119 19302 18128
rect 19352 18034 19380 22374
rect 20180 22094 20208 24006
rect 20364 23798 20392 25350
rect 20444 25356 20496 25362
rect 20444 25298 20496 25304
rect 20548 24993 20576 26250
rect 20640 25906 20668 27610
rect 20732 27130 20760 28086
rect 20996 27872 21048 27878
rect 20996 27814 21048 27820
rect 21008 27713 21036 27814
rect 20994 27704 21050 27713
rect 20994 27639 21050 27648
rect 20810 27568 20866 27577
rect 20810 27503 20866 27512
rect 20824 27470 20852 27503
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 21008 27062 21036 27338
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 20902 26480 20958 26489
rect 20902 26415 20958 26424
rect 20916 26382 20944 26415
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20812 26240 20864 26246
rect 20810 26208 20812 26217
rect 20864 26208 20866 26217
rect 20810 26143 20866 26152
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20628 25764 20680 25770
rect 20628 25706 20680 25712
rect 20640 25158 20668 25706
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20732 25294 20760 25434
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20534 24984 20590 24993
rect 20534 24919 20590 24928
rect 20442 24848 20498 24857
rect 20548 24818 20576 24919
rect 20628 24880 20680 24886
rect 20628 24822 20680 24828
rect 20732 24834 20760 25230
rect 20824 24954 20852 25638
rect 20812 24948 20864 24954
rect 20812 24890 20864 24896
rect 20442 24783 20498 24792
rect 20536 24812 20588 24818
rect 20456 24206 20484 24783
rect 20536 24754 20588 24760
rect 20548 24274 20576 24754
rect 20640 24585 20668 24822
rect 20732 24806 20852 24834
rect 20916 24818 20944 26318
rect 20626 24576 20682 24585
rect 20626 24511 20682 24520
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20626 24168 20682 24177
rect 20626 24103 20682 24112
rect 20640 24070 20668 24103
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20640 23746 20668 24006
rect 20718 23760 20774 23769
rect 20536 23724 20588 23730
rect 20640 23718 20718 23746
rect 20824 23730 20852 24806
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 21008 24750 21036 26998
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 21100 24614 21128 27406
rect 21192 26382 21220 29446
rect 21284 29034 21312 29815
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21284 27674 21312 28018
rect 21272 27668 21324 27674
rect 21272 27610 21324 27616
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21192 25537 21220 25842
rect 21178 25528 21234 25537
rect 21178 25463 21234 25472
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20718 23695 20774 23704
rect 20812 23724 20864 23730
rect 20536 23666 20588 23672
rect 20812 23666 20864 23672
rect 20442 23216 20498 23225
rect 20442 23151 20498 23160
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20272 22098 20300 22986
rect 20456 22642 20484 23151
rect 20548 23050 20576 23666
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20548 22506 20576 22986
rect 20640 22642 20668 23258
rect 20916 23225 20944 24006
rect 21008 23633 21036 24346
rect 20994 23624 21050 23633
rect 20994 23559 21050 23568
rect 20902 23216 20958 23225
rect 20902 23151 20958 23160
rect 20720 23112 20772 23118
rect 21008 23100 21036 23559
rect 21086 23488 21142 23497
rect 21192 23474 21220 25463
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21284 24410 21312 24754
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21376 24154 21404 30110
rect 21454 30016 21510 30025
rect 21454 29951 21510 29960
rect 21468 28014 21496 29951
rect 21560 29170 21588 31282
rect 21652 30054 21680 31436
rect 21744 30802 21772 32166
rect 21928 31736 21956 32982
rect 22008 32904 22060 32910
rect 22008 32846 22060 32852
rect 22020 32434 22048 32846
rect 22112 32609 22140 33526
rect 22204 32910 22232 34462
rect 22466 34439 22468 34448
rect 22520 34439 22522 34448
rect 22468 34410 22520 34416
rect 22468 34196 22520 34202
rect 22468 34138 22520 34144
rect 22376 33992 22428 33998
rect 22376 33934 22428 33940
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 22098 32600 22154 32609
rect 22204 32570 22232 32846
rect 22098 32535 22154 32544
rect 22192 32564 22244 32570
rect 22192 32506 22244 32512
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 21836 31708 21956 31736
rect 21732 30796 21784 30802
rect 21732 30738 21784 30744
rect 21836 30734 21864 31708
rect 21914 31648 21970 31657
rect 22020 31634 22048 31826
rect 22112 31804 22140 32370
rect 22296 32298 22324 33050
rect 22388 32842 22416 33934
rect 22376 32836 22428 32842
rect 22376 32778 22428 32784
rect 22388 32745 22416 32778
rect 22374 32736 22430 32745
rect 22374 32671 22430 32680
rect 22376 32564 22428 32570
rect 22376 32506 22428 32512
rect 22284 32292 22336 32298
rect 22284 32234 22336 32240
rect 22192 31816 22244 31822
rect 22112 31784 22192 31804
rect 22244 31784 22246 31793
rect 22112 31776 22190 31784
rect 22190 31719 22246 31728
rect 22020 31606 22140 31634
rect 21914 31583 21970 31592
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 21836 30394 21864 30670
rect 21824 30388 21876 30394
rect 21824 30330 21876 30336
rect 21640 30048 21692 30054
rect 21640 29990 21692 29996
rect 21548 29164 21600 29170
rect 21548 29106 21600 29112
rect 21456 28008 21508 28014
rect 21456 27950 21508 27956
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 21468 27538 21496 27814
rect 21456 27532 21508 27538
rect 21456 27474 21508 27480
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21468 25906 21496 26386
rect 21560 26314 21588 29106
rect 21652 27878 21680 29990
rect 21822 29880 21878 29889
rect 21822 29815 21878 29824
rect 21836 29782 21864 29815
rect 21824 29776 21876 29782
rect 21824 29718 21876 29724
rect 21928 29306 21956 31583
rect 22008 31476 22060 31482
rect 22008 31418 22060 31424
rect 22020 29782 22048 31418
rect 22112 31414 22140 31606
rect 22388 31498 22416 32506
rect 22480 31686 22508 34138
rect 22572 32026 22600 35634
rect 22652 35488 22704 35494
rect 22652 35430 22704 35436
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22664 35290 22692 35430
rect 22652 35284 22704 35290
rect 22652 35226 22704 35232
rect 22756 34406 22784 35430
rect 22940 35018 22968 36586
rect 23032 35737 23060 37828
rect 23112 37664 23164 37670
rect 23112 37606 23164 37612
rect 23124 37466 23152 37606
rect 23112 37460 23164 37466
rect 23112 37402 23164 37408
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23018 35728 23074 35737
rect 23018 35663 23074 35672
rect 22928 35012 22980 35018
rect 22928 34954 22980 34960
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22848 34746 22876 34886
rect 22926 34776 22982 34785
rect 22836 34740 22888 34746
rect 22926 34711 22982 34720
rect 22836 34682 22888 34688
rect 22940 34542 22968 34711
rect 22928 34536 22980 34542
rect 22928 34478 22980 34484
rect 22744 34400 22796 34406
rect 22744 34342 22796 34348
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 22664 32910 22692 33798
rect 22744 33584 22796 33590
rect 22744 33526 22796 33532
rect 22756 33046 22784 33526
rect 22836 33312 22888 33318
rect 22836 33254 22888 33260
rect 22744 33040 22796 33046
rect 22744 32982 22796 32988
rect 22848 32910 22876 33254
rect 23032 32994 23060 35663
rect 23124 35562 23152 37198
rect 23572 37188 23624 37194
rect 23572 37130 23624 37136
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 23112 35556 23164 35562
rect 23112 35498 23164 35504
rect 23110 35456 23166 35465
rect 23110 35391 23166 35400
rect 23124 35086 23152 35391
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23216 34950 23244 37062
rect 23584 36378 23612 37130
rect 23664 37120 23716 37126
rect 23664 37062 23716 37068
rect 23296 36372 23348 36378
rect 23296 36314 23348 36320
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23112 34944 23164 34950
rect 23112 34886 23164 34892
rect 23204 34944 23256 34950
rect 23204 34886 23256 34892
rect 23124 34524 23152 34886
rect 23204 34536 23256 34542
rect 23124 34496 23204 34524
rect 23204 34478 23256 34484
rect 23204 34400 23256 34406
rect 23204 34342 23256 34348
rect 23110 33144 23166 33153
rect 23110 33079 23166 33088
rect 22940 32966 23060 32994
rect 22652 32904 22704 32910
rect 22652 32846 22704 32852
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22744 32768 22796 32774
rect 22744 32710 22796 32716
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 22664 32473 22692 32506
rect 22650 32464 22706 32473
rect 22756 32434 22784 32710
rect 22940 32434 22968 32966
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 23032 32570 23060 32846
rect 23124 32774 23152 33079
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 23020 32564 23072 32570
rect 23020 32506 23072 32512
rect 23112 32496 23164 32502
rect 23112 32438 23164 32444
rect 22650 32399 22706 32408
rect 22744 32428 22796 32434
rect 22744 32370 22796 32376
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 22652 32360 22704 32366
rect 22652 32302 22704 32308
rect 23020 32360 23072 32366
rect 23020 32302 23072 32308
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22560 31816 22612 31822
rect 22560 31758 22612 31764
rect 22468 31680 22520 31686
rect 22468 31622 22520 31628
rect 22388 31470 22508 31498
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 22388 30598 22416 30670
rect 22376 30592 22428 30598
rect 22376 30534 22428 30540
rect 22480 30410 22508 31470
rect 22204 30382 22508 30410
rect 22008 29776 22060 29782
rect 22060 29736 22140 29764
rect 22008 29718 22060 29724
rect 22112 29617 22140 29736
rect 22098 29608 22154 29617
rect 22008 29572 22060 29578
rect 22098 29543 22154 29552
rect 22008 29514 22060 29520
rect 22020 29306 22048 29514
rect 21916 29300 21968 29306
rect 21916 29242 21968 29248
rect 22008 29300 22060 29306
rect 22008 29242 22060 29248
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22020 28490 22048 29106
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 22008 28484 22060 28490
rect 22008 28426 22060 28432
rect 22112 28218 22140 28970
rect 22008 28212 22060 28218
rect 22008 28154 22060 28160
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 21824 28144 21876 28150
rect 21824 28086 21876 28092
rect 21732 28008 21784 28014
rect 21732 27950 21784 27956
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21548 26308 21600 26314
rect 21548 26250 21600 26256
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21548 25220 21600 25226
rect 21548 25162 21600 25168
rect 21376 24126 21496 24154
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21284 23594 21312 24006
rect 21376 23798 21404 24006
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21468 23730 21496 24126
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21272 23588 21324 23594
rect 21272 23530 21324 23536
rect 21192 23446 21312 23474
rect 21086 23423 21142 23432
rect 20720 23054 20772 23060
rect 20916 23072 21036 23100
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20364 22234 20392 22374
rect 20548 22273 20576 22442
rect 20534 22264 20590 22273
rect 20352 22228 20404 22234
rect 20534 22199 20590 22208
rect 20352 22170 20404 22176
rect 19996 22066 20208 22094
rect 20260 22092 20312 22098
rect 20640 22094 20668 22578
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21672 19472 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21690 20024 22066
rect 20260 22034 20312 22040
rect 20456 22066 20668 22094
rect 19984 21684 20036 21690
rect 19444 21644 19564 21672
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19444 21010 19472 21422
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19432 20868 19484 20874
rect 19536 20856 19564 21644
rect 19984 21626 20036 21632
rect 19708 21412 19760 21418
rect 19708 21354 19760 21360
rect 20168 21412 20220 21418
rect 20168 21354 20220 21360
rect 19484 20828 19564 20856
rect 19432 20810 19484 20816
rect 19720 20806 19748 21354
rect 20180 21010 20208 21354
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19444 19378 19472 19858
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19378 20024 20266
rect 20088 19990 20116 20402
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19444 18970 19472 19314
rect 20088 19258 20116 19926
rect 20180 19922 20208 20742
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20166 19544 20222 19553
rect 20166 19479 20222 19488
rect 20180 19446 20208 19479
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 20272 19394 20300 20402
rect 20364 20058 20392 20402
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20272 19366 20392 19394
rect 20260 19304 20312 19310
rect 19996 19230 20208 19258
rect 20260 19246 20312 19252
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19904 18737 19932 19110
rect 19890 18728 19946 18737
rect 19890 18663 19946 18672
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 19260 18006 19380 18034
rect 19260 17524 19288 18006
rect 19720 17921 19748 18294
rect 19798 18184 19854 18193
rect 19798 18119 19854 18128
rect 19338 17912 19394 17921
rect 19338 17847 19394 17856
rect 19706 17912 19762 17921
rect 19706 17847 19762 17856
rect 19352 17678 19380 17847
rect 19812 17746 19840 18119
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19616 17536 19668 17542
rect 19260 17496 19380 17524
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18840 13824 18920 13852
rect 18972 13864 19024 13870
rect 18788 13806 18840 13812
rect 18972 13806 19024 13812
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18708 12102 18736 13330
rect 18800 12306 18828 13806
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18524 10674 18552 11086
rect 18984 11014 19012 13806
rect 19076 12850 19104 14418
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19260 14074 19288 14282
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19352 12442 19380 17496
rect 19444 17496 19616 17524
rect 19444 16590 19472 17496
rect 19904 17524 19932 17682
rect 19904 17496 19948 17524
rect 19616 17478 19668 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19920 17338 19948 17496
rect 19892 17332 19948 17338
rect 19944 17292 19948 17332
rect 19892 17274 19944 17280
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19798 17096 19854 17105
rect 19904 17082 19932 17138
rect 19996 17082 20024 19230
rect 20180 18970 20208 19230
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20272 18816 20300 19246
rect 20180 18788 20300 18816
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 20088 18290 20116 18634
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 20088 17678 20116 18226
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20088 17202 20116 17614
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 19904 17066 20116 17082
rect 19798 17031 19854 17040
rect 19892 17060 20116 17066
rect 19616 16720 19668 16726
rect 19616 16662 19668 16668
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19628 16522 19656 16662
rect 19812 16590 19840 17031
rect 19944 17054 20116 17060
rect 19892 17002 19944 17008
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15094 20024 16526
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19628 14618 19656 14758
rect 20088 14618 20116 17054
rect 20180 15162 20208 18788
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20272 17746 20300 18226
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20272 17338 20300 17546
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20364 17218 20392 19366
rect 20456 17377 20484 22066
rect 20732 21622 20760 23054
rect 20916 22642 20944 23072
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20824 22234 20852 22374
rect 21008 22234 21036 22918
rect 21100 22778 21128 23423
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21192 22642 21220 23122
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21178 22536 21234 22545
rect 21178 22471 21180 22480
rect 21232 22471 21234 22480
rect 21180 22442 21232 22448
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 21284 22030 21312 23446
rect 21362 23352 21418 23361
rect 21362 23287 21418 23296
rect 21376 23254 21404 23287
rect 21364 23248 21416 23254
rect 21364 23190 21416 23196
rect 21468 22778 21496 23666
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20732 20942 20760 21422
rect 20824 20942 20852 21422
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21100 20942 21128 21354
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20732 20466 20760 20878
rect 20824 20466 20852 20878
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20548 18834 20576 19654
rect 20640 18970 20668 19654
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20548 17678 20576 18770
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20442 17368 20498 17377
rect 20442 17303 20498 17312
rect 20272 17190 20392 17218
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20180 14414 20208 14826
rect 20272 14822 20300 17190
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20364 16726 20392 17002
rect 20456 16794 20484 17002
rect 20548 16794 20576 17614
rect 20640 17338 20668 18566
rect 20732 18426 20760 20402
rect 21100 20262 21128 20878
rect 21284 20466 21312 21558
rect 21376 21486 21404 22374
rect 21468 22030 21496 22510
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21468 21894 21496 21966
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21376 20924 21404 21422
rect 21456 20936 21508 20942
rect 21376 20896 21456 20924
rect 21456 20878 21508 20884
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21468 20058 21496 20878
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21560 19334 21588 25162
rect 21652 24138 21680 27814
rect 21744 25498 21772 27950
rect 21836 27470 21864 28086
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 21824 26784 21876 26790
rect 21824 26726 21876 26732
rect 21732 25492 21784 25498
rect 21732 25434 21784 25440
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21652 23322 21680 23462
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21640 23180 21692 23186
rect 21744 23168 21772 23666
rect 21836 23662 21864 26726
rect 22020 24274 22048 28154
rect 22112 27441 22140 28154
rect 22204 27470 22232 30382
rect 22468 29572 22520 29578
rect 22468 29514 22520 29520
rect 22480 29306 22508 29514
rect 22572 29306 22600 31758
rect 22664 30122 22692 32302
rect 23032 32201 23060 32302
rect 23018 32192 23074 32201
rect 23018 32127 23074 32136
rect 22742 32056 22798 32065
rect 22742 31991 22798 32000
rect 22756 31822 22784 31991
rect 22744 31816 22796 31822
rect 22744 31758 22796 31764
rect 23124 31754 23152 32438
rect 22848 31726 23152 31754
rect 22848 30734 22876 31726
rect 23020 31680 23072 31686
rect 23020 31622 23072 31628
rect 23112 31680 23164 31686
rect 23216 31668 23244 34342
rect 23308 33590 23336 36314
rect 23572 35624 23624 35630
rect 23572 35566 23624 35572
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 23400 35222 23428 35430
rect 23388 35216 23440 35222
rect 23388 35158 23440 35164
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23400 34950 23428 35022
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23478 34640 23534 34649
rect 23584 34610 23612 35566
rect 23478 34575 23480 34584
rect 23532 34575 23534 34584
rect 23572 34604 23624 34610
rect 23480 34546 23532 34552
rect 23572 34546 23624 34552
rect 23388 34536 23440 34542
rect 23388 34478 23440 34484
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 23400 33454 23428 34478
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 23296 32836 23348 32842
rect 23296 32778 23348 32784
rect 23164 31640 23244 31668
rect 23112 31622 23164 31628
rect 22928 31476 22980 31482
rect 22928 31418 22980 31424
rect 22940 31346 22968 31418
rect 23032 31346 23060 31622
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 23020 31340 23072 31346
rect 23020 31282 23072 31288
rect 22940 31142 22968 31282
rect 23124 31226 23152 31622
rect 23308 31482 23336 32778
rect 23400 32502 23428 33390
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 23492 32502 23520 32710
rect 23388 32496 23440 32502
rect 23388 32438 23440 32444
rect 23480 32496 23532 32502
rect 23480 32438 23532 32444
rect 23388 32360 23440 32366
rect 23388 32302 23440 32308
rect 23400 31929 23428 32302
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23572 32224 23624 32230
rect 23572 32166 23624 32172
rect 23386 31920 23442 31929
rect 23386 31855 23442 31864
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 23032 31198 23152 31226
rect 22928 31136 22980 31142
rect 22928 31078 22980 31084
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22652 30116 22704 30122
rect 22652 30058 22704 30064
rect 22468 29300 22520 29306
rect 22468 29242 22520 29248
rect 22560 29300 22612 29306
rect 22560 29242 22612 29248
rect 22664 29170 22692 30058
rect 22284 29164 22336 29170
rect 22284 29106 22336 29112
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22296 28393 22324 29106
rect 22282 28384 22338 28393
rect 22282 28319 22338 28328
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22192 27464 22244 27470
rect 22098 27432 22154 27441
rect 22192 27406 22244 27412
rect 22098 27367 22154 27376
rect 22296 26790 22324 28018
rect 22388 27946 22416 29106
rect 22376 27940 22428 27946
rect 22376 27882 22428 27888
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22204 25906 22232 26522
rect 22480 26518 22508 29106
rect 22572 28150 22600 29106
rect 22652 28960 22704 28966
rect 22652 28902 22704 28908
rect 22664 28422 22692 28902
rect 22756 28529 22784 30330
rect 22848 30025 22876 30670
rect 22928 30592 22980 30598
rect 22928 30534 22980 30540
rect 22940 30433 22968 30534
rect 22926 30424 22982 30433
rect 22926 30359 22982 30368
rect 22928 30048 22980 30054
rect 22834 30016 22890 30025
rect 22928 29990 22980 29996
rect 22834 29951 22890 29960
rect 22940 29646 22968 29990
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22848 29306 22876 29446
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22940 29186 22968 29582
rect 22848 29158 22968 29186
rect 22742 28520 22798 28529
rect 22742 28455 22798 28464
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22756 28218 22784 28455
rect 22744 28212 22796 28218
rect 22744 28154 22796 28160
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22650 28112 22706 28121
rect 22650 28047 22706 28056
rect 22558 27976 22614 27985
rect 22664 27946 22692 28047
rect 22558 27911 22614 27920
rect 22652 27940 22704 27946
rect 22572 27470 22600 27911
rect 22652 27882 22704 27888
rect 22560 27464 22612 27470
rect 22560 27406 22612 27412
rect 22468 26512 22520 26518
rect 22468 26454 22520 26460
rect 22560 26240 22612 26246
rect 22560 26182 22612 26188
rect 22572 25906 22600 26182
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22468 25764 22520 25770
rect 22468 25706 22520 25712
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 22204 25294 22232 25638
rect 22284 25424 22336 25430
rect 22284 25366 22336 25372
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22296 24993 22324 25366
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 22388 25129 22416 25230
rect 22374 25120 22430 25129
rect 22374 25055 22430 25064
rect 22282 24984 22338 24993
rect 22282 24919 22338 24928
rect 22100 24812 22152 24818
rect 22284 24812 22336 24818
rect 22100 24754 22152 24760
rect 22204 24772 22284 24800
rect 22112 24410 22140 24754
rect 22204 24721 22232 24772
rect 22284 24754 22336 24760
rect 22190 24712 22246 24721
rect 22190 24647 22246 24656
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22204 24313 22232 24550
rect 22190 24304 22246 24313
rect 22008 24268 22060 24274
rect 21928 24228 22008 24256
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 21928 23594 21956 24228
rect 22190 24239 22246 24248
rect 22008 24210 22060 24216
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22008 24132 22060 24138
rect 22008 24074 22060 24080
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 21692 23140 21772 23168
rect 21640 23122 21692 23128
rect 21652 22030 21680 23122
rect 21916 23112 21968 23118
rect 21836 23072 21916 23100
rect 21836 23066 21864 23072
rect 21744 23038 21864 23066
rect 21916 23054 21968 23060
rect 21744 22438 21772 23038
rect 21822 22808 21878 22817
rect 21822 22743 21878 22752
rect 21916 22772 21968 22778
rect 21836 22710 21864 22743
rect 21916 22714 21968 22720
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21836 22234 21864 22374
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21928 21078 21956 22714
rect 22020 22545 22048 24074
rect 22112 23866 22140 24142
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22204 23866 22232 24006
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 22204 23746 22232 23802
rect 22112 23718 22232 23746
rect 22112 23118 22140 23718
rect 22388 23526 22416 25055
rect 22480 24954 22508 25706
rect 22560 25424 22612 25430
rect 22560 25366 22612 25372
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22480 24177 22508 24754
rect 22572 24206 22600 25366
rect 22664 24596 22692 27882
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22756 25974 22784 26454
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22744 25764 22796 25770
rect 22744 25706 22796 25712
rect 22756 25498 22784 25706
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22848 24721 22876 29158
rect 22926 28792 22982 28801
rect 23032 28778 23060 31198
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 23216 30938 23244 31078
rect 23204 30932 23256 30938
rect 23204 30874 23256 30880
rect 23308 30818 23336 31282
rect 23124 30790 23336 30818
rect 23124 30054 23152 30790
rect 23296 30592 23348 30598
rect 23296 30534 23348 30540
rect 23202 30288 23258 30297
rect 23202 30223 23258 30232
rect 23216 30122 23244 30223
rect 23204 30116 23256 30122
rect 23204 30058 23256 30064
rect 23112 30048 23164 30054
rect 23112 29990 23164 29996
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23124 29481 23152 29582
rect 23110 29472 23166 29481
rect 23110 29407 23166 29416
rect 23216 28994 23244 30058
rect 23308 29782 23336 30534
rect 23296 29776 23348 29782
rect 23296 29718 23348 29724
rect 22982 28750 23060 28778
rect 23124 28966 23244 28994
rect 22926 28727 22982 28736
rect 22940 28472 22968 28727
rect 23020 28484 23072 28490
rect 22940 28444 23020 28472
rect 23020 28426 23072 28432
rect 22926 28384 22982 28393
rect 22926 28319 22982 28328
rect 22940 28218 22968 28319
rect 22928 28212 22980 28218
rect 22928 28154 22980 28160
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22940 27946 22968 28018
rect 22928 27940 22980 27946
rect 22928 27882 22980 27888
rect 23032 27334 23060 28426
rect 23124 28082 23152 28966
rect 23400 28626 23428 31758
rect 23492 30938 23520 32166
rect 23480 30932 23532 30938
rect 23480 30874 23532 30880
rect 23584 30580 23612 32166
rect 23676 30734 23704 37062
rect 23860 36922 23888 37198
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23756 34944 23808 34950
rect 23756 34886 23808 34892
rect 23768 33522 23796 34886
rect 23756 33516 23808 33522
rect 23756 33458 23808 33464
rect 23768 32366 23796 33458
rect 23848 33108 23900 33114
rect 23848 33050 23900 33056
rect 23860 32910 23888 33050
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23848 32428 23900 32434
rect 23952 32416 23980 37946
rect 24412 36922 24440 38354
rect 24780 38214 24808 38898
rect 24952 38752 25004 38758
rect 24952 38694 25004 38700
rect 24964 38418 24992 38694
rect 25056 38554 25084 38898
rect 26148 38888 26200 38894
rect 26148 38830 26200 38836
rect 25044 38548 25096 38554
rect 25044 38490 25096 38496
rect 25042 38448 25098 38457
rect 24952 38412 25004 38418
rect 26160 38418 26188 38830
rect 27080 38729 27108 38898
rect 31208 38752 31260 38758
rect 27066 38720 27122 38729
rect 27066 38655 27122 38664
rect 31206 38720 31208 38729
rect 31260 38720 31262 38729
rect 31206 38655 31262 38664
rect 33060 38554 33088 38898
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35636 38554 35664 38898
rect 37922 38856 37978 38865
rect 37922 38791 37978 38800
rect 37936 38554 37964 38791
rect 27896 38548 27948 38554
rect 27896 38490 27948 38496
rect 30288 38548 30340 38554
rect 30288 38490 30340 38496
rect 33048 38548 33100 38554
rect 33048 38490 33100 38496
rect 35624 38548 35676 38554
rect 35624 38490 35676 38496
rect 37924 38548 37976 38554
rect 37924 38490 37976 38496
rect 27540 38418 27660 38434
rect 25042 38383 25098 38392
rect 26148 38412 26200 38418
rect 24952 38354 25004 38360
rect 24860 38276 24912 38282
rect 24860 38218 24912 38224
rect 24952 38276 25004 38282
rect 24952 38218 25004 38224
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 24676 37324 24728 37330
rect 24676 37266 24728 37272
rect 24400 36916 24452 36922
rect 24400 36858 24452 36864
rect 24582 36816 24638 36825
rect 24582 36751 24638 36760
rect 24596 36650 24624 36751
rect 24584 36644 24636 36650
rect 24584 36586 24636 36592
rect 24124 36168 24176 36174
rect 24124 36110 24176 36116
rect 24032 35556 24084 35562
rect 24032 35498 24084 35504
rect 24044 32842 24072 35498
rect 24032 32836 24084 32842
rect 24032 32778 24084 32784
rect 24136 32434 24164 36110
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24216 35148 24268 35154
rect 24216 35090 24268 35096
rect 23900 32388 23980 32416
rect 24124 32428 24176 32434
rect 23848 32370 23900 32376
rect 24124 32370 24176 32376
rect 23756 32360 23808 32366
rect 23860 32337 23888 32370
rect 23756 32302 23808 32308
rect 23846 32328 23902 32337
rect 23846 32263 23902 32272
rect 23940 32292 23992 32298
rect 23940 32234 23992 32240
rect 23848 32224 23900 32230
rect 23754 32192 23810 32201
rect 23848 32166 23900 32172
rect 23754 32127 23810 32136
rect 23768 32026 23796 32127
rect 23756 32020 23808 32026
rect 23756 31962 23808 31968
rect 23860 31754 23888 32166
rect 23952 32065 23980 32234
rect 23938 32056 23994 32065
rect 23938 31991 23994 32000
rect 23768 31726 23888 31754
rect 23768 30734 23796 31726
rect 23848 31272 23900 31278
rect 23848 31214 23900 31220
rect 23664 30728 23716 30734
rect 23664 30670 23716 30676
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23664 30592 23716 30598
rect 23584 30552 23664 30580
rect 23716 30552 23796 30580
rect 23664 30534 23716 30540
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23676 29170 23704 29446
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23664 29164 23716 29170
rect 23664 29106 23716 29112
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23388 28620 23440 28626
rect 23388 28562 23440 28568
rect 23296 28484 23348 28490
rect 23296 28426 23348 28432
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23124 27146 23152 28018
rect 23216 27470 23244 28358
rect 23308 28082 23336 28426
rect 23296 28076 23348 28082
rect 23296 28018 23348 28024
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 23308 27538 23336 27814
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23400 27402 23428 28018
rect 23388 27396 23440 27402
rect 23388 27338 23440 27344
rect 23032 27118 23152 27146
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 22940 25158 22968 25298
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 22834 24712 22890 24721
rect 22834 24647 22890 24656
rect 22664 24568 22876 24596
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22560 24200 22612 24206
rect 22466 24168 22522 24177
rect 22560 24142 22612 24148
rect 22466 24103 22522 24112
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22006 22536 22062 22545
rect 22006 22471 22062 22480
rect 22020 21418 22048 22471
rect 22112 22030 22140 22918
rect 22204 22166 22232 23122
rect 22388 22982 22416 23122
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22480 22642 22508 24103
rect 22664 23730 22692 24346
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22756 24070 22784 24142
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 22652 23724 22704 23730
rect 22572 23684 22652 23712
rect 22572 23118 22600 23684
rect 22652 23666 22704 23672
rect 22650 23624 22706 23633
rect 22650 23559 22706 23568
rect 22664 23526 22692 23559
rect 22652 23520 22704 23526
rect 22652 23462 22704 23468
rect 22664 23186 22692 23462
rect 22652 23180 22704 23186
rect 22652 23122 22704 23128
rect 22756 23118 22784 23734
rect 22848 23202 22876 24568
rect 22940 23322 22968 25094
rect 23032 23594 23060 27118
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 23204 26036 23256 26042
rect 23204 25978 23256 25984
rect 23216 25945 23244 25978
rect 23202 25936 23258 25945
rect 23112 25900 23164 25906
rect 23308 25906 23336 26318
rect 23202 25871 23258 25880
rect 23296 25900 23348 25906
rect 23112 25842 23164 25848
rect 23296 25842 23348 25848
rect 23124 25362 23152 25842
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 23112 25356 23164 25362
rect 23112 25298 23164 25304
rect 23308 25294 23336 25706
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23110 24848 23166 24857
rect 23308 24834 23336 25230
rect 23166 24806 23336 24834
rect 23110 24783 23166 24792
rect 23400 24342 23428 27338
rect 23492 26042 23520 28902
rect 23584 28150 23612 29106
rect 23768 28994 23796 30552
rect 23860 29646 23888 31214
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 23952 30734 23980 30874
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23860 29306 23888 29582
rect 23848 29300 23900 29306
rect 23848 29242 23900 29248
rect 24044 29170 24072 31078
rect 24032 29164 24084 29170
rect 24032 29106 24084 29112
rect 23676 28966 23796 28994
rect 23572 28144 23624 28150
rect 23572 28086 23624 28092
rect 23584 27577 23612 28086
rect 23570 27568 23626 27577
rect 23570 27503 23626 27512
rect 23676 27470 23704 28966
rect 23754 28656 23810 28665
rect 23810 28614 23980 28642
rect 23754 28591 23810 28600
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 23768 27538 23796 27814
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23480 26036 23532 26042
rect 23480 25978 23532 25984
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23124 23798 23152 24142
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23400 23866 23428 24006
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23020 23588 23072 23594
rect 23020 23530 23072 23536
rect 23112 23588 23164 23594
rect 23112 23530 23164 23536
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 22848 23174 22968 23202
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22192 22160 22244 22166
rect 22192 22102 22244 22108
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22112 21690 22140 21966
rect 22204 21894 22232 22102
rect 22296 22030 22324 22374
rect 22388 22166 22416 22510
rect 22466 22400 22522 22409
rect 22466 22335 22522 22344
rect 22376 22160 22428 22166
rect 22376 22102 22428 22108
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22204 21554 22232 21830
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22296 21486 22324 21966
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22388 21554 22416 21898
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22008 21412 22060 21418
rect 22008 21354 22060 21360
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 21916 21072 21968 21078
rect 21916 21014 21968 21020
rect 22296 20466 22324 21286
rect 22388 21010 22416 21286
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22190 19952 22246 19961
rect 22190 19887 22246 19896
rect 22204 19378 22232 19887
rect 22192 19372 22244 19378
rect 21560 19306 21680 19334
rect 22192 19314 22244 19320
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20824 18290 20852 18702
rect 20916 18358 20944 19178
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20732 17270 20760 17750
rect 20916 17678 20944 18294
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20352 16720 20404 16726
rect 20352 16662 20404 16668
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20444 16584 20496 16590
rect 20442 16552 20444 16561
rect 20496 16552 20498 16561
rect 20442 16487 20498 16496
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20456 15502 20484 16050
rect 20444 15496 20496 15502
rect 20350 15464 20406 15473
rect 20548 15484 20576 16594
rect 20640 16182 20668 17138
rect 20732 16590 20760 17206
rect 21008 17202 21036 17818
rect 21284 17610 21312 18566
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20640 15978 20668 16118
rect 20916 16114 20944 17138
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20916 15502 20944 15642
rect 21008 15570 21036 16730
rect 21100 16574 21128 17070
rect 21192 16998 21220 17138
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 16794 21220 16934
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21180 16584 21232 16590
rect 21100 16546 21180 16574
rect 21180 16526 21232 16532
rect 21284 16522 21312 17546
rect 21376 17338 21404 18634
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21284 15502 21312 16458
rect 20628 15496 20680 15502
rect 20548 15456 20628 15484
rect 20444 15438 20496 15444
rect 20628 15438 20680 15444
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 20350 15399 20406 15408
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19444 12434 19472 13738
rect 20180 13394 20208 14350
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20364 13258 20392 15399
rect 20456 15026 20484 15438
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20456 14414 20484 14962
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 13530 20484 14350
rect 20548 14074 20576 14758
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19444 12406 19564 12434
rect 19444 12170 19472 12406
rect 19536 12374 19564 12406
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19246 11656 19302 11665
rect 19246 11591 19248 11600
rect 19300 11591 19302 11600
rect 19248 11562 19300 11568
rect 19352 11082 19380 12106
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19614 11792 19670 11801
rect 19614 11727 19616 11736
rect 19668 11727 19670 11736
rect 19984 11756 20036 11762
rect 19616 11698 19668 11704
rect 19984 11698 20036 11704
rect 19996 11558 20024 11698
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 18972 11008 19024 11014
rect 18602 10976 18658 10985
rect 18972 10950 19024 10956
rect 18602 10911 18658 10920
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18524 10130 18552 10610
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18616 10062 18644 10911
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18800 10062 18828 10406
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18524 9178 18552 9522
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18340 8566 18368 8842
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 19168 8430 19196 10474
rect 19248 10124 19300 10130
rect 19352 10112 19380 11018
rect 19444 10742 19472 11086
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19300 10084 19380 10112
rect 19248 10066 19300 10072
rect 19352 8956 19380 10084
rect 19892 10056 19944 10062
rect 19890 10024 19892 10033
rect 19944 10024 19946 10033
rect 19890 9959 19946 9968
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19444 9654 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19996 9518 20024 11494
rect 20088 9722 20116 12038
rect 20180 11354 20208 12310
rect 20640 11354 20668 15438
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 15094 20760 15302
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20732 14550 20760 15030
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20916 14482 20944 14962
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20916 13938 20944 14418
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20732 13326 20760 13466
rect 20916 13410 20944 13874
rect 20824 13394 20944 13410
rect 20812 13388 20944 13394
rect 20864 13382 20944 13388
rect 20812 13330 20864 13336
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 12646 20760 13262
rect 20812 12844 20864 12850
rect 20916 12832 20944 13382
rect 21008 13258 21036 14826
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 13938 21128 14758
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21008 12918 21036 13194
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20864 12804 20944 12832
rect 20812 12786 20864 12792
rect 20916 12714 20944 12804
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 21100 12646 21128 13874
rect 21192 13258 21220 14418
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21178 12200 21234 12209
rect 21178 12135 21234 12144
rect 21192 11898 21220 12135
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20260 11280 20312 11286
rect 20260 11222 20312 11228
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20180 10810 20208 10950
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 19984 9512 20036 9518
rect 19798 9480 19854 9489
rect 19984 9454 20036 9460
rect 19798 9415 19800 9424
rect 19852 9415 19854 9424
rect 19800 9386 19852 9392
rect 19524 8968 19576 8974
rect 19352 8928 19524 8956
rect 19524 8910 19576 8916
rect 20180 8838 20208 10746
rect 20272 10538 20300 11222
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20260 10532 20312 10538
rect 20260 10474 20312 10480
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20272 10010 20300 10134
rect 20456 10062 20484 10610
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20444 10056 20496 10062
rect 20272 9982 20392 10010
rect 20444 9998 20496 10004
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19982 8664 20038 8673
rect 19982 8599 19984 8608
rect 20036 8599 20038 8608
rect 20076 8628 20128 8634
rect 19984 8570 20036 8576
rect 20076 8570 20128 8576
rect 20088 8498 20116 8570
rect 20180 8498 20208 8774
rect 20272 8498 20300 9862
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18064 6662 18092 6734
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6458 18092 6598
rect 18432 6458 18460 6802
rect 18616 6798 18644 6938
rect 18694 6896 18750 6905
rect 18694 6831 18750 6840
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18708 6780 18736 6831
rect 18788 6792 18840 6798
rect 18708 6752 18788 6780
rect 18524 6458 18552 6734
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18616 6254 18644 6734
rect 18708 6662 18736 6752
rect 18788 6734 18840 6740
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 19168 6322 19196 8366
rect 19352 7290 19380 8434
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19444 7546 19472 7958
rect 19904 7732 19932 8298
rect 19996 7886 20024 8366
rect 20088 7886 20116 8434
rect 20180 7886 20208 8434
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20364 7750 20392 9982
rect 20548 9518 20576 10542
rect 20640 10130 20668 10746
rect 20916 10674 20944 11222
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20824 10198 20852 10474
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20824 9722 20852 10134
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20916 9586 20944 10610
rect 21088 10192 21140 10198
rect 21086 10160 21088 10169
rect 21140 10160 21142 10169
rect 21086 10095 21142 10104
rect 21086 10024 21142 10033
rect 21086 9959 21142 9968
rect 21100 9654 21128 9959
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20548 9160 20576 9454
rect 20548 9132 20668 9160
rect 20640 9042 20668 9132
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20548 7954 20576 8910
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8498 20668 8774
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20536 7948 20588 7954
rect 20456 7908 20536 7936
rect 20352 7744 20404 7750
rect 19904 7704 20024 7732
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19904 7410 19932 7482
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19352 7262 19472 7290
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 6866 19380 7142
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19352 6458 19380 6802
rect 19444 6458 19472 7262
rect 19904 7002 19932 7346
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 18340 5302 18368 6054
rect 19352 5370 19380 6054
rect 19996 5914 20024 7704
rect 20352 7686 20404 7692
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20180 7206 20208 7346
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20180 7002 20208 7142
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19168 4826 19196 4966
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19260 4622 19288 5238
rect 19352 5234 19380 5306
rect 19996 5302 20024 5850
rect 20088 5710 20116 6938
rect 20272 6934 20300 7346
rect 20352 7268 20404 7274
rect 20352 7210 20404 7216
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20168 5636 20220 5642
rect 20168 5578 20220 5584
rect 20180 5302 20208 5578
rect 19984 5296 20036 5302
rect 19984 5238 20036 5244
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 19352 4690 19380 5170
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19628 4690 19656 4966
rect 20088 4826 20116 5034
rect 20272 4826 20300 5170
rect 20364 5166 20392 7210
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 20088 4486 20116 4762
rect 20364 4554 20392 5102
rect 20456 4690 20484 7908
rect 20536 7890 20588 7896
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20548 7546 20576 7754
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20640 5030 20668 7686
rect 20732 7206 20760 9522
rect 20916 9042 20944 9522
rect 21284 9518 21312 10746
rect 21376 10418 21404 17274
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21560 15706 21588 17070
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21468 11898 21496 12038
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21652 11286 21680 19306
rect 21822 19136 21878 19145
rect 21822 19071 21878 19080
rect 21836 18834 21864 19071
rect 21914 19000 21970 19009
rect 21914 18935 21916 18944
rect 21968 18935 21970 18944
rect 21916 18906 21968 18912
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21836 18426 21864 18770
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21928 18358 21956 18906
rect 22192 18760 22244 18766
rect 22190 18728 22192 18737
rect 22244 18728 22246 18737
rect 22190 18663 22246 18672
rect 21916 18352 21968 18358
rect 21916 18294 21968 18300
rect 22204 18222 22232 18663
rect 22388 18612 22416 20946
rect 22480 18834 22508 22335
rect 22572 22273 22600 22918
rect 22756 22778 22784 23054
rect 22744 22772 22796 22778
rect 22664 22732 22744 22760
rect 22558 22264 22614 22273
rect 22558 22199 22614 22208
rect 22572 19854 22600 22199
rect 22664 21622 22692 22732
rect 22744 22714 22796 22720
rect 22744 22500 22796 22506
rect 22744 22442 22796 22448
rect 22652 21616 22704 21622
rect 22652 21558 22704 21564
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22572 19378 22600 19790
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22652 19304 22704 19310
rect 22650 19272 22652 19281
rect 22704 19272 22706 19281
rect 22650 19207 22706 19216
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22468 18624 22520 18630
rect 22388 18584 22468 18612
rect 22192 18216 22244 18222
rect 22192 18158 22244 18164
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17921 21864 18022
rect 21822 17912 21878 17921
rect 21822 17847 21878 17856
rect 21914 16552 21970 16561
rect 21914 16487 21970 16496
rect 22008 16516 22060 16522
rect 21928 15570 21956 16487
rect 22008 16458 22060 16464
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 22020 14006 22048 16458
rect 22284 15428 22336 15434
rect 22284 15370 22336 15376
rect 22296 14498 22324 15370
rect 22112 14470 22324 14498
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 22112 13462 22140 14470
rect 22192 14340 22244 14346
rect 22192 14282 22244 14288
rect 22204 14074 22232 14282
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22204 13326 22232 14010
rect 22388 13410 22416 18584
rect 22468 18566 22520 18572
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22664 17066 22692 17614
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22572 15706 22600 16458
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22296 13382 22416 13410
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21744 12782 21772 13126
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21836 12730 21864 13126
rect 22296 12968 22324 13382
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22020 12940 22324 12968
rect 21744 12288 21772 12718
rect 21836 12702 21956 12730
rect 21824 12300 21876 12306
rect 21744 12260 21824 12288
rect 21824 12242 21876 12248
rect 21836 12102 21864 12242
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21836 10674 21864 11630
rect 21928 10742 21956 12702
rect 22020 11558 22048 12940
rect 22098 12880 22154 12889
rect 22098 12815 22154 12824
rect 22112 12782 22140 12815
rect 22388 12782 22416 13262
rect 22480 12850 22508 14350
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22572 13530 22600 13806
rect 22664 13716 22692 17002
rect 22756 14278 22784 22442
rect 22940 22094 22968 23174
rect 23124 23118 23152 23530
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23124 22574 23152 23054
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 23204 22094 23256 22098
rect 22940 22092 23256 22094
rect 22940 22066 23204 22092
rect 23492 22094 23520 25638
rect 23584 23730 23612 27270
rect 23756 27124 23808 27130
rect 23756 27066 23808 27072
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23676 22982 23704 25842
rect 23768 24138 23796 27066
rect 23860 26382 23888 28494
rect 23952 28150 23980 28614
rect 23940 28144 23992 28150
rect 23940 28086 23992 28092
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 23848 25832 23900 25838
rect 23848 25774 23900 25780
rect 23860 25362 23888 25774
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23756 24132 23808 24138
rect 23756 24074 23808 24080
rect 23952 23662 23980 28086
rect 24044 26382 24072 29106
rect 24136 28540 24164 32370
rect 24228 31482 24256 35090
rect 24596 34678 24624 35430
rect 24584 34672 24636 34678
rect 24584 34614 24636 34620
rect 24492 34536 24544 34542
rect 24490 34504 24492 34513
rect 24688 34513 24716 37266
rect 24780 34950 24808 37606
rect 24872 37466 24900 38218
rect 24964 38010 24992 38218
rect 24952 38004 25004 38010
rect 24952 37946 25004 37952
rect 24952 37868 25004 37874
rect 25056 37856 25084 38383
rect 26148 38354 26200 38360
rect 27344 38412 27396 38418
rect 27344 38354 27396 38360
rect 27540 38412 27672 38418
rect 27540 38406 27620 38412
rect 27356 38282 27384 38354
rect 27252 38276 27304 38282
rect 27252 38218 27304 38224
rect 27344 38276 27396 38282
rect 27344 38218 27396 38224
rect 26424 38208 26476 38214
rect 26424 38150 26476 38156
rect 26436 38010 26464 38150
rect 27264 38010 27292 38218
rect 26424 38004 26476 38010
rect 26424 37946 26476 37952
rect 27252 38004 27304 38010
rect 27252 37946 27304 37952
rect 25410 37904 25466 37913
rect 25004 37828 25084 37856
rect 25228 37868 25280 37874
rect 24952 37810 25004 37816
rect 25410 37839 25412 37848
rect 25228 37810 25280 37816
rect 25464 37839 25466 37848
rect 25412 37810 25464 37816
rect 25240 37738 25268 37810
rect 25228 37732 25280 37738
rect 25228 37674 25280 37680
rect 24860 37460 24912 37466
rect 24860 37402 24912 37408
rect 25044 37392 25096 37398
rect 25044 37334 25096 37340
rect 24952 36848 25004 36854
rect 24952 36790 25004 36796
rect 24964 36174 24992 36790
rect 25056 36378 25084 37334
rect 25240 37262 25268 37674
rect 25412 37664 25464 37670
rect 25412 37606 25464 37612
rect 26240 37664 26292 37670
rect 26240 37606 26292 37612
rect 25228 37256 25280 37262
rect 25228 37198 25280 37204
rect 25320 36780 25372 36786
rect 25240 36740 25320 36768
rect 25044 36372 25096 36378
rect 25044 36314 25096 36320
rect 24952 36168 25004 36174
rect 24952 36110 25004 36116
rect 25136 36032 25188 36038
rect 25240 36009 25268 36740
rect 25320 36722 25372 36728
rect 25318 36272 25374 36281
rect 25318 36207 25320 36216
rect 25372 36207 25374 36216
rect 25320 36178 25372 36184
rect 25320 36100 25372 36106
rect 25320 36042 25372 36048
rect 25136 35974 25188 35980
rect 25226 36000 25282 36009
rect 25148 35086 25176 35974
rect 25226 35935 25282 35944
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 24768 34944 24820 34950
rect 24768 34886 24820 34892
rect 24544 34504 24546 34513
rect 24490 34439 24546 34448
rect 24674 34504 24730 34513
rect 24674 34439 24730 34448
rect 24308 34060 24360 34066
rect 24584 34060 24636 34066
rect 24360 34020 24584 34048
rect 24308 34002 24360 34008
rect 24584 34002 24636 34008
rect 24320 33658 24348 34002
rect 24676 33924 24728 33930
rect 24676 33866 24728 33872
rect 24308 33652 24360 33658
rect 24308 33594 24360 33600
rect 24308 32836 24360 32842
rect 24308 32778 24360 32784
rect 24216 31476 24268 31482
rect 24216 31418 24268 31424
rect 24228 29714 24256 31418
rect 24320 30122 24348 32778
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24490 32328 24546 32337
rect 24490 32263 24546 32272
rect 24308 30116 24360 30122
rect 24308 30058 24360 30064
rect 24216 29708 24268 29714
rect 24216 29650 24268 29656
rect 24216 29028 24268 29034
rect 24216 28970 24268 28976
rect 24228 28694 24256 28970
rect 24216 28688 24268 28694
rect 24216 28630 24268 28636
rect 24504 28558 24532 32263
rect 24596 31822 24624 32370
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 24688 30122 24716 33866
rect 24780 31754 24808 34886
rect 24872 32298 24900 35022
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 24964 34746 24992 34886
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 24964 33590 24992 34682
rect 25056 34610 25084 34886
rect 25240 34610 25268 35935
rect 25332 35562 25360 36042
rect 25320 35556 25372 35562
rect 25320 35498 25372 35504
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25228 34604 25280 34610
rect 25228 34546 25280 34552
rect 25044 34400 25096 34406
rect 25044 34342 25096 34348
rect 25056 33862 25084 34342
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 25136 33856 25188 33862
rect 25136 33798 25188 33804
rect 24952 33584 25004 33590
rect 24952 33526 25004 33532
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 24860 32292 24912 32298
rect 24860 32234 24912 32240
rect 24964 31890 24992 32370
rect 25056 32366 25084 33798
rect 25044 32360 25096 32366
rect 25044 32302 25096 32308
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 24780 31726 24992 31754
rect 24676 30116 24728 30122
rect 24676 30058 24728 30064
rect 24688 28665 24716 30058
rect 24674 28656 24730 28665
rect 24674 28591 24730 28600
rect 24216 28552 24268 28558
rect 24136 28512 24216 28540
rect 24216 28494 24268 28500
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24124 28076 24176 28082
rect 24124 28018 24176 28024
rect 24136 27470 24164 28018
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 24136 26858 24164 27406
rect 24124 26852 24176 26858
rect 24124 26794 24176 26800
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 24136 25838 24164 26794
rect 24124 25832 24176 25838
rect 24122 25800 24124 25809
rect 24176 25800 24178 25809
rect 24122 25735 24178 25744
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 24044 25498 24072 25638
rect 24032 25492 24084 25498
rect 24032 25434 24084 25440
rect 24228 24818 24256 28494
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24412 27062 24440 27270
rect 24400 27056 24452 27062
rect 24400 26998 24452 27004
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 24398 24440 24454 24449
rect 24398 24375 24400 24384
rect 24452 24375 24454 24384
rect 24400 24346 24452 24352
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24136 23730 24164 24006
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24504 23186 24532 27610
rect 24584 27532 24636 27538
rect 24584 27474 24636 27480
rect 24596 25401 24624 27474
rect 24860 27056 24912 27062
rect 24860 26998 24912 27004
rect 24676 26308 24728 26314
rect 24676 26250 24728 26256
rect 24688 26042 24716 26250
rect 24766 26208 24822 26217
rect 24766 26143 24822 26152
rect 24676 26036 24728 26042
rect 24676 25978 24728 25984
rect 24780 25906 24808 26143
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 24688 25498 24716 25842
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24582 25392 24638 25401
rect 24582 25327 24584 25336
rect 24636 25327 24638 25336
rect 24676 25356 24728 25362
rect 24584 25298 24636 25304
rect 24676 25298 24728 25304
rect 24582 24984 24638 24993
rect 24582 24919 24638 24928
rect 24596 24886 24624 24919
rect 24584 24880 24636 24886
rect 24584 24822 24636 24828
rect 24688 24052 24716 25298
rect 24780 25265 24808 25706
rect 24766 25256 24822 25265
rect 24766 25191 24822 25200
rect 24780 24206 24808 25191
rect 24872 24585 24900 26998
rect 24964 26042 24992 31726
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 25056 27674 25084 30330
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 25148 26194 25176 33798
rect 25240 31754 25268 34546
rect 25332 33980 25360 35498
rect 25424 35222 25452 37606
rect 25872 37120 25924 37126
rect 25872 37062 25924 37068
rect 25688 36576 25740 36582
rect 25688 36518 25740 36524
rect 25780 36576 25832 36582
rect 25780 36518 25832 36524
rect 25504 36168 25556 36174
rect 25700 36156 25728 36518
rect 25556 36128 25728 36156
rect 25504 36110 25556 36116
rect 25596 36032 25648 36038
rect 25502 36000 25558 36009
rect 25558 35980 25596 35986
rect 25558 35974 25648 35980
rect 25558 35958 25636 35974
rect 25502 35935 25558 35944
rect 25596 35760 25648 35766
rect 25596 35702 25648 35708
rect 25502 35592 25558 35601
rect 25502 35527 25504 35536
rect 25556 35527 25558 35536
rect 25504 35498 25556 35504
rect 25608 35222 25636 35702
rect 25700 35680 25728 36128
rect 25792 35834 25820 36518
rect 25780 35828 25832 35834
rect 25780 35770 25832 35776
rect 25780 35692 25832 35698
rect 25700 35652 25780 35680
rect 25780 35634 25832 35640
rect 25412 35216 25464 35222
rect 25412 35158 25464 35164
rect 25596 35216 25648 35222
rect 25596 35158 25648 35164
rect 25424 34785 25452 35158
rect 25780 35080 25832 35086
rect 25780 35022 25832 35028
rect 25596 35012 25648 35018
rect 25596 34954 25648 34960
rect 25410 34776 25466 34785
rect 25410 34711 25466 34720
rect 25504 34468 25556 34474
rect 25504 34410 25556 34416
rect 25516 34241 25544 34410
rect 25608 34406 25636 34954
rect 25792 34746 25820 35022
rect 25780 34740 25832 34746
rect 25780 34682 25832 34688
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25596 34400 25648 34406
rect 25596 34342 25648 34348
rect 25688 34400 25740 34406
rect 25688 34342 25740 34348
rect 25502 34232 25558 34241
rect 25502 34167 25558 34176
rect 25700 33998 25728 34342
rect 25792 34218 25820 34546
rect 25884 34388 25912 37062
rect 25964 36780 26016 36786
rect 25964 36722 26016 36728
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 25976 36174 26004 36722
rect 26056 36304 26108 36310
rect 26054 36272 26056 36281
rect 26108 36272 26110 36281
rect 26054 36207 26110 36216
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 26054 36136 26110 36145
rect 25976 35057 26004 36110
rect 26054 36071 26056 36080
rect 26108 36071 26110 36080
rect 26056 36042 26108 36048
rect 26160 35766 26188 36722
rect 26252 36378 26280 37606
rect 26436 36378 26464 37946
rect 27344 37868 27396 37874
rect 27344 37810 27396 37816
rect 26976 37800 27028 37806
rect 26976 37742 27028 37748
rect 26988 37482 27016 37742
rect 26988 37454 27108 37482
rect 27080 37398 27108 37454
rect 27068 37392 27120 37398
rect 27068 37334 27120 37340
rect 26976 37324 27028 37330
rect 26976 37266 27028 37272
rect 26792 36644 26844 36650
rect 26792 36586 26844 36592
rect 26804 36378 26832 36586
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 26424 36372 26476 36378
rect 26424 36314 26476 36320
rect 26792 36372 26844 36378
rect 26792 36314 26844 36320
rect 26252 36258 26280 36314
rect 26252 36230 26464 36258
rect 26436 36174 26464 36230
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26424 36168 26476 36174
rect 26988 36122 27016 37266
rect 26424 36110 26476 36116
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26148 35760 26200 35766
rect 26148 35702 26200 35708
rect 26252 35698 26280 36042
rect 26056 35692 26108 35698
rect 26056 35634 26108 35640
rect 26240 35692 26292 35698
rect 26240 35634 26292 35640
rect 25962 35048 26018 35057
rect 25962 34983 26018 34992
rect 25976 34610 26004 34983
rect 25964 34604 26016 34610
rect 25964 34546 26016 34552
rect 25884 34360 26004 34388
rect 25792 34190 25912 34218
rect 25412 33992 25464 33998
rect 25332 33952 25412 33980
rect 25412 33934 25464 33940
rect 25688 33992 25740 33998
rect 25688 33934 25740 33940
rect 25424 32910 25452 33934
rect 25688 33516 25740 33522
rect 25688 33458 25740 33464
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25596 32768 25648 32774
rect 25596 32710 25648 32716
rect 25608 32570 25636 32710
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 25700 32434 25728 33458
rect 25780 32904 25832 32910
rect 25780 32846 25832 32852
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25688 32428 25740 32434
rect 25688 32370 25740 32376
rect 25228 31748 25280 31754
rect 25228 31690 25280 31696
rect 25332 31657 25360 32370
rect 25504 32360 25556 32366
rect 25504 32302 25556 32308
rect 25516 31906 25544 32302
rect 25424 31878 25544 31906
rect 25318 31648 25374 31657
rect 25318 31583 25374 31592
rect 25332 31346 25360 31583
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25228 31136 25280 31142
rect 25228 31078 25280 31084
rect 25240 29850 25268 31078
rect 25320 30728 25372 30734
rect 25424 30716 25452 31878
rect 25504 31748 25556 31754
rect 25504 31690 25556 31696
rect 25372 30688 25452 30716
rect 25320 30670 25372 30676
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 25332 29034 25360 30670
rect 25516 30258 25544 31690
rect 25700 31414 25728 32370
rect 25688 31408 25740 31414
rect 25688 31350 25740 31356
rect 25596 31136 25648 31142
rect 25596 31078 25648 31084
rect 25608 30870 25636 31078
rect 25596 30864 25648 30870
rect 25596 30806 25648 30812
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25608 30410 25636 30670
rect 25608 30394 25728 30410
rect 25608 30388 25740 30394
rect 25608 30382 25688 30388
rect 25688 30330 25740 30336
rect 25504 30252 25556 30258
rect 25688 30252 25740 30258
rect 25556 30212 25636 30240
rect 25504 30194 25556 30200
rect 25410 29880 25466 29889
rect 25410 29815 25466 29824
rect 25424 29646 25452 29815
rect 25412 29640 25464 29646
rect 25412 29582 25464 29588
rect 25504 29504 25556 29510
rect 25504 29446 25556 29452
rect 25412 29300 25464 29306
rect 25412 29242 25464 29248
rect 25424 29170 25452 29242
rect 25516 29170 25544 29446
rect 25412 29164 25464 29170
rect 25412 29106 25464 29112
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25228 29028 25280 29034
rect 25228 28970 25280 28976
rect 25320 29028 25372 29034
rect 25320 28970 25372 28976
rect 25056 26166 25176 26194
rect 24952 26036 25004 26042
rect 24952 25978 25004 25984
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24964 25226 24992 25842
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24858 24576 24914 24585
rect 24858 24511 24914 24520
rect 24860 24336 24912 24342
rect 24860 24278 24912 24284
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24768 24064 24820 24070
rect 24688 24024 24768 24052
rect 24768 24006 24820 24012
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24676 23656 24728 23662
rect 24780 23644 24808 24006
rect 24728 23616 24808 23644
rect 24676 23598 24728 23604
rect 24596 23322 24624 23598
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 24400 22976 24452 22982
rect 24400 22918 24452 22924
rect 24412 22166 24440 22918
rect 24400 22160 24452 22166
rect 24400 22102 24452 22108
rect 23492 22066 23612 22094
rect 23204 22034 23256 22040
rect 23110 21992 23166 22001
rect 22836 21956 22888 21962
rect 23110 21927 23166 21936
rect 22836 21898 22888 21904
rect 22848 21554 22876 21898
rect 23018 21720 23074 21729
rect 23018 21655 23074 21664
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22848 18766 22876 21490
rect 23032 21350 23060 21655
rect 23124 21554 23152 21927
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22940 19378 22968 19722
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 23032 19281 23060 20402
rect 23386 20360 23442 20369
rect 23386 20295 23388 20304
rect 23440 20295 23442 20304
rect 23388 20266 23440 20272
rect 23204 20256 23256 20262
rect 23204 20198 23256 20204
rect 23216 20058 23244 20198
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23018 19272 23074 19281
rect 22940 19230 23018 19258
rect 22940 18902 22968 19230
rect 23018 19207 23074 19216
rect 23296 19236 23348 19242
rect 23296 19178 23348 19184
rect 23202 19000 23258 19009
rect 23308 18970 23336 19178
rect 23202 18935 23258 18944
rect 23296 18964 23348 18970
rect 22928 18896 22980 18902
rect 22928 18838 22980 18844
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22848 18057 22876 18702
rect 22834 18048 22890 18057
rect 22834 17983 22890 17992
rect 22940 17785 22968 18702
rect 23032 18329 23060 18770
rect 23124 18714 23152 18838
rect 23216 18834 23244 18935
rect 23296 18906 23348 18912
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23400 18850 23428 18906
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23308 18822 23428 18850
rect 23308 18714 23336 18822
rect 23124 18686 23336 18714
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23018 18320 23074 18329
rect 23018 18255 23074 18264
rect 22926 17776 22982 17785
rect 22926 17711 22982 17720
rect 23032 17134 23060 18255
rect 23110 17912 23166 17921
rect 23110 17847 23166 17856
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23124 16658 23152 17847
rect 23308 17814 23336 18686
rect 23400 18290 23428 18702
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23400 18086 23428 18226
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 23400 17202 23428 18022
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 22926 16552 22982 16561
rect 22926 16487 22982 16496
rect 22940 16454 22968 16487
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 23492 15502 23520 19314
rect 23584 15502 23612 22066
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23768 21146 23796 21830
rect 24676 21616 24728 21622
rect 23938 21584 23994 21593
rect 24676 21558 24728 21564
rect 23938 21519 23994 21528
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23676 18970 23704 20470
rect 23952 20466 23980 21519
rect 24124 21004 24176 21010
rect 24044 20964 24124 20992
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23756 20392 23808 20398
rect 24044 20346 24072 20964
rect 24124 20946 24176 20952
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 24136 20602 24164 20810
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 23756 20334 23808 20340
rect 23768 18970 23796 20334
rect 23860 20318 24072 20346
rect 23860 19378 23888 20318
rect 24228 19990 24256 20742
rect 24216 19984 24268 19990
rect 24216 19926 24268 19932
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23952 19417 23980 19654
rect 23938 19408 23994 19417
rect 23848 19372 23900 19378
rect 23938 19343 23994 19352
rect 23848 19314 23900 19320
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23860 18834 23888 19110
rect 23940 18964 23992 18970
rect 23940 18906 23992 18912
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23860 17746 23888 18294
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23860 17377 23888 17682
rect 23952 17542 23980 18906
rect 24044 18766 24072 19790
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24214 19544 24270 19553
rect 24214 19479 24270 19488
rect 24228 19446 24256 19479
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24412 19378 24440 19654
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24124 19236 24176 19242
rect 24124 19178 24176 19184
rect 24308 19236 24360 19242
rect 24308 19178 24360 19184
rect 24136 18970 24164 19178
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24122 18864 24178 18873
rect 24178 18834 24256 18850
rect 24178 18828 24268 18834
rect 24178 18822 24216 18828
rect 24122 18799 24178 18808
rect 24216 18770 24268 18776
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23846 17368 23902 17377
rect 23846 17303 23902 17312
rect 24136 16998 24164 18702
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24228 17134 24256 17614
rect 24320 17202 24348 19178
rect 24400 18896 24452 18902
rect 24400 18838 24452 18844
rect 24308 17196 24360 17202
rect 24308 17138 24360 17144
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24136 16658 24164 16934
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24306 16552 24362 16561
rect 24306 16487 24362 16496
rect 24320 16114 24348 16487
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24320 15745 24348 16050
rect 24306 15736 24362 15745
rect 24306 15671 24362 15680
rect 23204 15496 23256 15502
rect 23202 15464 23204 15473
rect 23480 15496 23532 15502
rect 23256 15464 23258 15473
rect 23480 15438 23532 15444
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23202 15399 23258 15408
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22744 13728 22796 13734
rect 22664 13688 22744 13716
rect 22744 13670 22796 13676
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21454 10432 21510 10441
rect 21376 10390 21454 10418
rect 21454 10367 21510 10376
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21180 9376 21232 9382
rect 21376 9364 21404 10066
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21232 9336 21404 9364
rect 21180 9318 21232 9324
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20824 8634 20852 8910
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20916 8498 20944 8978
rect 21364 8832 21416 8838
rect 21468 8820 21496 9454
rect 21560 9382 21588 10542
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21652 10130 21680 10406
rect 21914 10160 21970 10169
rect 21640 10124 21692 10130
rect 21914 10095 21970 10104
rect 21640 10066 21692 10072
rect 21928 9994 21956 10095
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21416 8792 21496 8820
rect 21364 8774 21416 8780
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20824 5642 20852 8230
rect 21376 7342 21404 8774
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21192 6798 21220 7210
rect 21652 7002 21680 7414
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21652 6798 21680 6938
rect 21744 6934 21772 7278
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 21928 6798 21956 9318
rect 22112 7528 22140 12718
rect 22296 11694 22324 12718
rect 22388 12306 22416 12718
rect 22480 12442 22508 12786
rect 22756 12714 22784 13670
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22664 12374 22692 12582
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22480 11626 22508 12106
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22468 11620 22520 11626
rect 22468 11562 22520 11568
rect 22572 10674 22600 12038
rect 22664 11762 22692 12310
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22848 11642 22876 13942
rect 23032 13138 23060 14010
rect 23216 13530 23244 15399
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23400 14618 23428 14962
rect 23492 14958 23520 15438
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23480 14952 23532 14958
rect 23480 14894 23532 14900
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23492 14362 23520 14894
rect 23492 14334 23612 14362
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23400 13326 23428 13738
rect 23492 13326 23520 14214
rect 23388 13320 23440 13326
rect 23110 13288 23166 13297
rect 23110 13223 23112 13232
rect 23164 13223 23166 13232
rect 23308 13280 23388 13308
rect 23112 13194 23164 13200
rect 23032 13110 23152 13138
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22928 12096 22980 12102
rect 22926 12064 22928 12073
rect 22980 12064 22982 12073
rect 22926 11999 22982 12008
rect 22664 11614 22876 11642
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22376 10464 22428 10470
rect 22190 10432 22246 10441
rect 22376 10406 22428 10412
rect 22190 10367 22246 10376
rect 22204 10198 22232 10367
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22296 9722 22324 9862
rect 22388 9722 22416 10406
rect 22468 10056 22520 10062
rect 22466 10024 22468 10033
rect 22520 10024 22522 10033
rect 22466 9959 22522 9968
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22466 9344 22522 9353
rect 22466 9279 22522 9288
rect 22480 9178 22508 9279
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22572 8974 22600 10610
rect 22664 10198 22692 11614
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 22652 10192 22704 10198
rect 22652 10134 22704 10140
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22664 8498 22692 10134
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22756 9722 22784 9998
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22848 9586 22876 9862
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22756 9178 22784 9318
rect 22848 9178 22876 9318
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22836 8968 22888 8974
rect 22940 8956 22968 11494
rect 23032 10062 23060 12922
rect 23124 10674 23152 13110
rect 23308 12374 23336 13280
rect 23388 13262 23440 13268
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12986 23428 13126
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23492 12594 23520 13262
rect 23400 12566 23520 12594
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23400 12238 23428 12566
rect 23584 12458 23612 14334
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23676 13734 23704 13874
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23662 13424 23718 13433
rect 23662 13359 23718 13368
rect 23676 13326 23704 13359
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23492 12430 23612 12458
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23216 10062 23244 12174
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23308 10674 23336 11018
rect 23400 10742 23428 11698
rect 23492 11014 23520 12430
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23584 11150 23612 12242
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23584 10810 23612 11086
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 22888 8928 22968 8956
rect 22836 8910 22888 8916
rect 22848 8634 22876 8910
rect 23032 8838 23060 9998
rect 23124 9908 23152 9998
rect 23308 9908 23336 10610
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23492 9926 23520 9998
rect 23124 9880 23336 9908
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23492 9738 23520 9862
rect 23400 9710 23520 9738
rect 23400 9178 23428 9710
rect 23584 9382 23612 10474
rect 23676 10033 23704 13262
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23768 12714 23796 13194
rect 23756 12708 23808 12714
rect 23756 12650 23808 12656
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23768 10062 23796 10406
rect 23756 10056 23808 10062
rect 23662 10024 23718 10033
rect 23756 9998 23808 10004
rect 23662 9959 23718 9968
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22376 7540 22428 7546
rect 22020 7500 22324 7528
rect 22020 7410 22048 7500
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22112 6866 22140 7346
rect 22296 6934 22324 7500
rect 22376 7482 22428 7488
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20456 4146 20484 4626
rect 20640 4146 20668 4966
rect 21284 4826 21312 5170
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21376 4690 21404 6598
rect 21928 6322 21956 6734
rect 22388 6458 22416 7482
rect 22480 7410 22508 7890
rect 22756 7546 22784 8366
rect 23032 8362 23060 8774
rect 23124 8498 23152 8978
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 23216 8362 23244 8570
rect 23308 8566 23336 8978
rect 23584 8634 23612 9318
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23020 8356 23072 8362
rect 23020 8298 23072 8304
rect 23204 8356 23256 8362
rect 23204 8298 23256 8304
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23584 7886 23612 8230
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 23032 7546 23060 7686
rect 23492 7546 23520 7822
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22480 7002 22508 7346
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 22572 6118 22600 6598
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5710 22600 6054
rect 22756 5914 22784 6258
rect 22848 6118 22876 6598
rect 22940 6458 22968 7414
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 23124 6866 23152 7278
rect 23676 7274 23704 9114
rect 23768 8922 23796 9998
rect 23860 9625 23888 10950
rect 23846 9616 23902 9625
rect 23846 9551 23902 9560
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 23860 9194 23888 9386
rect 23952 9382 23980 15302
rect 24320 15162 24348 15671
rect 24412 15638 24440 18838
rect 24504 18358 24532 20878
rect 24688 19854 24716 21558
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24780 19514 24808 23616
rect 24872 23118 24900 24278
rect 24964 24177 24992 24754
rect 24950 24168 25006 24177
rect 24950 24103 25006 24112
rect 24964 24070 24992 24103
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24952 22160 25004 22166
rect 24858 22128 24914 22137
rect 24952 22102 25004 22108
rect 24858 22063 24914 22072
rect 24872 22030 24900 22063
rect 24964 22030 24992 22102
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24964 21350 24992 21966
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 25056 21010 25084 26166
rect 25136 26036 25188 26042
rect 25136 25978 25188 25984
rect 25148 22030 25176 25978
rect 25240 23118 25268 28970
rect 25424 28218 25452 29106
rect 25608 28608 25636 30212
rect 25688 30194 25740 30200
rect 25700 28994 25728 30194
rect 25792 29850 25820 32846
rect 25884 31822 25912 34190
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25870 31512 25926 31521
rect 25870 31447 25926 31456
rect 25884 31414 25912 31447
rect 25872 31408 25924 31414
rect 25872 31350 25924 31356
rect 25872 30796 25924 30802
rect 25872 30738 25924 30744
rect 25884 30433 25912 30738
rect 25870 30424 25926 30433
rect 25870 30359 25926 30368
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25884 29850 25912 29990
rect 25780 29844 25832 29850
rect 25780 29786 25832 29792
rect 25872 29844 25924 29850
rect 25872 29786 25924 29792
rect 25778 29608 25834 29617
rect 25778 29543 25834 29552
rect 25792 29510 25820 29543
rect 25780 29504 25832 29510
rect 25780 29446 25832 29452
rect 25700 28966 25912 28994
rect 25608 28580 25820 28608
rect 25504 28552 25556 28558
rect 25504 28494 25556 28500
rect 25516 28393 25544 28494
rect 25688 28484 25740 28490
rect 25688 28426 25740 28432
rect 25502 28384 25558 28393
rect 25502 28319 25558 28328
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25700 27878 25728 28426
rect 25792 28422 25820 28580
rect 25884 28558 25912 28966
rect 25872 28552 25924 28558
rect 25872 28494 25924 28500
rect 25780 28416 25832 28422
rect 25780 28358 25832 28364
rect 25688 27872 25740 27878
rect 25688 27814 25740 27820
rect 25596 27328 25648 27334
rect 25596 27270 25648 27276
rect 25608 26994 25636 27270
rect 25792 26994 25820 28358
rect 25884 27130 25912 28494
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 25318 26208 25374 26217
rect 25318 26143 25374 26152
rect 25332 25498 25360 26143
rect 25424 26081 25452 26250
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25410 26072 25466 26081
rect 25410 26007 25466 26016
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 25424 25378 25452 26007
rect 25332 25350 25452 25378
rect 25332 23798 25360 25350
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25424 25129 25452 25162
rect 25516 25158 25544 26182
rect 25504 25152 25556 25158
rect 25410 25120 25466 25129
rect 25504 25094 25556 25100
rect 25608 25106 25636 26726
rect 25688 25968 25740 25974
rect 25688 25910 25740 25916
rect 25700 25702 25728 25910
rect 25688 25696 25740 25702
rect 25688 25638 25740 25644
rect 25700 25294 25728 25638
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25686 25120 25742 25129
rect 25410 25055 25466 25064
rect 25516 24818 25544 25094
rect 25608 25078 25686 25106
rect 25686 25055 25742 25064
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25516 24410 25544 24754
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25608 23526 25636 24210
rect 25700 24206 25728 25055
rect 25792 24954 25820 26930
rect 25872 26444 25924 26450
rect 25872 26386 25924 26392
rect 25884 26042 25912 26386
rect 25872 26036 25924 26042
rect 25872 25978 25924 25984
rect 25780 24948 25832 24954
rect 25780 24890 25832 24896
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25778 23624 25834 23633
rect 25778 23559 25834 23568
rect 25596 23520 25648 23526
rect 25596 23462 25648 23468
rect 25320 23180 25372 23186
rect 25320 23122 25372 23128
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25148 21554 25176 21626
rect 25240 21554 25268 23054
rect 25332 21962 25360 23122
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25516 22234 25544 22986
rect 25608 22642 25636 23054
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25608 22094 25636 22578
rect 25516 22066 25636 22094
rect 25516 22030 25544 22066
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 25148 21010 25176 21490
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 25044 21004 25096 21010
rect 25044 20946 25096 20952
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24872 19174 24900 20810
rect 25056 20466 25084 20946
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24952 20324 25004 20330
rect 24952 20266 25004 20272
rect 24964 19854 24992 20266
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24596 17338 24624 17614
rect 24780 17610 24808 18770
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24872 16522 24900 18634
rect 24952 17808 25004 17814
rect 24952 17750 25004 17756
rect 24964 17610 24992 17750
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24964 16114 24992 16662
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24400 15632 24452 15638
rect 24400 15574 24452 15580
rect 24308 15156 24360 15162
rect 24308 15098 24360 15104
rect 24596 15026 24624 16050
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24688 15502 24716 15846
rect 24964 15502 24992 16050
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24136 13870 24164 14894
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24228 13938 24256 14350
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24044 12442 24072 13670
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23860 9166 23980 9194
rect 23952 8974 23980 9166
rect 23940 8968 23992 8974
rect 23768 8906 23888 8922
rect 23940 8910 23992 8916
rect 23768 8900 23900 8906
rect 23768 8894 23848 8900
rect 23768 8498 23796 8894
rect 23848 8842 23900 8848
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23664 7268 23716 7274
rect 23664 7210 23716 7216
rect 23860 6934 23888 8570
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 23952 7002 23980 8230
rect 24044 7886 24072 12378
rect 24136 10062 24164 13806
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 12442 24440 12786
rect 24492 12640 24544 12646
rect 24492 12582 24544 12588
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24320 11762 24348 12174
rect 24504 11830 24532 12582
rect 24596 12238 24624 12854
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24688 11830 24716 15438
rect 25056 14890 25084 18702
rect 25148 18426 25176 19110
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25148 17746 25176 18362
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25148 16810 25176 17682
rect 25240 16946 25268 21286
rect 25332 18426 25360 21490
rect 25424 21457 25452 21966
rect 25410 21448 25466 21457
rect 25410 21383 25466 21392
rect 25412 21004 25464 21010
rect 25412 20946 25464 20952
rect 25424 20913 25452 20946
rect 25410 20904 25466 20913
rect 25410 20839 25466 20848
rect 25410 20496 25466 20505
rect 25516 20466 25544 21966
rect 25688 21956 25740 21962
rect 25688 21898 25740 21904
rect 25594 20632 25650 20641
rect 25594 20567 25650 20576
rect 25410 20431 25412 20440
rect 25464 20431 25466 20440
rect 25504 20460 25556 20466
rect 25412 20402 25464 20408
rect 25504 20402 25556 20408
rect 25608 19854 25636 20567
rect 25700 20466 25728 21898
rect 25792 21554 25820 23559
rect 25976 22030 26004 34360
rect 26068 33998 26096 35634
rect 26238 35456 26294 35465
rect 26344 35442 26372 36110
rect 26516 36100 26568 36106
rect 26516 36042 26568 36048
rect 26804 36094 27016 36122
rect 26528 35494 26556 36042
rect 26294 35414 26372 35442
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 26238 35391 26294 35400
rect 26516 34604 26568 34610
rect 26516 34546 26568 34552
rect 26528 34202 26556 34546
rect 26516 34196 26568 34202
rect 26516 34138 26568 34144
rect 26056 33992 26108 33998
rect 26108 33952 26188 33980
rect 26056 33934 26108 33940
rect 26160 32910 26188 33952
rect 26516 33856 26568 33862
rect 26516 33798 26568 33804
rect 26240 33448 26292 33454
rect 26240 33390 26292 33396
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 26068 32026 26096 32846
rect 26252 32502 26280 33390
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26344 32570 26372 32846
rect 26424 32768 26476 32774
rect 26424 32710 26476 32716
rect 26436 32570 26464 32710
rect 26332 32564 26384 32570
rect 26332 32506 26384 32512
rect 26424 32564 26476 32570
rect 26424 32506 26476 32512
rect 26240 32496 26292 32502
rect 26240 32438 26292 32444
rect 26528 32366 26556 33798
rect 26516 32360 26568 32366
rect 26344 32320 26516 32348
rect 26148 32292 26200 32298
rect 26148 32234 26200 32240
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 26068 30258 26096 31758
rect 26160 31346 26188 32234
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 26252 32026 26280 32166
rect 26240 32020 26292 32026
rect 26240 31962 26292 31968
rect 26344 31754 26372 32320
rect 26516 32302 26568 32308
rect 26608 32360 26660 32366
rect 26608 32302 26660 32308
rect 26620 31754 26648 32302
rect 26344 31726 26464 31754
rect 26620 31726 26740 31754
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 26160 30394 26188 31282
rect 26148 30388 26200 30394
rect 26148 30330 26200 30336
rect 26056 30252 26108 30258
rect 26056 30194 26108 30200
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 26068 29850 26096 29990
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 26054 29744 26110 29753
rect 26160 29730 26188 30330
rect 26332 30184 26384 30190
rect 26332 30126 26384 30132
rect 26344 29850 26372 30126
rect 26332 29844 26384 29850
rect 26332 29786 26384 29792
rect 26110 29702 26188 29730
rect 26054 29679 26110 29688
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 26068 28218 26096 28358
rect 26056 28212 26108 28218
rect 26056 28154 26108 28160
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 26160 27674 26188 28018
rect 26148 27668 26200 27674
rect 26148 27610 26200 27616
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 26068 26353 26096 26930
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26054 26344 26110 26353
rect 26054 26279 26110 26288
rect 26160 25906 26188 26726
rect 26252 26042 26280 28494
rect 26344 27946 26372 28494
rect 26332 27940 26384 27946
rect 26332 27882 26384 27888
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 26148 25492 26200 25498
rect 26148 25434 26200 25440
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 26068 24585 26096 24754
rect 26054 24576 26110 24585
rect 26054 24511 26110 24520
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 25976 21690 26004 21966
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 25962 21584 26018 21593
rect 25780 21548 25832 21554
rect 25962 21519 25964 21528
rect 25780 21490 25832 21496
rect 26016 21519 26018 21528
rect 25964 21490 26016 21496
rect 25792 21321 25820 21490
rect 25778 21312 25834 21321
rect 25778 21247 25834 21256
rect 26056 20868 26108 20874
rect 26056 20810 26108 20816
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25700 19786 25728 20402
rect 25792 20210 25820 20402
rect 25792 20182 25912 20210
rect 25884 19854 25912 20182
rect 25872 19848 25924 19854
rect 25778 19816 25834 19825
rect 25688 19780 25740 19786
rect 25872 19790 25924 19796
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 25778 19751 25780 19760
rect 25688 19722 25740 19728
rect 25832 19751 25834 19760
rect 25780 19722 25832 19728
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25608 18698 25636 19654
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25700 19281 25728 19314
rect 25686 19272 25742 19281
rect 25686 19207 25742 19216
rect 25596 18692 25648 18698
rect 25596 18634 25648 18640
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25332 18193 25360 18362
rect 25318 18184 25374 18193
rect 25318 18119 25374 18128
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 25608 17338 25636 17614
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25700 17134 25728 19207
rect 25778 18864 25834 18873
rect 25778 18799 25834 18808
rect 25792 18766 25820 18799
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25884 18630 25912 19790
rect 25976 19514 26004 19790
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 26068 19378 26096 20810
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 26160 18766 26188 25434
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26252 23866 26280 24006
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 26344 22642 26372 26250
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26332 20868 26384 20874
rect 26332 20810 26384 20816
rect 26344 19378 26372 20810
rect 26436 19514 26464 31726
rect 26712 30190 26740 31726
rect 26700 30184 26752 30190
rect 26700 30126 26752 30132
rect 26514 29880 26570 29889
rect 26514 29815 26570 29824
rect 26528 29714 26556 29815
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 26516 29572 26568 29578
rect 26516 29514 26568 29520
rect 26528 28694 26556 29514
rect 26700 28960 26752 28966
rect 26700 28902 26752 28908
rect 26516 28688 26568 28694
rect 26516 28630 26568 28636
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26516 27668 26568 27674
rect 26516 27610 26568 27616
rect 26528 26518 26556 27610
rect 26516 26512 26568 26518
rect 26516 26454 26568 26460
rect 26528 25702 26556 26454
rect 26620 26042 26648 28494
rect 26712 28082 26740 28902
rect 26804 28082 26832 36094
rect 26976 36032 27028 36038
rect 26976 35974 27028 35980
rect 26988 35086 27016 35974
rect 27356 35698 27384 37810
rect 27540 37806 27568 38406
rect 27620 38354 27672 38360
rect 27620 38208 27672 38214
rect 27672 38168 27752 38196
rect 27620 38150 27672 38156
rect 27528 37800 27580 37806
rect 27528 37742 27580 37748
rect 27528 37664 27580 37670
rect 27528 37606 27580 37612
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27448 36310 27476 36518
rect 27436 36304 27488 36310
rect 27436 36246 27488 36252
rect 27436 36168 27488 36174
rect 27436 36110 27488 36116
rect 27448 35834 27476 36110
rect 27436 35828 27488 35834
rect 27436 35770 27488 35776
rect 27344 35692 27396 35698
rect 27344 35634 27396 35640
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 26976 35080 27028 35086
rect 26976 35022 27028 35028
rect 27264 34678 27292 35226
rect 27252 34672 27304 34678
rect 27252 34614 27304 34620
rect 27252 34400 27304 34406
rect 27252 34342 27304 34348
rect 27264 34066 27292 34342
rect 27252 34060 27304 34066
rect 27252 34002 27304 34008
rect 27068 32904 27120 32910
rect 27068 32846 27120 32852
rect 27080 31278 27108 32846
rect 27160 32768 27212 32774
rect 27160 32710 27212 32716
rect 27172 32570 27200 32710
rect 27160 32564 27212 32570
rect 27160 32506 27212 32512
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 27172 31929 27200 31962
rect 27158 31920 27214 31929
rect 27158 31855 27214 31864
rect 27356 31754 27384 35634
rect 27436 35624 27488 35630
rect 27436 35566 27488 35572
rect 27448 35086 27476 35566
rect 27436 35080 27488 35086
rect 27436 35022 27488 35028
rect 27436 34196 27488 34202
rect 27436 34138 27488 34144
rect 27448 33862 27476 34138
rect 27540 34066 27568 37606
rect 27724 35086 27752 38168
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27816 37330 27844 37742
rect 27804 37324 27856 37330
rect 27804 37266 27856 37272
rect 27804 36236 27856 36242
rect 27804 36178 27856 36184
rect 27816 35630 27844 36178
rect 27804 35624 27856 35630
rect 27804 35566 27856 35572
rect 27712 35080 27764 35086
rect 27712 35022 27764 35028
rect 27528 34060 27580 34066
rect 27528 34002 27580 34008
rect 27724 33930 27752 35022
rect 27908 34678 27936 38490
rect 30300 38282 30328 38490
rect 31208 38344 31260 38350
rect 31036 38304 31208 38332
rect 29828 38276 29880 38282
rect 29828 38218 29880 38224
rect 30288 38276 30340 38282
rect 30288 38218 30340 38224
rect 29276 38208 29328 38214
rect 29276 38150 29328 38156
rect 29288 38010 29316 38150
rect 29840 38010 29868 38218
rect 29276 38004 29328 38010
rect 29276 37946 29328 37952
rect 29828 38004 29880 38010
rect 29828 37946 29880 37952
rect 27988 37868 28040 37874
rect 27988 37810 28040 37816
rect 29184 37868 29236 37874
rect 29184 37810 29236 37816
rect 27896 34672 27948 34678
rect 27896 34614 27948 34620
rect 27908 34542 27936 34614
rect 27896 34536 27948 34542
rect 27896 34478 27948 34484
rect 27712 33924 27764 33930
rect 27712 33866 27764 33872
rect 27436 33856 27488 33862
rect 27436 33798 27488 33804
rect 27896 32836 27948 32842
rect 27896 32778 27948 32784
rect 27172 31726 27384 31754
rect 27908 31754 27936 32778
rect 28000 32026 28028 37810
rect 29196 37330 29224 37810
rect 29184 37324 29236 37330
rect 29184 37266 29236 37272
rect 28264 36916 28316 36922
rect 28264 36858 28316 36864
rect 28276 36106 28304 36858
rect 28724 36712 28776 36718
rect 28724 36654 28776 36660
rect 28264 36100 28316 36106
rect 28264 36042 28316 36048
rect 28276 35290 28304 36042
rect 28736 36038 28764 36654
rect 29288 36530 29316 37946
rect 30300 37942 30328 38218
rect 30288 37936 30340 37942
rect 30288 37878 30340 37884
rect 29736 36848 29788 36854
rect 29736 36790 29788 36796
rect 29012 36502 29316 36530
rect 28724 36032 28776 36038
rect 28724 35974 28776 35980
rect 28264 35284 28316 35290
rect 28264 35226 28316 35232
rect 28264 35148 28316 35154
rect 28264 35090 28316 35096
rect 27988 32020 28040 32026
rect 27988 31962 28040 31968
rect 27908 31726 28212 31754
rect 27068 31272 27120 31278
rect 27068 31214 27120 31220
rect 27080 30734 27108 31214
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 26976 30592 27028 30598
rect 26976 30534 27028 30540
rect 26988 30190 27016 30534
rect 27172 30326 27200 31726
rect 27896 31340 27948 31346
rect 27896 31282 27948 31288
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 27712 31136 27764 31142
rect 27712 31078 27764 31084
rect 27160 30320 27212 30326
rect 27160 30262 27212 30268
rect 26884 30184 26936 30190
rect 26884 30126 26936 30132
rect 26976 30184 27028 30190
rect 26976 30126 27028 30132
rect 26896 30036 26924 30126
rect 26896 30008 27016 30036
rect 26988 28994 27016 30008
rect 26896 28966 27016 28994
rect 26700 28076 26752 28082
rect 26700 28018 26752 28024
rect 26792 28076 26844 28082
rect 26792 28018 26844 28024
rect 26712 26518 26740 28018
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 26608 26036 26660 26042
rect 26608 25978 26660 25984
rect 26516 25696 26568 25702
rect 26516 25638 26568 25644
rect 26620 25294 26648 25978
rect 26712 25294 26740 26454
rect 26516 25288 26568 25294
rect 26516 25230 26568 25236
rect 26608 25288 26660 25294
rect 26608 25230 26660 25236
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26528 24750 26556 25230
rect 26712 24886 26740 25230
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 26516 24744 26568 24750
rect 26516 24686 26568 24692
rect 26700 24744 26752 24750
rect 26700 24686 26752 24692
rect 26608 24676 26660 24682
rect 26608 24618 26660 24624
rect 26620 24313 26648 24618
rect 26712 24410 26740 24686
rect 26700 24404 26752 24410
rect 26700 24346 26752 24352
rect 26606 24304 26662 24313
rect 26606 24239 26662 24248
rect 26620 24206 26648 24239
rect 26804 24206 26832 28018
rect 26896 25945 26924 28966
rect 27068 28960 27120 28966
rect 27068 28902 27120 28908
rect 27080 28626 27108 28902
rect 27068 28620 27120 28626
rect 27068 28562 27120 28568
rect 27068 28484 27120 28490
rect 27068 28426 27120 28432
rect 26974 28384 27030 28393
rect 26974 28319 27030 28328
rect 26988 28150 27016 28319
rect 27080 28218 27108 28426
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 26976 28144 27028 28150
rect 26976 28086 27028 28092
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 27080 26042 27108 26318
rect 27068 26036 27120 26042
rect 27068 25978 27120 25984
rect 26882 25936 26938 25945
rect 26882 25871 26938 25880
rect 26896 25498 26924 25871
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 26884 25356 26936 25362
rect 26884 25298 26936 25304
rect 26896 24274 26924 25298
rect 27066 24848 27122 24857
rect 27066 24783 27122 24792
rect 26884 24268 26936 24274
rect 26884 24210 26936 24216
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26516 24132 26568 24138
rect 26516 24074 26568 24080
rect 26976 24132 27028 24138
rect 26976 24074 27028 24080
rect 26528 23798 26556 24074
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 26528 23186 26556 23734
rect 26988 23497 27016 24074
rect 27080 23730 27108 24783
rect 27068 23724 27120 23730
rect 27068 23666 27120 23672
rect 26974 23488 27030 23497
rect 26974 23423 27030 23432
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26608 23112 26660 23118
rect 26608 23054 26660 23060
rect 26620 20058 26648 23054
rect 27068 23044 27120 23050
rect 27068 22986 27120 22992
rect 27080 22817 27108 22986
rect 27066 22808 27122 22817
rect 27066 22743 27122 22752
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 26988 22098 27016 22578
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 26884 21956 26936 21962
rect 26884 21898 26936 21904
rect 26792 21548 26844 21554
rect 26792 21490 26844 21496
rect 26804 20942 26832 21490
rect 26896 21146 26924 21898
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 26884 21140 26936 21146
rect 26884 21082 26936 21088
rect 26792 20936 26844 20942
rect 26844 20896 26924 20924
rect 26792 20878 26844 20884
rect 26608 20052 26660 20058
rect 26608 19994 26660 20000
rect 26896 19854 26924 20896
rect 26988 20874 27016 21422
rect 27172 21146 27200 30262
rect 27252 30184 27304 30190
rect 27252 30126 27304 30132
rect 27264 29850 27292 30126
rect 27252 29844 27304 29850
rect 27252 29786 27304 29792
rect 27252 28076 27304 28082
rect 27252 28018 27304 28024
rect 27264 27674 27292 28018
rect 27252 27668 27304 27674
rect 27252 27610 27304 27616
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 27448 26450 27476 26726
rect 27436 26444 27488 26450
rect 27436 26386 27488 26392
rect 27540 26330 27568 27406
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27448 26302 27568 26330
rect 27448 25906 27476 26302
rect 27632 26042 27660 26930
rect 27620 26036 27672 26042
rect 27620 25978 27672 25984
rect 27436 25900 27488 25906
rect 27436 25842 27488 25848
rect 27448 24886 27476 25842
rect 27436 24880 27488 24886
rect 27436 24822 27488 24828
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27356 23730 27384 24142
rect 27252 23724 27304 23730
rect 27252 23666 27304 23672
rect 27344 23724 27396 23730
rect 27344 23666 27396 23672
rect 27264 23361 27292 23666
rect 27250 23352 27306 23361
rect 27250 23287 27306 23296
rect 27252 23180 27304 23186
rect 27252 23122 27304 23128
rect 27264 22778 27292 23122
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27250 22672 27306 22681
rect 27356 22642 27384 23666
rect 27250 22607 27252 22616
rect 27304 22607 27306 22616
rect 27344 22636 27396 22642
rect 27252 22578 27304 22584
rect 27344 22578 27396 22584
rect 27448 22094 27476 24822
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27264 22066 27476 22094
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 27264 20942 27292 22066
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27356 21554 27384 21966
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27160 20936 27212 20942
rect 27160 20878 27212 20884
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 26976 20868 27028 20874
rect 26976 20810 27028 20816
rect 26884 19848 26936 19854
rect 26884 19790 26936 19796
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26608 19372 26660 19378
rect 26608 19314 26660 19320
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26620 18834 26648 19314
rect 26804 18970 26832 19314
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26424 18692 26476 18698
rect 26424 18634 26476 18640
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25688 17128 25740 17134
rect 25688 17070 25740 17076
rect 25240 16918 25452 16946
rect 25148 16782 25268 16810
rect 25134 16144 25190 16153
rect 25134 16079 25136 16088
rect 25188 16079 25190 16088
rect 25136 16050 25188 16056
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24780 12628 24808 14350
rect 24964 14074 24992 14418
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25056 14074 25084 14350
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 25148 13938 25176 15642
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 25136 13932 25188 13938
rect 25136 13874 25188 13880
rect 24872 13841 24900 13874
rect 24858 13832 24914 13841
rect 24914 13790 24992 13818
rect 24858 13767 24914 13776
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 24872 12782 24900 13398
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24780 12600 24900 12628
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 11898 24808 12174
rect 24872 12170 24900 12600
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24492 11824 24544 11830
rect 24490 11792 24492 11801
rect 24676 11824 24728 11830
rect 24544 11792 24546 11801
rect 24308 11756 24360 11762
rect 24676 11766 24728 11772
rect 24490 11727 24546 11736
rect 24308 11698 24360 11704
rect 24320 11014 24348 11698
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 24136 8634 24164 8910
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24228 8514 24256 10406
rect 24320 9110 24348 10950
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24398 10024 24454 10033
rect 24504 9994 24532 10202
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24398 9959 24454 9968
rect 24492 9988 24544 9994
rect 24308 9104 24360 9110
rect 24308 9046 24360 9052
rect 24412 8974 24440 9959
rect 24492 9930 24544 9936
rect 24492 9716 24544 9722
rect 24492 9658 24544 9664
rect 24504 9489 24532 9658
rect 24490 9480 24546 9489
rect 24490 9415 24546 9424
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24136 8486 24256 8514
rect 24306 8528 24362 8537
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23112 6860 23164 6866
rect 23112 6802 23164 6808
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 23124 6322 23152 6802
rect 23204 6724 23256 6730
rect 23204 6666 23256 6672
rect 23216 6458 23244 6666
rect 23204 6452 23256 6458
rect 23204 6394 23256 6400
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22848 5574 22876 6054
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22940 5234 22968 5714
rect 23400 5234 23428 5714
rect 23860 5710 23888 6190
rect 23952 5710 23980 6938
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23940 5704 23992 5710
rect 24044 5692 24072 7822
rect 24136 7410 24164 8486
rect 24306 8463 24362 8472
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24136 6458 24164 7346
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24124 5704 24176 5710
rect 24044 5664 24124 5692
rect 23940 5646 23992 5652
rect 24124 5646 24176 5652
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23492 5302 23520 5510
rect 23480 5296 23532 5302
rect 23480 5238 23532 5244
rect 23860 5234 23888 5646
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23216 4826 23244 5170
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23400 4690 23428 5170
rect 23952 5030 23980 5646
rect 24320 5302 24348 8463
rect 24412 6322 24440 8910
rect 24504 8838 24532 9415
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24596 7410 24624 9998
rect 24780 9926 24808 11834
rect 24872 11626 24900 12106
rect 24860 11620 24912 11626
rect 24860 11562 24912 11568
rect 24872 10538 24900 11562
rect 24964 11150 24992 13790
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25056 12889 25084 13262
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25042 12880 25098 12889
rect 25042 12815 25098 12824
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24860 10532 24912 10538
rect 24860 10474 24912 10480
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 25056 9586 25084 12718
rect 25148 12306 25176 12922
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25240 10606 25268 16782
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25332 12850 25360 14010
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 25332 11898 25360 12242
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25320 11620 25372 11626
rect 25320 11562 25372 11568
rect 25332 11354 25360 11562
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 25044 9580 25096 9586
rect 25044 9522 25096 9528
rect 24688 8906 24716 9522
rect 24964 9382 24992 9522
rect 25044 9444 25096 9450
rect 25044 9386 25096 9392
rect 24952 9376 25004 9382
rect 25056 9353 25084 9386
rect 24952 9318 25004 9324
rect 25042 9344 25098 9353
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24676 8900 24728 8906
rect 24676 8842 24728 8848
rect 24780 7410 24808 8978
rect 24964 8566 24992 9318
rect 25042 9279 25098 9288
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24964 7478 24992 8298
rect 24952 7472 25004 7478
rect 24952 7414 25004 7420
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 25148 7206 25176 8774
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 24964 6866 24992 7142
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25148 6458 25176 6734
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24952 6316 25004 6322
rect 24952 6258 25004 6264
rect 24596 5914 24624 6258
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24964 5710 24992 6258
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24676 5568 24728 5574
rect 24676 5510 24728 5516
rect 24308 5296 24360 5302
rect 24308 5238 24360 5244
rect 23940 5024 23992 5030
rect 23940 4966 23992 4972
rect 24688 4826 24716 5510
rect 24964 5098 24992 5646
rect 24952 5092 25004 5098
rect 24952 5034 25004 5040
rect 25136 5024 25188 5030
rect 25136 4966 25188 4972
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 22940 3942 22968 4558
rect 24032 4548 24084 4554
rect 24032 4490 24084 4496
rect 24044 4214 24072 4490
rect 25148 4282 25176 4966
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 25228 4752 25280 4758
rect 25228 4694 25280 4700
rect 25240 4622 25268 4694
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25332 4282 25360 4762
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 25320 4276 25372 4282
rect 25320 4218 25372 4224
rect 24032 4208 24084 4214
rect 25332 4185 25360 4218
rect 24032 4150 24084 4156
rect 25318 4176 25374 4185
rect 24044 4010 24072 4150
rect 25318 4111 25374 4120
rect 24032 4004 24084 4010
rect 24032 3946 24084 3952
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 25424 3058 25452 16918
rect 25884 16590 25912 18566
rect 26436 17241 26464 18634
rect 26620 18086 26648 18770
rect 27172 18290 27200 20878
rect 27540 20330 27568 24754
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27632 23730 27660 24006
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27724 22642 27752 31078
rect 27908 30190 27936 31282
rect 28000 30938 28028 31282
rect 28092 31249 28120 31282
rect 28078 31240 28134 31249
rect 28184 31226 28212 31726
rect 28276 31346 28304 35090
rect 28540 34536 28592 34542
rect 28540 34478 28592 34484
rect 28446 34232 28502 34241
rect 28446 34167 28502 34176
rect 28460 33862 28488 34167
rect 28356 33856 28408 33862
rect 28356 33798 28408 33804
rect 28448 33856 28500 33862
rect 28448 33798 28500 33804
rect 28368 33658 28396 33798
rect 28356 33652 28408 33658
rect 28356 33594 28408 33600
rect 28552 33590 28580 34478
rect 28632 34060 28684 34066
rect 28632 34002 28684 34008
rect 28540 33584 28592 33590
rect 28540 33526 28592 33532
rect 28448 33448 28500 33454
rect 28448 33390 28500 33396
rect 28460 33114 28488 33390
rect 28448 33108 28500 33114
rect 28448 33050 28500 33056
rect 28448 32836 28500 32842
rect 28448 32778 28500 32784
rect 28356 32020 28408 32026
rect 28356 31962 28408 31968
rect 28368 31657 28396 31962
rect 28354 31648 28410 31657
rect 28354 31583 28410 31592
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28184 31198 28304 31226
rect 28078 31175 28134 31184
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 27988 30932 28040 30938
rect 27988 30874 28040 30880
rect 27896 30184 27948 30190
rect 27896 30126 27948 30132
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 28000 29034 28028 29446
rect 27988 29028 28040 29034
rect 27988 28970 28040 28976
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 27804 27396 27856 27402
rect 27804 27338 27856 27344
rect 27816 27062 27844 27338
rect 27804 27056 27856 27062
rect 27804 26998 27856 27004
rect 27804 26308 27856 26314
rect 27908 26296 27936 28358
rect 27856 26268 27936 26296
rect 27804 26250 27856 26256
rect 27816 26081 27844 26250
rect 28000 26194 28028 28970
rect 27908 26166 28028 26194
rect 27802 26072 27858 26081
rect 27802 26007 27858 26016
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27632 22166 27660 22578
rect 27620 22160 27672 22166
rect 27620 22102 27672 22108
rect 27816 21962 27844 24142
rect 27804 21956 27856 21962
rect 27804 21898 27856 21904
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27632 21146 27660 21830
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26608 18080 26660 18086
rect 26608 18022 26660 18028
rect 26608 17604 26660 17610
rect 26712 17592 26740 18158
rect 27172 17882 27200 18226
rect 27160 17876 27212 17882
rect 27160 17818 27212 17824
rect 26660 17564 26740 17592
rect 26608 17546 26660 17552
rect 26422 17232 26478 17241
rect 26422 17167 26478 17176
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 26240 16040 26292 16046
rect 26424 16040 26476 16046
rect 26240 15982 26292 15988
rect 26344 16000 26424 16028
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25516 15162 25544 15438
rect 26252 15434 26280 15982
rect 26344 15502 26372 16000
rect 26424 15982 26476 15988
rect 26516 15972 26568 15978
rect 26516 15914 26568 15920
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26240 15428 26292 15434
rect 26240 15370 26292 15376
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 26252 15094 26280 15370
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25780 14816 25832 14822
rect 25780 14758 25832 14764
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25516 13530 25544 13874
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25608 12986 25636 14758
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25700 12918 25728 13874
rect 25792 13326 25820 14758
rect 25884 14074 25912 14894
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 25872 13796 25924 13802
rect 25872 13738 25924 13744
rect 25884 13433 25912 13738
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 25870 13424 25926 13433
rect 25870 13359 25926 13368
rect 25976 13326 26004 13670
rect 26252 13326 26280 13670
rect 26436 13410 26464 15574
rect 26528 15094 26556 15914
rect 26620 15586 26648 17546
rect 27068 17128 27120 17134
rect 27068 17070 27120 17076
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 26896 15978 26924 16730
rect 26884 15972 26936 15978
rect 26884 15914 26936 15920
rect 26896 15638 26924 15914
rect 26884 15632 26936 15638
rect 26620 15558 26832 15586
rect 26884 15574 26936 15580
rect 26516 15088 26568 15094
rect 26516 15030 26568 15036
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26712 13938 26740 14758
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26436 13382 26556 13410
rect 26528 13326 26556 13382
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26516 13320 26568 13326
rect 26568 13280 26648 13308
rect 26516 13262 26568 13268
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 25688 12912 25740 12918
rect 25688 12854 25740 12860
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25700 12238 25728 12582
rect 25884 12306 25912 13126
rect 26344 12850 26372 13126
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25792 11898 25820 12038
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25596 11144 25648 11150
rect 25594 11112 25596 11121
rect 25648 11112 25650 11121
rect 25792 11082 25820 11834
rect 25884 11150 25912 12242
rect 26344 12238 26372 12650
rect 26436 12594 26464 13262
rect 26620 12850 26648 13280
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26608 12640 26660 12646
rect 26436 12566 26556 12594
rect 26608 12582 26660 12588
rect 26422 12472 26478 12481
rect 26422 12407 26478 12416
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 25976 12073 26004 12106
rect 25962 12064 26018 12073
rect 25962 11999 26018 12008
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25594 11047 25650 11056
rect 25780 11076 25832 11082
rect 26436 11064 26464 12407
rect 26528 11801 26556 12566
rect 26514 11792 26570 11801
rect 26514 11727 26570 11736
rect 25780 11018 25832 11024
rect 26344 11036 26464 11064
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25608 9489 25636 9522
rect 25594 9480 25650 9489
rect 25594 9415 25650 9424
rect 25792 9042 25820 11018
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 26240 11008 26292 11014
rect 26240 10950 26292 10956
rect 25884 10810 25912 10950
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 26252 10062 26280 10950
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 25870 9616 25926 9625
rect 25870 9551 25872 9560
rect 25924 9551 25926 9560
rect 25964 9580 26016 9586
rect 25872 9522 25924 9528
rect 25964 9522 26016 9528
rect 25976 9489 26004 9522
rect 25962 9480 26018 9489
rect 25962 9415 26018 9424
rect 26344 9382 26372 11036
rect 26424 10600 26476 10606
rect 26528 10588 26556 11727
rect 26620 10810 26648 12582
rect 26712 12306 26740 13874
rect 26804 13818 26832 15558
rect 26896 13938 26924 15574
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26988 15162 27016 15438
rect 27080 15162 27108 17070
rect 27264 16658 27292 19314
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27160 16176 27212 16182
rect 27160 16118 27212 16124
rect 27172 15910 27200 16118
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27172 15638 27200 15846
rect 27160 15632 27212 15638
rect 27160 15574 27212 15580
rect 26976 15156 27028 15162
rect 26976 15098 27028 15104
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27264 14618 27292 16594
rect 27252 14612 27304 14618
rect 27252 14554 27304 14560
rect 27356 14521 27384 19450
rect 27724 18222 27752 21490
rect 27816 21486 27844 21898
rect 27908 21690 27936 26166
rect 27988 24948 28040 24954
rect 27988 24890 28040 24896
rect 28000 23798 28028 24890
rect 27988 23792 28040 23798
rect 27988 23734 28040 23740
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 27908 19378 27936 19858
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 28000 19334 28028 21966
rect 28092 19854 28120 31078
rect 28276 28994 28304 31198
rect 28184 28966 28304 28994
rect 28184 22166 28212 28966
rect 28356 26240 28408 26246
rect 28356 26182 28408 26188
rect 28264 25968 28316 25974
rect 28264 25910 28316 25916
rect 28276 24818 28304 25910
rect 28368 25906 28396 26182
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 28356 24948 28408 24954
rect 28356 24890 28408 24896
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28368 24664 28396 24890
rect 28276 24636 28396 24664
rect 28276 23798 28304 24636
rect 28460 24562 28488 32778
rect 28552 32502 28580 33526
rect 28644 32978 28672 34002
rect 28632 32972 28684 32978
rect 28632 32914 28684 32920
rect 28540 32496 28592 32502
rect 28540 32438 28592 32444
rect 28632 32496 28684 32502
rect 28632 32438 28684 32444
rect 28552 30326 28580 32438
rect 28644 31754 28672 32438
rect 28632 31748 28684 31754
rect 28632 31690 28684 31696
rect 28632 31408 28684 31414
rect 28632 31350 28684 31356
rect 28644 31113 28672 31350
rect 28630 31104 28686 31113
rect 28630 31039 28686 31048
rect 28540 30320 28592 30326
rect 28540 30262 28592 30268
rect 28736 29306 28764 35974
rect 29012 35562 29040 36502
rect 29092 36372 29144 36378
rect 29092 36314 29144 36320
rect 29000 35556 29052 35562
rect 29000 35498 29052 35504
rect 29104 34610 29132 36314
rect 29288 36174 29316 36502
rect 29368 36372 29420 36378
rect 29368 36314 29420 36320
rect 29380 36174 29408 36314
rect 29460 36304 29512 36310
rect 29460 36246 29512 36252
rect 29276 36168 29328 36174
rect 29276 36110 29328 36116
rect 29368 36168 29420 36174
rect 29368 36110 29420 36116
rect 29368 36032 29420 36038
rect 29368 35974 29420 35980
rect 29184 35692 29236 35698
rect 29184 35634 29236 35640
rect 29092 34604 29144 34610
rect 29092 34546 29144 34552
rect 28908 32972 28960 32978
rect 28908 32914 28960 32920
rect 28816 31476 28868 31482
rect 28816 31418 28868 31424
rect 28828 31346 28856 31418
rect 28816 31340 28868 31346
rect 28816 31282 28868 31288
rect 28814 31240 28870 31249
rect 28814 31175 28870 31184
rect 28828 31142 28856 31175
rect 28816 31136 28868 31142
rect 28816 31078 28868 31084
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 28828 29850 28856 30670
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28920 29714 28948 32914
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 29012 32366 29040 32846
rect 29104 32570 29132 34546
rect 29196 34474 29224 35634
rect 29380 35494 29408 35974
rect 29472 35698 29500 36246
rect 29748 36174 29776 36790
rect 30012 36644 30064 36650
rect 30012 36586 30064 36592
rect 30024 36174 30052 36586
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 30012 36168 30064 36174
rect 30012 36110 30064 36116
rect 30932 36168 30984 36174
rect 30932 36110 30984 36116
rect 29460 35692 29512 35698
rect 29460 35634 29512 35640
rect 29552 35692 29604 35698
rect 29552 35634 29604 35640
rect 29276 35488 29328 35494
rect 29276 35430 29328 35436
rect 29368 35488 29420 35494
rect 29368 35430 29420 35436
rect 29184 34468 29236 34474
rect 29184 34410 29236 34416
rect 29092 32564 29144 32570
rect 29092 32506 29144 32512
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 29012 31890 29040 32302
rect 29000 31884 29052 31890
rect 29000 31826 29052 31832
rect 29288 31754 29316 35430
rect 29380 34678 29408 35430
rect 29460 35080 29512 35086
rect 29460 35022 29512 35028
rect 29368 34672 29420 34678
rect 29368 34614 29420 34620
rect 29472 34610 29500 35022
rect 29564 35018 29592 35634
rect 29552 35012 29604 35018
rect 29552 34954 29604 34960
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 29564 34066 29592 34954
rect 29920 34672 29972 34678
rect 29920 34614 29972 34620
rect 29736 34400 29788 34406
rect 29736 34342 29788 34348
rect 29552 34060 29604 34066
rect 29552 34002 29604 34008
rect 29748 33998 29776 34342
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29736 33312 29788 33318
rect 29736 33254 29788 33260
rect 29748 32774 29776 33254
rect 29736 32768 29788 32774
rect 29736 32710 29788 32716
rect 29644 32564 29696 32570
rect 29644 32506 29696 32512
rect 29656 32434 29684 32506
rect 29748 32434 29776 32710
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29656 31754 29684 32370
rect 29932 32348 29960 34614
rect 30024 34610 30052 36110
rect 30380 36032 30432 36038
rect 30380 35974 30432 35980
rect 30748 36032 30800 36038
rect 30748 35974 30800 35980
rect 30392 35766 30420 35974
rect 30380 35760 30432 35766
rect 30380 35702 30432 35708
rect 30472 35760 30524 35766
rect 30472 35702 30524 35708
rect 30484 35290 30512 35702
rect 30760 35630 30788 35974
rect 30840 35760 30892 35766
rect 30840 35702 30892 35708
rect 30852 35630 30880 35702
rect 30748 35624 30800 35630
rect 30748 35566 30800 35572
rect 30840 35624 30892 35630
rect 30840 35566 30892 35572
rect 30944 35290 30972 36110
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 30932 35284 30984 35290
rect 30932 35226 30984 35232
rect 30012 34604 30064 34610
rect 30012 34546 30064 34552
rect 30380 34604 30432 34610
rect 30380 34546 30432 34552
rect 30024 32858 30052 34546
rect 30392 34202 30420 34546
rect 30656 34400 30708 34406
rect 30656 34342 30708 34348
rect 30668 34202 30696 34342
rect 30380 34196 30432 34202
rect 30380 34138 30432 34144
rect 30656 34196 30708 34202
rect 30656 34138 30708 34144
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30196 33312 30248 33318
rect 30196 33254 30248 33260
rect 30024 32830 30144 32858
rect 30116 32434 30144 32830
rect 30208 32502 30236 33254
rect 30392 32570 30420 33934
rect 30472 33924 30524 33930
rect 30472 33866 30524 33872
rect 30380 32564 30432 32570
rect 30380 32506 30432 32512
rect 30196 32496 30248 32502
rect 30196 32438 30248 32444
rect 30104 32428 30156 32434
rect 30104 32370 30156 32376
rect 30012 32360 30064 32366
rect 29932 32320 30012 32348
rect 30012 32302 30064 32308
rect 29104 31726 29316 31754
rect 29472 31726 29684 31754
rect 29000 31680 29052 31686
rect 29000 31622 29052 31628
rect 29012 31482 29040 31622
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 29104 31346 29132 31726
rect 29000 31340 29052 31346
rect 29000 31282 29052 31288
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 29012 30938 29040 31282
rect 29288 31142 29316 31282
rect 29276 31136 29328 31142
rect 29276 31078 29328 31084
rect 29000 30932 29052 30938
rect 29000 30874 29052 30880
rect 29276 30864 29328 30870
rect 29276 30806 29328 30812
rect 29184 30728 29236 30734
rect 29184 30670 29236 30676
rect 29000 30660 29052 30666
rect 29000 30602 29052 30608
rect 28908 29708 28960 29714
rect 28828 29668 28908 29696
rect 28724 29300 28776 29306
rect 28724 29242 28776 29248
rect 28540 28416 28592 28422
rect 28540 28358 28592 28364
rect 28552 27062 28580 28358
rect 28828 28014 28856 29668
rect 28908 29650 28960 29656
rect 28908 29504 28960 29510
rect 28908 29446 28960 29452
rect 28920 29102 28948 29446
rect 28908 29096 28960 29102
rect 28908 29038 28960 29044
rect 29012 28966 29040 30602
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 29104 30190 29132 30534
rect 29092 30184 29144 30190
rect 29092 30126 29144 30132
rect 29000 28960 29052 28966
rect 29000 28902 29052 28908
rect 28954 28688 29006 28694
rect 28954 28630 29006 28636
rect 29090 28656 29146 28665
rect 28966 28540 28994 28630
rect 29196 28642 29224 30670
rect 29288 30326 29316 30806
rect 29276 30320 29328 30326
rect 29276 30262 29328 30268
rect 29472 29646 29500 31726
rect 29920 31340 29972 31346
rect 29920 31282 29972 31288
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 29840 29646 29868 29990
rect 29460 29640 29512 29646
rect 29460 29582 29512 29588
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29146 28614 29408 28642
rect 29090 28591 29146 28600
rect 29104 28558 29132 28591
rect 29092 28552 29144 28558
rect 28966 28529 29040 28540
rect 28966 28520 29054 28529
rect 28966 28512 28998 28520
rect 29092 28494 29144 28500
rect 29184 28552 29236 28558
rect 29184 28494 29236 28500
rect 28998 28455 29054 28464
rect 29196 28218 29224 28494
rect 29184 28212 29236 28218
rect 29184 28154 29236 28160
rect 28998 28112 29054 28121
rect 28998 28048 29000 28056
rect 29052 28048 29054 28056
rect 28998 28047 29054 28048
rect 29092 28076 29144 28082
rect 29000 28042 29052 28047
rect 29144 28036 29200 28064
rect 29092 28018 29144 28024
rect 28816 28008 28868 28014
rect 28816 27950 28868 27956
rect 29172 27962 29200 28036
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28540 27056 28592 27062
rect 28540 26998 28592 27004
rect 28644 26994 28672 27270
rect 28632 26988 28684 26994
rect 28632 26930 28684 26936
rect 28724 26988 28776 26994
rect 28724 26930 28776 26936
rect 28540 25152 28592 25158
rect 28644 25129 28672 26930
rect 28736 26246 28764 26930
rect 28724 26240 28776 26246
rect 28724 26182 28776 26188
rect 28828 25838 28856 27950
rect 29172 27934 29224 27962
rect 29196 27674 29224 27934
rect 29184 27668 29236 27674
rect 29184 27610 29236 27616
rect 28908 27600 28960 27606
rect 28908 27542 28960 27548
rect 28920 26994 28948 27542
rect 29092 27464 29144 27470
rect 29092 27406 29144 27412
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 29104 26382 29132 27406
rect 29092 26376 29144 26382
rect 28920 26324 29092 26330
rect 28920 26318 29144 26324
rect 28920 26302 29132 26318
rect 28920 25974 28948 26302
rect 29092 26240 29144 26246
rect 29092 26182 29144 26188
rect 28908 25968 28960 25974
rect 28908 25910 28960 25916
rect 29000 25900 29052 25906
rect 29000 25842 29052 25848
rect 28816 25832 28868 25838
rect 28816 25774 28868 25780
rect 28540 25094 28592 25100
rect 28630 25120 28686 25129
rect 28368 24534 28488 24562
rect 28264 23792 28316 23798
rect 28264 23734 28316 23740
rect 28368 22234 28396 24534
rect 28552 24070 28580 25094
rect 28630 25055 28686 25064
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28644 24410 28672 24754
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28736 23866 28764 24346
rect 28828 24274 28856 25774
rect 29012 25498 29040 25842
rect 29104 25838 29132 26182
rect 29092 25832 29144 25838
rect 29092 25774 29144 25780
rect 29000 25492 29052 25498
rect 29000 25434 29052 25440
rect 29196 25378 29224 27610
rect 29380 27470 29408 28614
rect 29472 28082 29500 29582
rect 29932 29306 29960 31282
rect 30024 29578 30052 32302
rect 30116 29714 30144 32370
rect 30484 31822 30512 33866
rect 30748 32836 30800 32842
rect 30748 32778 30800 32784
rect 30760 32570 30788 32778
rect 30748 32564 30800 32570
rect 30748 32506 30800 32512
rect 30564 32292 30616 32298
rect 30564 32234 30616 32240
rect 30576 31958 30604 32234
rect 30760 32026 30788 32506
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 30564 31952 30616 31958
rect 30564 31894 30616 31900
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30472 31816 30524 31822
rect 30472 31758 30524 31764
rect 30208 31482 30236 31758
rect 30392 31668 30420 31758
rect 30392 31640 30512 31668
rect 30196 31476 30248 31482
rect 30196 31418 30248 31424
rect 30208 30938 30236 31418
rect 30484 31142 30512 31640
rect 30576 31346 30604 31894
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 30472 31136 30524 31142
rect 30472 31078 30524 31084
rect 30196 30932 30248 30938
rect 30196 30874 30248 30880
rect 30104 29708 30156 29714
rect 30104 29650 30156 29656
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 29920 29300 29972 29306
rect 29920 29242 29972 29248
rect 30024 28994 30052 29514
rect 29932 28966 30052 28994
rect 29552 28960 29604 28966
rect 29552 28902 29604 28908
rect 29460 28076 29512 28082
rect 29460 28018 29512 28024
rect 29368 27464 29420 27470
rect 29368 27406 29420 27412
rect 29472 27334 29500 28018
rect 29460 27328 29512 27334
rect 29460 27270 29512 27276
rect 29564 27130 29592 28902
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 29748 28082 29776 28358
rect 29932 28150 29960 28966
rect 29920 28144 29972 28150
rect 30012 28144 30064 28150
rect 29920 28086 29972 28092
rect 30010 28112 30012 28121
rect 30064 28112 30066 28121
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29932 27606 29960 28086
rect 30116 28082 30144 29650
rect 30484 29628 30512 31078
rect 30852 30326 30880 32370
rect 31036 31754 31064 38304
rect 31208 38286 31260 38292
rect 32036 38344 32088 38350
rect 32036 38286 32088 38292
rect 34520 38344 34572 38350
rect 34520 38286 34572 38292
rect 31944 38208 31996 38214
rect 31944 38150 31996 38156
rect 31956 38010 31984 38150
rect 31944 38004 31996 38010
rect 31944 37946 31996 37952
rect 32048 37738 32076 38286
rect 32312 37868 32364 37874
rect 32312 37810 32364 37816
rect 32036 37732 32088 37738
rect 32036 37674 32088 37680
rect 31760 37664 31812 37670
rect 31760 37606 31812 37612
rect 31208 37324 31260 37330
rect 31208 37266 31260 37272
rect 31300 37324 31352 37330
rect 31300 37266 31352 37272
rect 31220 37126 31248 37266
rect 31116 37120 31168 37126
rect 31116 37062 31168 37068
rect 31208 37120 31260 37126
rect 31208 37062 31260 37068
rect 31128 36854 31156 37062
rect 31116 36848 31168 36854
rect 31116 36790 31168 36796
rect 31312 35154 31340 37266
rect 31772 36922 31800 37606
rect 32324 37194 32352 37810
rect 34532 37262 34560 38286
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34520 37256 34572 37262
rect 34520 37198 34572 37204
rect 37278 37224 37334 37233
rect 32312 37188 32364 37194
rect 37278 37159 37280 37168
rect 32312 37130 32364 37136
rect 37332 37159 37334 37168
rect 37280 37130 37332 37136
rect 33140 37120 33192 37126
rect 33140 37062 33192 37068
rect 37832 37120 37884 37126
rect 37832 37062 37884 37068
rect 31760 36916 31812 36922
rect 31760 36858 31812 36864
rect 32956 36780 33008 36786
rect 32956 36722 33008 36728
rect 32772 36576 32824 36582
rect 32772 36518 32824 36524
rect 32784 36242 32812 36518
rect 32772 36236 32824 36242
rect 32772 36178 32824 36184
rect 32680 36100 32732 36106
rect 32680 36042 32732 36048
rect 32692 35834 32720 36042
rect 32772 36032 32824 36038
rect 32772 35974 32824 35980
rect 32680 35828 32732 35834
rect 32680 35770 32732 35776
rect 31852 35488 31904 35494
rect 31852 35430 31904 35436
rect 31300 35148 31352 35154
rect 31300 35090 31352 35096
rect 31864 35086 31892 35430
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 31116 34944 31168 34950
rect 31116 34886 31168 34892
rect 31128 34542 31156 34886
rect 31116 34536 31168 34542
rect 31116 34478 31168 34484
rect 31392 34536 31444 34542
rect 31392 34478 31444 34484
rect 31404 34202 31432 34478
rect 31392 34196 31444 34202
rect 31392 34138 31444 34144
rect 31404 33862 31432 34138
rect 32692 33998 32720 35770
rect 32784 33998 32812 35974
rect 32968 35834 32996 36722
rect 33152 35834 33180 37062
rect 37844 36825 37872 37062
rect 37830 36816 37886 36825
rect 37830 36751 37886 36760
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34244 36032 34296 36038
rect 34244 35974 34296 35980
rect 34256 35834 34284 35974
rect 32956 35828 33008 35834
rect 32956 35770 33008 35776
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 34244 35828 34296 35834
rect 34244 35770 34296 35776
rect 33152 35714 33180 35770
rect 33152 35686 33548 35714
rect 33324 35624 33376 35630
rect 33324 35566 33376 35572
rect 33336 34542 33364 35566
rect 33324 34536 33376 34542
rect 33376 34496 33456 34524
rect 33324 34478 33376 34484
rect 32864 34196 32916 34202
rect 32864 34138 32916 34144
rect 32680 33992 32732 33998
rect 32680 33934 32732 33940
rect 32772 33992 32824 33998
rect 32772 33934 32824 33940
rect 31392 33856 31444 33862
rect 31392 33798 31444 33804
rect 31668 33584 31720 33590
rect 31668 33526 31720 33532
rect 31484 33040 31536 33046
rect 31484 32982 31536 32988
rect 31496 32502 31524 32982
rect 31484 32496 31536 32502
rect 31484 32438 31536 32444
rect 31484 32224 31536 32230
rect 31484 32166 31536 32172
rect 31116 31884 31168 31890
rect 31116 31826 31168 31832
rect 30944 31726 31064 31754
rect 30840 30320 30892 30326
rect 30840 30262 30892 30268
rect 30748 30252 30800 30258
rect 30748 30194 30800 30200
rect 30760 29850 30788 30194
rect 30748 29844 30800 29850
rect 30748 29786 30800 29792
rect 30656 29640 30708 29646
rect 30484 29600 30656 29628
rect 30708 29600 30788 29628
rect 30656 29582 30708 29588
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 30392 29306 30420 29514
rect 30380 29300 30432 29306
rect 30380 29242 30432 29248
rect 30380 28144 30432 28150
rect 30300 28104 30380 28132
rect 30010 28047 30066 28056
rect 30104 28076 30156 28082
rect 30104 28018 30156 28024
rect 29920 27600 29972 27606
rect 29920 27542 29972 27548
rect 29552 27124 29604 27130
rect 29552 27066 29604 27072
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 29288 26382 29316 26726
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29012 25350 29224 25378
rect 28908 24744 28960 24750
rect 28908 24686 28960 24692
rect 28920 24342 28948 24686
rect 28908 24336 28960 24342
rect 28908 24278 28960 24284
rect 28816 24268 28868 24274
rect 28816 24210 28868 24216
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28828 23322 28856 24210
rect 28816 23316 28868 23322
rect 28816 23258 28868 23264
rect 28724 22636 28776 22642
rect 28724 22578 28776 22584
rect 28356 22228 28408 22234
rect 28356 22170 28408 22176
rect 28172 22160 28224 22166
rect 28172 22102 28224 22108
rect 28736 22030 28764 22578
rect 28816 22568 28868 22574
rect 28816 22510 28868 22516
rect 28828 22098 28856 22510
rect 28816 22092 28868 22098
rect 28816 22034 28868 22040
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28724 22024 28776 22030
rect 28724 21966 28776 21972
rect 28356 21956 28408 21962
rect 28356 21898 28408 21904
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28368 21078 28396 21898
rect 28460 21486 28488 21898
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28356 21072 28408 21078
rect 28356 21014 28408 21020
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 28276 19718 28304 19994
rect 28460 19922 28488 20198
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28172 19712 28224 19718
rect 28172 19654 28224 19660
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 28184 19514 28212 19654
rect 28172 19508 28224 19514
rect 28172 19450 28224 19456
rect 28000 19306 28120 19334
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27632 17649 27660 17682
rect 27988 17672 28040 17678
rect 27618 17640 27674 17649
rect 27988 17614 28040 17620
rect 27618 17575 27674 17584
rect 28000 17066 28028 17614
rect 28092 17338 28120 19306
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28368 18358 28396 19110
rect 28552 19009 28580 21966
rect 28736 21554 28764 21966
rect 29012 21894 29040 25350
rect 29184 24336 29236 24342
rect 29184 24278 29236 24284
rect 29196 23866 29224 24278
rect 29184 23860 29236 23866
rect 29184 23802 29236 23808
rect 29656 23798 29684 25910
rect 29932 24818 29960 27542
rect 30116 26994 30144 28018
rect 30300 27878 30328 28104
rect 30380 28086 30432 28092
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 30392 27606 30420 27814
rect 30380 27600 30432 27606
rect 30656 27600 30708 27606
rect 30380 27542 30432 27548
rect 30484 27548 30656 27554
rect 30484 27542 30708 27548
rect 30484 27526 30696 27542
rect 30104 26988 30156 26994
rect 30104 26930 30156 26936
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 30300 26382 30328 26862
rect 30484 26382 30512 27526
rect 30760 27470 30788 29600
rect 30852 28082 30880 30262
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 30852 27606 30880 28018
rect 30840 27600 30892 27606
rect 30840 27542 30892 27548
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30760 26994 30788 27406
rect 30840 27396 30892 27402
rect 30840 27338 30892 27344
rect 30748 26988 30800 26994
rect 30748 26930 30800 26936
rect 30656 26512 30708 26518
rect 30656 26454 30708 26460
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 30472 26376 30524 26382
rect 30472 26318 30524 26324
rect 30380 25832 30432 25838
rect 30380 25774 30432 25780
rect 30392 25294 30420 25774
rect 30196 25288 30248 25294
rect 30196 25230 30248 25236
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 29920 24812 29972 24818
rect 29920 24754 29972 24760
rect 30208 24206 30236 25230
rect 30484 24682 30512 26318
rect 30564 26240 30616 26246
rect 30564 26182 30616 26188
rect 30472 24676 30524 24682
rect 30472 24618 30524 24624
rect 30576 24410 30604 26182
rect 30668 24954 30696 26454
rect 30748 26376 30800 26382
rect 30746 26344 30748 26353
rect 30800 26344 30802 26353
rect 30746 26279 30802 26288
rect 30656 24948 30708 24954
rect 30656 24890 30708 24896
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30380 24200 30432 24206
rect 30576 24188 30604 24346
rect 30668 24206 30696 24550
rect 30852 24206 30880 27338
rect 30432 24160 30604 24188
rect 30656 24200 30708 24206
rect 30380 24142 30432 24148
rect 30656 24142 30708 24148
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30748 24064 30800 24070
rect 30748 24006 30800 24012
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 29644 23792 29696 23798
rect 29644 23734 29696 23740
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29092 22432 29144 22438
rect 29092 22374 29144 22380
rect 29104 22094 29132 22374
rect 29472 22234 29500 22578
rect 30012 22568 30064 22574
rect 30012 22510 30064 22516
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 29104 22066 29224 22094
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 29104 20618 29132 21830
rect 29196 21554 29224 22066
rect 29748 22030 29776 22374
rect 29736 22024 29788 22030
rect 29736 21966 29788 21972
rect 29748 21690 29776 21966
rect 29920 21888 29972 21894
rect 29920 21830 29972 21836
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 29932 21486 29960 21830
rect 29920 21480 29972 21486
rect 29920 21422 29972 21428
rect 29460 21344 29512 21350
rect 29460 21286 29512 21292
rect 29920 21344 29972 21350
rect 29920 21286 29972 21292
rect 29012 20590 29132 20618
rect 29012 20534 29040 20590
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28632 20256 28684 20262
rect 28632 20198 28684 20204
rect 28644 19378 28672 20198
rect 28920 20058 28948 20402
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28538 19000 28594 19009
rect 28736 18970 28764 19790
rect 28920 19357 28948 19994
rect 29012 19922 29040 20470
rect 29472 20466 29500 21286
rect 29932 20942 29960 21286
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29092 20256 29144 20262
rect 29092 20198 29144 20204
rect 29276 20256 29328 20262
rect 29276 20198 29328 20204
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 29104 19802 29132 20198
rect 29288 19990 29316 20198
rect 29276 19984 29328 19990
rect 29276 19926 29328 19932
rect 29012 19774 29132 19802
rect 29012 19378 29040 19774
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 29196 19446 29224 19654
rect 29184 19440 29236 19446
rect 29184 19382 29236 19388
rect 29288 19378 29316 19926
rect 29000 19372 29052 19378
rect 28906 19348 28962 19357
rect 29000 19314 29052 19320
rect 29276 19372 29328 19378
rect 29276 19314 29328 19320
rect 28906 19283 28962 19292
rect 29380 19174 29408 20402
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29472 19378 29500 20198
rect 29564 19854 29592 20402
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29184 19168 29236 19174
rect 28906 19136 28962 19145
rect 29184 19110 29236 19116
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 28906 19071 28962 19080
rect 28538 18935 28594 18944
rect 28724 18964 28776 18970
rect 28356 18352 28408 18358
rect 28356 18294 28408 18300
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 28368 17338 28396 18158
rect 28552 18034 28580 18935
rect 28724 18906 28776 18912
rect 28816 18760 28868 18766
rect 28920 18748 28948 19071
rect 29196 18766 29224 19110
rect 29274 18864 29330 18873
rect 29380 18850 29408 19110
rect 29330 18822 29408 18850
rect 29274 18799 29330 18808
rect 28868 18720 28948 18748
rect 29184 18760 29236 18766
rect 28816 18702 28868 18708
rect 29184 18702 29236 18708
rect 28630 18048 28686 18057
rect 28552 18006 28630 18034
rect 28630 17983 28686 17992
rect 28908 17808 28960 17814
rect 28908 17750 28960 17756
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 28080 17332 28132 17338
rect 28080 17274 28132 17280
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 27988 17060 28040 17066
rect 27988 17002 28040 17008
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 27908 15502 27936 15914
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 27712 15428 27764 15434
rect 27712 15370 27764 15376
rect 27342 14512 27398 14521
rect 27342 14447 27398 14456
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26804 13790 26924 13818
rect 26792 13252 26844 13258
rect 26792 13194 26844 13200
rect 26804 12986 26832 13194
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 26896 12306 26924 13790
rect 27252 13728 27304 13734
rect 27252 13670 27304 13676
rect 27264 13530 27292 13670
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 26988 13382 27108 13410
rect 26988 13326 27016 13382
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26896 12209 26924 12242
rect 26882 12200 26938 12209
rect 26882 12135 26938 12144
rect 26700 12096 26752 12102
rect 26700 12038 26752 12044
rect 26712 11286 26740 12038
rect 26988 11830 27016 12786
rect 26792 11824 26844 11830
rect 26792 11766 26844 11772
rect 26976 11824 27028 11830
rect 26976 11766 27028 11772
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26804 11218 26832 11766
rect 26884 11756 26936 11762
rect 26884 11698 26936 11704
rect 26792 11212 26844 11218
rect 26792 11154 26844 11160
rect 26608 10804 26660 10810
rect 26608 10746 26660 10752
rect 26476 10560 26556 10588
rect 26424 10542 26476 10548
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25608 8430 25636 8910
rect 25700 8838 25728 8910
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25700 8090 25728 8774
rect 25792 8498 25820 8978
rect 26252 8974 26280 9318
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26344 8974 26372 9114
rect 26436 9110 26464 10542
rect 26896 10470 26924 11698
rect 26976 11552 27028 11558
rect 26976 11494 27028 11500
rect 26884 10464 26936 10470
rect 26884 10406 26936 10412
rect 26988 10062 27016 11494
rect 27080 10062 27108 13382
rect 27264 13326 27292 13466
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27264 12850 27292 13262
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27250 11928 27306 11937
rect 27250 11863 27306 11872
rect 27264 11830 27292 11863
rect 27252 11824 27304 11830
rect 27252 11766 27304 11772
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 27172 11354 27200 11494
rect 27264 11354 27292 11766
rect 27356 11762 27384 14447
rect 27528 13184 27580 13190
rect 27528 13126 27580 13132
rect 27540 11778 27568 13126
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27632 12442 27660 12786
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27448 11750 27568 11778
rect 27448 11354 27476 11750
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27172 11234 27200 11290
rect 27344 11280 27396 11286
rect 27172 11228 27344 11234
rect 27172 11222 27396 11228
rect 27172 11206 27384 11222
rect 27356 11150 27384 11206
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 27344 11144 27396 11150
rect 27540 11132 27568 11562
rect 27620 11144 27672 11150
rect 27540 11104 27620 11132
rect 27344 11086 27396 11092
rect 27620 11086 27672 11092
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 27068 10056 27120 10062
rect 27068 9998 27120 10004
rect 26516 9920 26568 9926
rect 26516 9862 26568 9868
rect 26424 9104 26476 9110
rect 26424 9046 26476 9052
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25976 7886 26004 8774
rect 26252 8634 26280 8774
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26528 8294 26556 9862
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26804 8974 26832 9318
rect 27172 9178 27200 11086
rect 27724 11014 27752 15370
rect 27804 15360 27856 15366
rect 27804 15302 27856 15308
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 27816 11626 27844 15302
rect 28000 15094 28028 15302
rect 27988 15088 28040 15094
rect 27988 15030 28040 15036
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27908 13530 27936 14962
rect 27988 14884 28040 14890
rect 27988 14826 28040 14832
rect 28000 14618 28028 14826
rect 27988 14612 28040 14618
rect 27988 14554 28040 14560
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 27896 13524 27948 13530
rect 27896 13466 27948 13472
rect 28000 13410 28028 14282
rect 28092 13818 28120 17274
rect 28736 17202 28764 17478
rect 28632 17196 28684 17202
rect 28632 17138 28684 17144
rect 28724 17196 28776 17202
rect 28724 17138 28776 17144
rect 28816 17196 28868 17202
rect 28920 17184 28948 17750
rect 29460 17740 29512 17746
rect 29460 17682 29512 17688
rect 29472 17338 29500 17682
rect 29840 17678 29868 20878
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29932 19854 29960 20334
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 30024 19666 30052 22510
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30392 22030 30420 22170
rect 30656 22160 30708 22166
rect 30656 22102 30708 22108
rect 30380 22024 30432 22030
rect 30208 21984 30380 22012
rect 30104 21684 30156 21690
rect 30104 21626 30156 21632
rect 30116 20466 30144 21626
rect 30208 21554 30236 21984
rect 30380 21966 30432 21972
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30196 21548 30248 21554
rect 30196 21490 30248 21496
rect 30484 21418 30512 21830
rect 30472 21412 30524 21418
rect 30472 21354 30524 21360
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 30116 19854 30144 20402
rect 30104 19848 30156 19854
rect 30104 19790 30156 19796
rect 30288 19780 30340 19786
rect 30288 19722 30340 19728
rect 29932 19638 30052 19666
rect 29932 17678 29960 19638
rect 30300 19514 30328 19722
rect 30472 19712 30524 19718
rect 30472 19654 30524 19660
rect 30484 19514 30512 19654
rect 30012 19508 30064 19514
rect 30012 19450 30064 19456
rect 30288 19508 30340 19514
rect 30288 19450 30340 19456
rect 30472 19508 30524 19514
rect 30472 19450 30524 19456
rect 30024 17814 30052 19450
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30484 19174 30512 19314
rect 30472 19168 30524 19174
rect 30472 19110 30524 19116
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30012 17808 30064 17814
rect 30012 17750 30064 17756
rect 29828 17672 29880 17678
rect 29828 17614 29880 17620
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 29460 17332 29512 17338
rect 29460 17274 29512 17280
rect 29092 17264 29144 17270
rect 29184 17264 29236 17270
rect 29092 17206 29144 17212
rect 29182 17232 29184 17241
rect 29236 17232 29238 17241
rect 29000 17196 29052 17202
rect 28920 17156 29000 17184
rect 28816 17138 28868 17144
rect 29000 17138 29052 17144
rect 28644 16658 28672 17138
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 28184 14618 28212 15506
rect 28724 15360 28776 15366
rect 28724 15302 28776 15308
rect 28356 15088 28408 15094
rect 28356 15030 28408 15036
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28172 14612 28224 14618
rect 28172 14554 28224 14560
rect 28172 14340 28224 14346
rect 28172 14282 28224 14288
rect 28184 13938 28212 14282
rect 28276 14074 28304 14962
rect 28368 14618 28396 15030
rect 28632 14952 28684 14958
rect 28632 14894 28684 14900
rect 28644 14822 28672 14894
rect 28632 14816 28684 14822
rect 28632 14758 28684 14764
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 28644 14074 28672 14758
rect 28736 14414 28764 15302
rect 28724 14408 28776 14414
rect 28724 14350 28776 14356
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28172 13932 28224 13938
rect 28172 13874 28224 13880
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28538 13832 28594 13841
rect 28092 13790 28212 13818
rect 27908 13382 28028 13410
rect 27804 11620 27856 11626
rect 27804 11562 27856 11568
rect 27528 11008 27580 11014
rect 27528 10950 27580 10956
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27540 10674 27568 10950
rect 27724 10826 27752 10950
rect 27632 10798 27752 10826
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27264 9654 27292 10542
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27160 9172 27212 9178
rect 27160 9114 27212 9120
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 26884 8968 26936 8974
rect 26884 8910 26936 8916
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 26528 7478 26556 8230
rect 26516 7472 26568 7478
rect 26516 7414 26568 7420
rect 26700 7472 26752 7478
rect 26804 7460 26832 8910
rect 26896 8634 26924 8910
rect 26988 8838 27016 8910
rect 27264 8838 27292 9590
rect 27356 9586 27384 10610
rect 27632 9586 27660 10798
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27724 10198 27752 10406
rect 27712 10192 27764 10198
rect 27712 10134 27764 10140
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 26976 8832 27028 8838
rect 26976 8774 27028 8780
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 26884 8628 26936 8634
rect 26884 8570 26936 8576
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26896 8090 26924 8366
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 26896 7478 26924 8026
rect 26988 7886 27016 8774
rect 27356 8090 27384 9522
rect 27712 9512 27764 9518
rect 27712 9454 27764 9460
rect 27724 8566 27752 9454
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 27172 7886 27200 8026
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 26752 7432 26832 7460
rect 26700 7414 26752 7420
rect 25596 7336 25648 7342
rect 25596 7278 25648 7284
rect 25608 7002 25636 7278
rect 26424 7268 26476 7274
rect 26424 7210 26476 7216
rect 25688 7200 25740 7206
rect 25688 7142 25740 7148
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25516 4622 25544 6734
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25608 6390 25636 6598
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25700 5710 25728 7142
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25700 4826 25728 4966
rect 26436 4826 26464 7210
rect 26804 6390 26832 7432
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 27172 7206 27200 7822
rect 27344 7744 27396 7750
rect 27344 7686 27396 7692
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27356 7546 27384 7686
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27252 7404 27304 7410
rect 27252 7346 27304 7352
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 27264 6934 27292 7346
rect 27252 6928 27304 6934
rect 27252 6870 27304 6876
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 26516 6384 26568 6390
rect 26516 6326 26568 6332
rect 26792 6384 26844 6390
rect 26792 6326 26844 6332
rect 26528 6118 26556 6326
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 25596 4820 25648 4826
rect 25596 4762 25648 4768
rect 25688 4820 25740 4826
rect 25688 4762 25740 4768
rect 25872 4820 25924 4826
rect 25872 4762 25924 4768
rect 26424 4820 26476 4826
rect 26424 4762 26476 4768
rect 25608 4622 25636 4762
rect 25504 4616 25556 4622
rect 25504 4558 25556 4564
rect 25596 4616 25648 4622
rect 25596 4558 25648 4564
rect 25516 4010 25544 4558
rect 25884 4214 25912 4762
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 25976 4078 26004 4558
rect 26436 4214 26464 4762
rect 27080 4690 27108 6734
rect 27068 4684 27120 4690
rect 27068 4626 27120 4632
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26516 4548 26568 4554
rect 26516 4490 26568 4496
rect 26528 4214 26556 4490
rect 26804 4282 26832 4558
rect 26884 4548 26936 4554
rect 26884 4490 26936 4496
rect 26792 4276 26844 4282
rect 26792 4218 26844 4224
rect 26424 4208 26476 4214
rect 26424 4150 26476 4156
rect 26516 4208 26568 4214
rect 26516 4150 26568 4156
rect 26896 4078 26924 4490
rect 27080 4282 27108 4626
rect 27068 4276 27120 4282
rect 27068 4218 27120 4224
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 27356 4010 27384 7346
rect 27448 5574 27476 7686
rect 27540 7002 27568 7686
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27632 6186 27660 8298
rect 27816 6934 27844 8978
rect 27804 6928 27856 6934
rect 27804 6870 27856 6876
rect 27908 6798 27936 13382
rect 27988 12300 28040 12306
rect 27988 12242 28040 12248
rect 28000 6934 28028 12242
rect 28078 11112 28134 11121
rect 28184 11098 28212 13790
rect 28538 13767 28540 13776
rect 28592 13767 28594 13776
rect 28540 13738 28592 13744
rect 28552 13326 28580 13738
rect 28644 13462 28672 13874
rect 28632 13456 28684 13462
rect 28632 13398 28684 13404
rect 28448 13320 28500 13326
rect 28446 13288 28448 13297
rect 28540 13320 28592 13326
rect 28500 13288 28502 13297
rect 28540 13262 28592 13268
rect 28446 13223 28502 13232
rect 28134 11070 28212 11098
rect 28078 11047 28134 11056
rect 28460 10674 28488 13223
rect 28552 10674 28580 13262
rect 28644 12986 28672 13398
rect 28632 12980 28684 12986
rect 28632 12922 28684 12928
rect 28828 12442 28856 17138
rect 29104 16980 29132 17206
rect 29182 17167 29238 17176
rect 29184 16992 29236 16998
rect 29104 16952 29184 16980
rect 29184 16934 29236 16940
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 29104 15502 29132 16050
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 28908 15428 28960 15434
rect 28908 15370 28960 15376
rect 28920 12918 28948 15370
rect 29104 15026 29132 15438
rect 29092 15020 29144 15026
rect 29092 14962 29144 14968
rect 29000 13320 29052 13326
rect 29052 13280 29132 13308
rect 29000 13262 29052 13268
rect 29000 13184 29052 13190
rect 28998 13152 29000 13161
rect 29052 13152 29054 13161
rect 28998 13087 29054 13096
rect 28998 13016 29054 13025
rect 28998 12951 29054 12960
rect 28908 12912 28960 12918
rect 28908 12854 28960 12860
rect 28816 12436 28868 12442
rect 28920 12434 28948 12854
rect 29012 12782 29040 12951
rect 29104 12850 29132 13280
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 28920 12406 29040 12434
rect 28816 12378 28868 12384
rect 29012 12374 29040 12406
rect 29000 12368 29052 12374
rect 29000 12310 29052 12316
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 28920 11898 28948 12174
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 28908 11892 28960 11898
rect 28908 11834 28960 11840
rect 28644 11286 28672 11834
rect 29104 11762 29132 12786
rect 29092 11756 29144 11762
rect 29092 11698 29144 11704
rect 28724 11552 28776 11558
rect 28724 11494 28776 11500
rect 28632 11280 28684 11286
rect 28632 11222 28684 11228
rect 28736 11098 28764 11494
rect 28644 11070 28764 11098
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 28460 10062 28488 10610
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28552 9722 28580 10610
rect 28644 10538 28672 11070
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28632 10532 28684 10538
rect 28632 10474 28684 10480
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28448 8968 28500 8974
rect 28552 8956 28580 9454
rect 28500 8928 28580 8956
rect 28448 8910 28500 8916
rect 28172 8628 28224 8634
rect 28224 8588 28488 8616
rect 28172 8570 28224 8576
rect 28356 8492 28408 8498
rect 28276 8452 28356 8480
rect 28276 8294 28304 8452
rect 28356 8434 28408 8440
rect 28264 8288 28316 8294
rect 28264 8230 28316 8236
rect 28356 8288 28408 8294
rect 28356 8230 28408 8236
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 28184 7478 28212 7822
rect 28172 7472 28224 7478
rect 28172 7414 28224 7420
rect 28276 7002 28304 8230
rect 28368 7954 28396 8230
rect 28460 7954 28488 8588
rect 28356 7948 28408 7954
rect 28356 7890 28408 7896
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28552 7818 28580 8928
rect 28644 8294 28672 10474
rect 28736 10062 28764 10610
rect 28724 10056 28776 10062
rect 29092 10056 29144 10062
rect 28724 9998 28776 10004
rect 29012 10004 29092 10010
rect 29012 9998 29144 10004
rect 29012 9982 29132 9998
rect 28908 9920 28960 9926
rect 28908 9862 28960 9868
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 28736 8906 28764 9114
rect 28828 8974 28856 9318
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28724 8900 28776 8906
rect 28724 8842 28776 8848
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28736 8090 28764 8434
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 28828 7886 28856 8434
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 28540 7812 28592 7818
rect 28540 7754 28592 7760
rect 28448 7404 28500 7410
rect 28448 7346 28500 7352
rect 28264 6996 28316 7002
rect 28264 6938 28316 6944
rect 27988 6928 28040 6934
rect 27988 6870 28040 6876
rect 28460 6798 28488 7346
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28356 6792 28408 6798
rect 28356 6734 28408 6740
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 27896 6248 27948 6254
rect 27948 6208 28120 6236
rect 27896 6190 27948 6196
rect 27620 6180 27672 6186
rect 27620 6122 27672 6128
rect 27632 5710 27660 6122
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 27620 5704 27672 5710
rect 27620 5646 27672 5652
rect 27436 5568 27488 5574
rect 27436 5510 27488 5516
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27436 4548 27488 4554
rect 27436 4490 27488 4496
rect 27448 4282 27476 4490
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 27724 4214 27752 4762
rect 27896 4480 27948 4486
rect 27896 4422 27948 4428
rect 27908 4282 27936 4422
rect 27896 4276 27948 4282
rect 27896 4218 27948 4224
rect 27712 4208 27764 4214
rect 27712 4150 27764 4156
rect 28000 4146 28028 5782
rect 28092 5710 28120 6208
rect 28184 5914 28212 6734
rect 28368 5914 28396 6734
rect 28460 6458 28488 6734
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28448 6452 28500 6458
rect 28448 6394 28500 6400
rect 28448 6316 28500 6322
rect 28448 6258 28500 6264
rect 28172 5908 28224 5914
rect 28172 5850 28224 5856
rect 28356 5908 28408 5914
rect 28356 5850 28408 5856
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 28092 4758 28120 5646
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 28184 5098 28212 5306
rect 28172 5092 28224 5098
rect 28172 5034 28224 5040
rect 28080 4752 28132 4758
rect 28080 4694 28132 4700
rect 28080 4276 28132 4282
rect 28080 4218 28132 4224
rect 28092 4185 28120 4218
rect 28078 4176 28134 4185
rect 27988 4140 28040 4146
rect 28184 4146 28212 5034
rect 28460 4826 28488 6258
rect 28448 4820 28500 4826
rect 28448 4762 28500 4768
rect 28540 4684 28592 4690
rect 28540 4626 28592 4632
rect 28552 4282 28580 4626
rect 28540 4276 28592 4282
rect 28540 4218 28592 4224
rect 28078 4111 28134 4120
rect 28172 4140 28224 4146
rect 27988 4082 28040 4088
rect 28172 4082 28224 4088
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 27344 4004 27396 4010
rect 27344 3946 27396 3952
rect 28644 3942 28672 6598
rect 28920 6390 28948 9862
rect 29012 9586 29040 9982
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 29104 9042 29132 9862
rect 29092 9036 29144 9042
rect 29092 8978 29144 8984
rect 29196 8922 29224 16934
rect 29368 16176 29420 16182
rect 29368 16118 29420 16124
rect 29380 15026 29408 16118
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29828 15904 29880 15910
rect 29828 15846 29880 15852
rect 29564 15706 29592 15846
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29840 15502 29868 15846
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29368 13184 29420 13190
rect 29274 13152 29330 13161
rect 29368 13126 29420 13132
rect 29274 13087 29330 13096
rect 29288 12850 29316 13087
rect 29380 13025 29408 13126
rect 29366 13016 29422 13025
rect 29366 12951 29422 12960
rect 29564 12866 29592 14894
rect 29932 13802 29960 17614
rect 30024 14958 30052 17750
rect 30116 16250 30144 18158
rect 30208 17610 30236 18226
rect 30668 18086 30696 22102
rect 30760 19446 30788 24006
rect 30852 23866 30880 24006
rect 30840 23860 30892 23866
rect 30840 23802 30892 23808
rect 30944 22982 30972 31726
rect 31024 30048 31076 30054
rect 31024 29990 31076 29996
rect 31036 29714 31064 29990
rect 31024 29708 31076 29714
rect 31024 29650 31076 29656
rect 31024 29300 31076 29306
rect 31024 29242 31076 29248
rect 31036 27470 31064 29242
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 31024 26988 31076 26994
rect 31024 26930 31076 26936
rect 31036 26382 31064 26930
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 31036 24342 31064 26318
rect 31024 24336 31076 24342
rect 31024 24278 31076 24284
rect 31024 23792 31076 23798
rect 31024 23734 31076 23740
rect 30932 22976 30984 22982
rect 30932 22918 30984 22924
rect 31036 22506 31064 23734
rect 31128 23594 31156 31826
rect 31496 31754 31524 32166
rect 31680 31770 31708 33526
rect 32876 33522 32904 34138
rect 33140 33924 33192 33930
rect 33140 33866 33192 33872
rect 32864 33516 32916 33522
rect 32864 33458 32916 33464
rect 33152 32586 33180 33866
rect 33232 33856 33284 33862
rect 33232 33798 33284 33804
rect 33324 33856 33376 33862
rect 33324 33798 33376 33804
rect 33244 32910 33272 33798
rect 33336 33658 33364 33798
rect 33324 33652 33376 33658
rect 33324 33594 33376 33600
rect 33336 33318 33364 33594
rect 33324 33312 33376 33318
rect 33324 33254 33376 33260
rect 33428 32978 33456 34496
rect 33416 32972 33468 32978
rect 33416 32914 33468 32920
rect 33232 32904 33284 32910
rect 33232 32846 33284 32852
rect 32496 32564 32548 32570
rect 32496 32506 32548 32512
rect 33152 32558 33272 32586
rect 32128 32224 32180 32230
rect 32128 32166 32180 32172
rect 32140 32026 32168 32166
rect 32508 32026 32536 32506
rect 32128 32020 32180 32026
rect 32128 31962 32180 31968
rect 32496 32020 32548 32026
rect 32496 31962 32548 31968
rect 31852 31884 31904 31890
rect 31852 31826 31904 31832
rect 31680 31754 31800 31770
rect 31496 31726 31616 31754
rect 31680 31748 31812 31754
rect 31680 31742 31760 31748
rect 31300 31476 31352 31482
rect 31300 31418 31352 31424
rect 31312 31346 31340 31418
rect 31588 31346 31616 31726
rect 31760 31690 31812 31696
rect 31772 31659 31800 31690
rect 31864 31482 31892 31826
rect 31852 31476 31904 31482
rect 31852 31418 31904 31424
rect 31300 31340 31352 31346
rect 31300 31282 31352 31288
rect 31576 31340 31628 31346
rect 31576 31282 31628 31288
rect 32312 31340 32364 31346
rect 32312 31282 32364 31288
rect 31312 29306 31340 31282
rect 32036 31136 32088 31142
rect 32036 31078 32088 31084
rect 31668 30048 31720 30054
rect 31668 29990 31720 29996
rect 31680 29306 31708 29990
rect 31760 29640 31812 29646
rect 31760 29582 31812 29588
rect 31300 29300 31352 29306
rect 31300 29242 31352 29248
rect 31668 29300 31720 29306
rect 31668 29242 31720 29248
rect 31772 29238 31800 29582
rect 31760 29232 31812 29238
rect 31760 29174 31812 29180
rect 31944 29232 31996 29238
rect 31944 29174 31996 29180
rect 31576 29164 31628 29170
rect 31576 29106 31628 29112
rect 31588 29073 31616 29106
rect 31574 29064 31630 29073
rect 31956 29034 31984 29174
rect 31574 28999 31630 29008
rect 31944 29028 31996 29034
rect 31944 28970 31996 28976
rect 31484 28960 31536 28966
rect 31484 28902 31536 28908
rect 31496 28558 31524 28902
rect 31484 28552 31536 28558
rect 31390 28520 31446 28529
rect 31484 28494 31536 28500
rect 31390 28455 31392 28464
rect 31444 28455 31446 28464
rect 31760 28484 31812 28490
rect 31392 28426 31444 28432
rect 31760 28426 31812 28432
rect 31208 27464 31260 27470
rect 31208 27406 31260 27412
rect 31220 26246 31248 27406
rect 31300 27396 31352 27402
rect 31300 27338 31352 27344
rect 31312 26858 31340 27338
rect 31300 26852 31352 26858
rect 31300 26794 31352 26800
rect 31404 26738 31432 28426
rect 31772 28218 31800 28426
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31312 26710 31432 26738
rect 31312 26314 31340 26710
rect 31392 26376 31444 26382
rect 31392 26318 31444 26324
rect 31300 26308 31352 26314
rect 31300 26250 31352 26256
rect 31208 26240 31260 26246
rect 31208 26182 31260 26188
rect 31312 26042 31340 26250
rect 31404 26042 31432 26318
rect 31760 26308 31812 26314
rect 31760 26250 31812 26256
rect 31772 26042 31800 26250
rect 31300 26036 31352 26042
rect 31300 25978 31352 25984
rect 31392 26036 31444 26042
rect 31392 25978 31444 25984
rect 31760 26036 31812 26042
rect 31760 25978 31812 25984
rect 31760 25696 31812 25702
rect 31760 25638 31812 25644
rect 31772 24886 31800 25638
rect 32048 25294 32076 31078
rect 32220 30592 32272 30598
rect 32220 30534 32272 30540
rect 32232 29646 32260 30534
rect 32220 29640 32272 29646
rect 32220 29582 32272 29588
rect 32324 29102 32352 31282
rect 32404 31136 32456 31142
rect 32404 31078 32456 31084
rect 32416 30190 32444 31078
rect 32496 30592 32548 30598
rect 32496 30534 32548 30540
rect 33048 30592 33100 30598
rect 33048 30534 33100 30540
rect 32508 30394 32536 30534
rect 32496 30388 32548 30394
rect 32496 30330 32548 30336
rect 32404 30184 32456 30190
rect 32404 30126 32456 30132
rect 32864 29572 32916 29578
rect 32864 29514 32916 29520
rect 32956 29572 33008 29578
rect 32956 29514 33008 29520
rect 32496 29504 32548 29510
rect 32496 29446 32548 29452
rect 32508 29238 32536 29446
rect 32496 29232 32548 29238
rect 32496 29174 32548 29180
rect 32312 29096 32364 29102
rect 32312 29038 32364 29044
rect 32772 29096 32824 29102
rect 32772 29038 32824 29044
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 32508 27674 32536 28018
rect 32784 28014 32812 29038
rect 32772 28008 32824 28014
rect 32772 27950 32824 27956
rect 32496 27668 32548 27674
rect 32496 27610 32548 27616
rect 32404 27464 32456 27470
rect 32404 27406 32456 27412
rect 32416 26042 32444 27406
rect 32588 26784 32640 26790
rect 32588 26726 32640 26732
rect 32600 26466 32628 26726
rect 32680 26512 32732 26518
rect 32600 26460 32680 26466
rect 32600 26454 32732 26460
rect 32600 26438 32720 26454
rect 32496 26240 32548 26246
rect 32496 26182 32548 26188
rect 32404 26036 32456 26042
rect 32404 25978 32456 25984
rect 32508 25974 32536 26182
rect 32600 26042 32628 26438
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32496 25968 32548 25974
rect 32496 25910 32548 25916
rect 32508 25702 32536 25910
rect 32784 25838 32812 27950
rect 32772 25832 32824 25838
rect 32772 25774 32824 25780
rect 32496 25696 32548 25702
rect 32496 25638 32548 25644
rect 32036 25288 32088 25294
rect 32036 25230 32088 25236
rect 32496 25288 32548 25294
rect 32496 25230 32548 25236
rect 32232 24942 32444 24970
rect 31760 24880 31812 24886
rect 31760 24822 31812 24828
rect 32128 24812 32180 24818
rect 32232 24800 32260 24942
rect 32416 24818 32444 24942
rect 32508 24886 32536 25230
rect 32496 24880 32548 24886
rect 32496 24822 32548 24828
rect 32180 24772 32260 24800
rect 32312 24812 32364 24818
rect 32128 24754 32180 24760
rect 32312 24754 32364 24760
rect 32404 24812 32456 24818
rect 32404 24754 32456 24760
rect 32036 24676 32088 24682
rect 32036 24618 32088 24624
rect 31484 24268 31536 24274
rect 31484 24210 31536 24216
rect 31208 24064 31260 24070
rect 31208 24006 31260 24012
rect 31116 23588 31168 23594
rect 31116 23530 31168 23536
rect 31220 23118 31248 24006
rect 31496 23662 31524 24210
rect 32048 24206 32076 24618
rect 32140 24342 32168 24754
rect 32220 24608 32272 24614
rect 32220 24550 32272 24556
rect 32128 24336 32180 24342
rect 32128 24278 32180 24284
rect 32036 24200 32088 24206
rect 32036 24142 32088 24148
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 31852 24064 31904 24070
rect 31852 24006 31904 24012
rect 31484 23656 31536 23662
rect 31484 23598 31536 23604
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31220 22778 31248 23054
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 31760 22568 31812 22574
rect 31760 22510 31812 22516
rect 31024 22500 31076 22506
rect 31024 22442 31076 22448
rect 31484 22432 31536 22438
rect 31484 22374 31536 22380
rect 31496 22234 31524 22374
rect 31484 22228 31536 22234
rect 31484 22170 31536 22176
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31220 21690 31248 21966
rect 31300 21888 31352 21894
rect 31300 21830 31352 21836
rect 31208 21684 31260 21690
rect 31208 21626 31260 21632
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30840 19780 30892 19786
rect 30840 19722 30892 19728
rect 30748 19440 30800 19446
rect 30748 19382 30800 19388
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30196 17604 30248 17610
rect 30196 17546 30248 17552
rect 30104 16244 30156 16250
rect 30104 16186 30156 16192
rect 30104 15360 30156 15366
rect 30104 15302 30156 15308
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 29920 13796 29972 13802
rect 29920 13738 29972 13744
rect 29828 13456 29880 13462
rect 29828 13398 29880 13404
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29276 12844 29328 12850
rect 29276 12786 29328 12792
rect 29380 12838 29592 12866
rect 29276 12096 29328 12102
rect 29276 12038 29328 12044
rect 29288 11898 29316 12038
rect 29276 11892 29328 11898
rect 29276 11834 29328 11840
rect 29380 10470 29408 12838
rect 29656 12714 29684 13194
rect 29840 12714 29868 13398
rect 29644 12708 29696 12714
rect 29828 12708 29880 12714
rect 29644 12650 29696 12656
rect 29748 12668 29828 12696
rect 29552 12640 29604 12646
rect 29472 12588 29552 12594
rect 29472 12582 29604 12588
rect 29472 12566 29592 12582
rect 29472 12442 29500 12566
rect 29460 12436 29512 12442
rect 29460 12378 29512 12384
rect 29552 12436 29604 12442
rect 29552 12378 29604 12384
rect 29472 12238 29500 12378
rect 29460 12232 29512 12238
rect 29460 12174 29512 12180
rect 29564 11762 29592 12378
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 29748 11354 29776 12668
rect 29828 12650 29880 12656
rect 30024 12434 30052 14894
rect 30116 13530 30144 15302
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 30116 13258 30144 13466
rect 30104 13252 30156 13258
rect 30104 13194 30156 13200
rect 30208 12442 30236 17546
rect 30392 16454 30420 17818
rect 30484 17678 30512 18022
rect 30472 17672 30524 17678
rect 30472 17614 30524 17620
rect 30484 17270 30512 17614
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 30288 16108 30340 16114
rect 30288 16050 30340 16056
rect 30300 14890 30328 16050
rect 30380 15972 30432 15978
rect 30380 15914 30432 15920
rect 30748 15972 30800 15978
rect 30748 15914 30800 15920
rect 30392 15638 30420 15914
rect 30656 15700 30708 15706
rect 30656 15642 30708 15648
rect 30380 15632 30432 15638
rect 30380 15574 30432 15580
rect 30668 15094 30696 15642
rect 30760 15570 30788 15914
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30656 15088 30708 15094
rect 30656 15030 30708 15036
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30472 14272 30524 14278
rect 30472 14214 30524 14220
rect 30380 13252 30432 13258
rect 30380 13194 30432 13200
rect 30392 12646 30420 13194
rect 30484 13190 30512 14214
rect 30576 13870 30604 14962
rect 30656 14544 30708 14550
rect 30656 14486 30708 14492
rect 30746 14512 30802 14521
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30576 12850 30604 13806
rect 30668 13326 30696 14486
rect 30852 14498 30880 19722
rect 30944 19310 30972 21286
rect 31312 20942 31340 21830
rect 31496 21554 31524 22170
rect 31576 22160 31628 22166
rect 31628 22137 31708 22148
rect 31628 22128 31722 22137
rect 31628 22120 31666 22128
rect 31576 22102 31628 22108
rect 31666 22063 31722 22072
rect 31576 22024 31628 22030
rect 31772 21978 31800 22510
rect 31864 22030 31892 24006
rect 31944 22160 31996 22166
rect 32048 22148 32076 24142
rect 32140 23866 32168 24142
rect 32232 24070 32260 24550
rect 32324 24290 32352 24754
rect 32508 24426 32536 24822
rect 32588 24676 32640 24682
rect 32588 24618 32640 24624
rect 32416 24398 32536 24426
rect 32416 24290 32444 24398
rect 32324 24262 32444 24290
rect 32496 24336 32548 24342
rect 32496 24278 32548 24284
rect 32220 24064 32272 24070
rect 32220 24006 32272 24012
rect 32324 23866 32352 24262
rect 32404 24200 32456 24206
rect 32404 24142 32456 24148
rect 32416 23866 32444 24142
rect 32128 23860 32180 23866
rect 32128 23802 32180 23808
rect 32312 23860 32364 23866
rect 32312 23802 32364 23808
rect 32404 23860 32456 23866
rect 32404 23802 32456 23808
rect 32140 23118 32168 23802
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 32140 22710 32168 23054
rect 32312 22976 32364 22982
rect 32312 22918 32364 22924
rect 32324 22778 32352 22918
rect 32312 22772 32364 22778
rect 32312 22714 32364 22720
rect 32128 22704 32180 22710
rect 32128 22646 32180 22652
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 31996 22120 32076 22148
rect 31944 22102 31996 22108
rect 32048 22030 32076 22120
rect 32140 22030 32168 22374
rect 32324 22166 32352 22578
rect 32312 22160 32364 22166
rect 32312 22102 32364 22108
rect 31628 21972 31800 21978
rect 31576 21966 31800 21972
rect 31852 22024 31904 22030
rect 31852 21966 31904 21972
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31588 21950 31800 21966
rect 32048 21554 32076 21966
rect 32140 21690 32168 21966
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 32324 21554 32352 22102
rect 32416 22030 32444 22578
rect 32508 22094 32536 24278
rect 32600 24206 32628 24618
rect 32588 24200 32640 24206
rect 32588 24142 32640 24148
rect 32784 23526 32812 25774
rect 32876 24970 32904 29514
rect 32968 29306 32996 29514
rect 32956 29300 33008 29306
rect 32956 29242 33008 29248
rect 33060 29073 33088 30534
rect 33152 30326 33180 32558
rect 33244 32502 33272 32558
rect 33232 32496 33284 32502
rect 33232 32438 33284 32444
rect 33140 30320 33192 30326
rect 33140 30262 33192 30268
rect 33046 29064 33102 29073
rect 33046 28999 33102 29008
rect 33060 28558 33088 28999
rect 33152 28626 33180 30262
rect 33428 29102 33456 32914
rect 33520 31906 33548 35686
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 33692 35148 33744 35154
rect 33692 35090 33744 35096
rect 33704 34066 33732 35090
rect 37556 34604 37608 34610
rect 37556 34546 37608 34552
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 33692 34060 33744 34066
rect 33692 34002 33744 34008
rect 33704 33946 33732 34002
rect 33704 33918 33824 33946
rect 33600 33584 33652 33590
rect 33600 33526 33652 33532
rect 33612 32026 33640 33526
rect 33692 32768 33744 32774
rect 33692 32710 33744 32716
rect 33704 32366 33732 32710
rect 33692 32360 33744 32366
rect 33692 32302 33744 32308
rect 33600 32020 33652 32026
rect 33600 31962 33652 31968
rect 33520 31890 33640 31906
rect 33520 31884 33652 31890
rect 33520 31878 33600 31884
rect 33600 31826 33652 31832
rect 33416 29096 33468 29102
rect 33416 29038 33468 29044
rect 33140 28620 33192 28626
rect 33140 28562 33192 28568
rect 33048 28552 33100 28558
rect 33048 28494 33100 28500
rect 33152 28422 33180 28562
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33140 28416 33192 28422
rect 33140 28358 33192 28364
rect 33232 28416 33284 28422
rect 33232 28358 33284 28364
rect 33244 28082 33272 28358
rect 33520 28082 33548 28426
rect 33232 28076 33284 28082
rect 33232 28018 33284 28024
rect 33508 28076 33560 28082
rect 33508 28018 33560 28024
rect 32956 25832 33008 25838
rect 32956 25774 33008 25780
rect 32968 25430 32996 25774
rect 33508 25696 33560 25702
rect 33508 25638 33560 25644
rect 33520 25498 33548 25638
rect 33508 25492 33560 25498
rect 33508 25434 33560 25440
rect 32956 25424 33008 25430
rect 32956 25366 33008 25372
rect 32876 24942 32996 24970
rect 32968 24818 32996 24942
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 32876 24410 32904 24754
rect 32864 24404 32916 24410
rect 32864 24346 32916 24352
rect 32968 24206 32996 24754
rect 32956 24200 33008 24206
rect 32956 24142 33008 24148
rect 32956 24064 33008 24070
rect 32956 24006 33008 24012
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 32968 22642 32996 24006
rect 33232 23588 33284 23594
rect 33232 23530 33284 23536
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 32680 22160 32732 22166
rect 32678 22128 32680 22137
rect 32732 22128 32734 22137
rect 32508 22066 32628 22094
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32416 21690 32444 21966
rect 32496 21888 32548 21894
rect 32496 21830 32548 21836
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31852 21548 31904 21554
rect 31852 21490 31904 21496
rect 32036 21548 32088 21554
rect 32036 21490 32088 21496
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31116 20800 31168 20806
rect 31116 20742 31168 20748
rect 30932 19304 30984 19310
rect 30932 19246 30984 19252
rect 31128 18222 31156 20742
rect 31208 19440 31260 19446
rect 31208 19382 31260 19388
rect 31220 18766 31248 19382
rect 31300 19168 31352 19174
rect 31300 19110 31352 19116
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31022 18048 31078 18057
rect 31022 17983 31078 17992
rect 30932 14816 30984 14822
rect 30932 14758 30984 14764
rect 30802 14470 30880 14498
rect 30746 14447 30802 14456
rect 30852 14414 30880 14470
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30944 14346 30972 14758
rect 30748 14340 30800 14346
rect 30748 14282 30800 14288
rect 30932 14340 30984 14346
rect 30932 14282 30984 14288
rect 30760 14074 30788 14282
rect 30748 14068 30800 14074
rect 30748 14010 30800 14016
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30840 13184 30892 13190
rect 30840 13126 30892 13132
rect 30564 12844 30616 12850
rect 30564 12786 30616 12792
rect 30472 12708 30524 12714
rect 30472 12650 30524 12656
rect 30380 12640 30432 12646
rect 30380 12582 30432 12588
rect 30196 12436 30248 12442
rect 30024 12406 30144 12434
rect 30012 12368 30064 12374
rect 30012 12310 30064 12316
rect 30116 12322 30144 12406
rect 30196 12378 30248 12384
rect 29828 12096 29880 12102
rect 29828 12038 29880 12044
rect 29840 11898 29868 12038
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 30024 11694 30052 12310
rect 30116 12294 30328 12322
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30104 12096 30156 12102
rect 30104 12038 30156 12044
rect 30012 11688 30064 11694
rect 30012 11630 30064 11636
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29828 11008 29880 11014
rect 29828 10950 29880 10956
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 29644 10464 29696 10470
rect 29644 10406 29696 10412
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 29380 9586 29408 9998
rect 29368 9580 29420 9586
rect 29368 9522 29420 9528
rect 29276 9376 29328 9382
rect 29276 9318 29328 9324
rect 29288 9178 29316 9318
rect 29276 9172 29328 9178
rect 29276 9114 29328 9120
rect 29104 8894 29224 8922
rect 29104 7342 29132 8894
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 29196 6798 29224 8774
rect 29380 8566 29408 9522
rect 29550 9480 29606 9489
rect 29550 9415 29552 9424
rect 29604 9415 29606 9424
rect 29552 9386 29604 9392
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29564 8634 29592 8910
rect 29552 8628 29604 8634
rect 29552 8570 29604 8576
rect 29368 8560 29420 8566
rect 29368 8502 29420 8508
rect 29368 8356 29420 8362
rect 29368 8298 29420 8304
rect 29380 7410 29408 8298
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29564 7886 29592 8230
rect 29552 7880 29604 7886
rect 29552 7822 29604 7828
rect 29276 7404 29328 7410
rect 29276 7346 29328 7352
rect 29368 7404 29420 7410
rect 29420 7364 29500 7392
rect 29368 7346 29420 7352
rect 29288 6866 29316 7346
rect 29368 7200 29420 7206
rect 29368 7142 29420 7148
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 28908 6384 28960 6390
rect 28908 6326 28960 6332
rect 28724 6180 28776 6186
rect 28724 6122 28776 6128
rect 28736 4758 28764 6122
rect 28724 4752 28776 4758
rect 28724 4694 28776 4700
rect 29288 4690 29316 6802
rect 29380 5914 29408 7142
rect 29368 5908 29420 5914
rect 29368 5850 29420 5856
rect 29472 5846 29500 7364
rect 29656 6254 29684 10406
rect 29840 10062 29868 10950
rect 29932 10198 29960 11086
rect 29920 10192 29972 10198
rect 29920 10134 29972 10140
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29932 8922 29960 10134
rect 30116 8974 30144 12038
rect 30208 9654 30236 12174
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 30104 8968 30156 8974
rect 29932 8894 30052 8922
rect 30104 8910 30156 8916
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 29932 8634 29960 8774
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 30024 8498 30052 8894
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30024 8090 30052 8434
rect 30012 8084 30064 8090
rect 30012 8026 30064 8032
rect 30300 7886 30328 12294
rect 30392 10010 30420 12582
rect 30484 12374 30512 12650
rect 30472 12368 30524 12374
rect 30472 12310 30524 12316
rect 30576 12238 30604 12786
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30668 11694 30696 12038
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 30484 10674 30512 11494
rect 30576 11150 30604 11630
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30576 10810 30604 11086
rect 30564 10804 30616 10810
rect 30564 10746 30616 10752
rect 30472 10668 30524 10674
rect 30472 10610 30524 10616
rect 30472 10464 30524 10470
rect 30472 10406 30524 10412
rect 30484 10198 30512 10406
rect 30472 10192 30524 10198
rect 30472 10134 30524 10140
rect 30472 10056 30524 10062
rect 30392 10004 30472 10010
rect 30392 9998 30524 10004
rect 30576 10010 30604 10746
rect 30748 10668 30800 10674
rect 30748 10610 30800 10616
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30668 10198 30696 10542
rect 30656 10192 30708 10198
rect 30656 10134 30708 10140
rect 30656 10056 30708 10062
rect 30576 10004 30656 10010
rect 30576 9998 30708 10004
rect 30392 9982 30512 9998
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30392 8974 30420 9862
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 30300 7410 30328 7822
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 29920 6996 29972 7002
rect 29920 6938 29972 6944
rect 29644 6248 29696 6254
rect 29644 6190 29696 6196
rect 29932 5846 29960 6938
rect 30484 6866 30512 9982
rect 30576 9982 30696 9998
rect 30576 9722 30604 9982
rect 30564 9716 30616 9722
rect 30564 9658 30616 9664
rect 30656 9512 30708 9518
rect 30656 9454 30708 9460
rect 30668 8634 30696 9454
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30564 8424 30616 8430
rect 30564 8366 30616 8372
rect 30576 8022 30604 8366
rect 30564 8016 30616 8022
rect 30564 7958 30616 7964
rect 30576 7886 30604 7958
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30656 7880 30708 7886
rect 30656 7822 30708 7828
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30576 6798 30604 7822
rect 30668 6798 30696 7822
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30656 6792 30708 6798
rect 30656 6734 30708 6740
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 30116 5914 30144 6258
rect 30104 5908 30156 5914
rect 30104 5850 30156 5856
rect 29460 5840 29512 5846
rect 29460 5782 29512 5788
rect 29920 5840 29972 5846
rect 29920 5782 29972 5788
rect 30012 5840 30064 5846
rect 30012 5782 30064 5788
rect 29472 5710 29500 5782
rect 29932 5710 29960 5782
rect 29460 5704 29512 5710
rect 29460 5646 29512 5652
rect 29920 5704 29972 5710
rect 29920 5646 29972 5652
rect 29736 5568 29788 5574
rect 29736 5510 29788 5516
rect 29748 5234 29776 5510
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 29736 5228 29788 5234
rect 29736 5170 29788 5176
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 29472 4826 29500 4966
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29276 4684 29328 4690
rect 29276 4626 29328 4632
rect 29564 4146 29592 5170
rect 29828 5160 29880 5166
rect 29828 5102 29880 5108
rect 29840 5030 29868 5102
rect 29828 5024 29880 5030
rect 29828 4966 29880 4972
rect 29932 4622 29960 5646
rect 30024 4826 30052 5782
rect 30392 5574 30420 6258
rect 30760 5794 30788 10610
rect 30852 10130 30880 13126
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30852 9926 30880 10066
rect 30840 9920 30892 9926
rect 30840 9862 30892 9868
rect 30932 9920 30984 9926
rect 30932 9862 30984 9868
rect 30944 9586 30972 9862
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 30932 9580 30984 9586
rect 30932 9522 30984 9528
rect 30852 9178 30880 9522
rect 30840 9172 30892 9178
rect 30840 9114 30892 9120
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30852 8362 30880 8774
rect 30840 8356 30892 8362
rect 30840 8298 30892 8304
rect 30852 7886 30880 8298
rect 30840 7880 30892 7886
rect 30840 7822 30892 7828
rect 31036 7478 31064 17983
rect 31208 17876 31260 17882
rect 31208 17818 31260 17824
rect 31220 17202 31248 17818
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31220 11898 31248 17138
rect 31312 14346 31340 19110
rect 31760 18896 31812 18902
rect 31760 18838 31812 18844
rect 31772 18222 31800 18838
rect 31760 18216 31812 18222
rect 31760 18158 31812 18164
rect 31772 17746 31800 18158
rect 31392 17740 31444 17746
rect 31392 17682 31444 17688
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 31404 17338 31432 17682
rect 31576 17672 31628 17678
rect 31576 17614 31628 17620
rect 31668 17672 31720 17678
rect 31668 17614 31720 17620
rect 31588 17338 31616 17614
rect 31680 17542 31708 17614
rect 31668 17536 31720 17542
rect 31668 17478 31720 17484
rect 31680 17338 31708 17478
rect 31392 17332 31444 17338
rect 31392 17274 31444 17280
rect 31576 17332 31628 17338
rect 31576 17274 31628 17280
rect 31668 17332 31720 17338
rect 31668 17274 31720 17280
rect 31588 17202 31616 17274
rect 31772 17202 31800 17682
rect 31864 17678 31892 21490
rect 32508 21010 32536 21830
rect 32600 21554 32628 22066
rect 32678 22063 32734 22072
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 32772 21888 32824 21894
rect 32772 21830 32824 21836
rect 32784 21554 32812 21830
rect 32876 21690 32904 21966
rect 32864 21684 32916 21690
rect 32864 21626 32916 21632
rect 33152 21554 33180 21966
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 33140 21548 33192 21554
rect 33140 21490 33192 21496
rect 32496 21004 32548 21010
rect 32496 20946 32548 20952
rect 33048 20800 33100 20806
rect 33048 20742 33100 20748
rect 31944 19372 31996 19378
rect 31944 19314 31996 19320
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 31956 18698 31984 19314
rect 32220 19304 32272 19310
rect 32220 19246 32272 19252
rect 32232 18766 32260 19246
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 31944 18692 31996 18698
rect 31944 18634 31996 18640
rect 32416 18630 32444 19314
rect 32600 18766 32628 19314
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32956 18692 33008 18698
rect 32876 18652 32956 18680
rect 32036 18624 32088 18630
rect 32036 18566 32088 18572
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32404 18624 32456 18630
rect 32404 18566 32456 18572
rect 32772 18624 32824 18630
rect 32772 18566 32824 18572
rect 32048 18426 32076 18566
rect 32036 18420 32088 18426
rect 32036 18362 32088 18368
rect 32220 18148 32272 18154
rect 32220 18090 32272 18096
rect 32232 17814 32260 18090
rect 32324 17882 32352 18566
rect 32416 18222 32444 18566
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32784 18086 32812 18566
rect 32772 18080 32824 18086
rect 32772 18022 32824 18028
rect 32312 17876 32364 17882
rect 32312 17818 32364 17824
rect 32220 17808 32272 17814
rect 32220 17750 32272 17756
rect 31852 17672 31904 17678
rect 31852 17614 31904 17620
rect 32496 17672 32548 17678
rect 32496 17614 32548 17620
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31760 17196 31812 17202
rect 31760 17138 31812 17144
rect 32404 17060 32456 17066
rect 32404 17002 32456 17008
rect 32416 16794 32444 17002
rect 32404 16788 32456 16794
rect 32404 16730 32456 16736
rect 32128 16584 32180 16590
rect 32128 16526 32180 16532
rect 32036 15564 32088 15570
rect 32036 15506 32088 15512
rect 31760 15020 31812 15026
rect 31760 14962 31812 14968
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 31300 14340 31352 14346
rect 31300 14282 31352 14288
rect 31312 12481 31340 14282
rect 31496 12986 31524 14350
rect 31588 14074 31616 14350
rect 31576 14068 31628 14074
rect 31576 14010 31628 14016
rect 31772 13870 31800 14962
rect 32048 14618 32076 15506
rect 32036 14612 32088 14618
rect 32036 14554 32088 14560
rect 31852 13932 31904 13938
rect 31852 13874 31904 13880
rect 31760 13864 31812 13870
rect 31760 13806 31812 13812
rect 31668 13728 31720 13734
rect 31864 13716 31892 13874
rect 31668 13670 31720 13676
rect 31772 13688 31892 13716
rect 31680 13326 31708 13670
rect 31772 13394 31800 13688
rect 32140 13530 32168 16526
rect 32416 15502 32444 16730
rect 32508 16658 32536 17614
rect 32784 17610 32812 18022
rect 32876 17678 32904 18652
rect 32956 18634 33008 18640
rect 33060 17728 33088 20742
rect 33244 19854 33272 23530
rect 33612 22982 33640 31826
rect 33796 30190 33824 33918
rect 34612 33924 34664 33930
rect 34612 33866 34664 33872
rect 34152 33856 34204 33862
rect 34152 33798 34204 33804
rect 34164 33522 34192 33798
rect 34152 33516 34204 33522
rect 34152 33458 34204 33464
rect 34624 32842 34652 33866
rect 37568 33658 37596 34546
rect 37924 34536 37976 34542
rect 37924 34478 37976 34484
rect 37936 34105 37964 34478
rect 37922 34096 37978 34105
rect 37922 34031 37978 34040
rect 37556 33652 37608 33658
rect 37556 33594 37608 33600
rect 37556 33516 37608 33522
rect 37556 33458 37608 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 37568 33114 37596 33458
rect 37556 33108 37608 33114
rect 37556 33050 37608 33056
rect 34796 32904 34848 32910
rect 34716 32864 34796 32892
rect 33968 32836 34020 32842
rect 33968 32778 34020 32784
rect 34612 32836 34664 32842
rect 34612 32778 34664 32784
rect 33980 32434 34008 32778
rect 33968 32428 34020 32434
rect 33968 32370 34020 32376
rect 34244 32360 34296 32366
rect 34244 32302 34296 32308
rect 33968 32224 34020 32230
rect 33968 32166 34020 32172
rect 34152 32224 34204 32230
rect 34152 32166 34204 32172
rect 33980 31890 34008 32166
rect 34164 32026 34192 32166
rect 34256 32026 34284 32302
rect 34152 32020 34204 32026
rect 34152 31962 34204 31968
rect 34244 32020 34296 32026
rect 34244 31962 34296 31968
rect 33968 31884 34020 31890
rect 33968 31826 34020 31832
rect 33980 31754 34008 31826
rect 33980 31726 34284 31754
rect 34256 30274 34284 31726
rect 34624 31346 34652 32778
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 34336 30728 34388 30734
rect 34336 30670 34388 30676
rect 34348 30394 34376 30670
rect 34520 30592 34572 30598
rect 34520 30534 34572 30540
rect 34336 30388 34388 30394
rect 34336 30330 34388 30336
rect 34532 30326 34560 30534
rect 34520 30320 34572 30326
rect 34256 30246 34376 30274
rect 34520 30262 34572 30268
rect 33784 30184 33836 30190
rect 33784 30126 33836 30132
rect 34244 30184 34296 30190
rect 34244 30126 34296 30132
rect 33692 28756 33744 28762
rect 33692 28698 33744 28704
rect 33704 27674 33732 28698
rect 33796 28014 33824 30126
rect 34256 29510 34284 30126
rect 34348 29714 34376 30246
rect 34532 29850 34560 30262
rect 34520 29844 34572 29850
rect 34520 29786 34572 29792
rect 34336 29708 34388 29714
rect 34336 29650 34388 29656
rect 34244 29504 34296 29510
rect 34244 29446 34296 29452
rect 34244 28416 34296 28422
rect 34244 28358 34296 28364
rect 34256 28218 34284 28358
rect 34244 28212 34296 28218
rect 34244 28154 34296 28160
rect 33968 28144 34020 28150
rect 33968 28086 34020 28092
rect 33784 28008 33836 28014
rect 33784 27950 33836 27956
rect 33692 27668 33744 27674
rect 33692 27610 33744 27616
rect 33796 27334 33824 27950
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 33784 26444 33836 26450
rect 33784 26386 33836 26392
rect 33690 26344 33746 26353
rect 33690 26279 33692 26288
rect 33744 26279 33746 26288
rect 33692 26250 33744 26256
rect 33796 25838 33824 26386
rect 33980 26042 34008 28086
rect 34348 27614 34376 29650
rect 34716 29646 34744 32864
rect 34796 32846 34848 32852
rect 34796 32768 34848 32774
rect 34796 32710 34848 32716
rect 35072 32768 35124 32774
rect 35072 32710 35124 32716
rect 34808 32570 34836 32710
rect 35084 32570 35112 32710
rect 34796 32564 34848 32570
rect 34796 32506 34848 32512
rect 35072 32564 35124 32570
rect 35072 32506 35124 32512
rect 36636 32360 36688 32366
rect 36636 32302 36688 32308
rect 35900 32224 35952 32230
rect 35900 32166 35952 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35912 31754 35940 32166
rect 35912 31726 36032 31754
rect 34796 31136 34848 31142
rect 34796 31078 34848 31084
rect 34808 30938 34836 31078
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30932 34848 30938
rect 34796 30874 34848 30880
rect 36004 30666 36032 31726
rect 36648 31686 36676 32302
rect 36636 31680 36688 31686
rect 36636 31622 36688 31628
rect 35992 30660 36044 30666
rect 35992 30602 36044 30608
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34716 29306 34744 29582
rect 34796 29504 34848 29510
rect 34796 29446 34848 29452
rect 34980 29504 35032 29510
rect 34980 29446 35032 29452
rect 36360 29504 36412 29510
rect 36360 29446 36412 29452
rect 34808 29306 34836 29446
rect 34704 29300 34756 29306
rect 34704 29242 34756 29248
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 34520 28416 34572 28422
rect 34520 28358 34572 28364
rect 34532 28218 34560 28358
rect 34520 28212 34572 28218
rect 34520 28154 34572 28160
rect 34256 27586 34376 27614
rect 34716 27606 34744 29242
rect 34888 29232 34940 29238
rect 34808 29180 34888 29186
rect 34808 29174 34940 29180
rect 34808 29158 34928 29174
rect 34808 28626 34836 29158
rect 34992 29102 35020 29446
rect 36372 29238 36400 29446
rect 36360 29232 36412 29238
rect 36360 29174 36412 29180
rect 36648 29170 36676 31622
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 36820 29164 36872 29170
rect 36820 29106 36872 29112
rect 34980 29096 35032 29102
rect 34980 29038 35032 29044
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 34808 28150 34836 28562
rect 34796 28144 34848 28150
rect 34796 28086 34848 28092
rect 34704 27600 34756 27606
rect 34256 26450 34284 27586
rect 34704 27542 34756 27548
rect 34716 27130 34744 27542
rect 34808 27130 34836 28086
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34704 27124 34756 27130
rect 34704 27066 34756 27072
rect 34796 27124 34848 27130
rect 34796 27066 34848 27072
rect 35348 27124 35400 27130
rect 35348 27066 35400 27072
rect 34336 26988 34388 26994
rect 34336 26930 34388 26936
rect 34348 26586 34376 26930
rect 34612 26784 34664 26790
rect 34612 26726 34664 26732
rect 34336 26580 34388 26586
rect 34336 26522 34388 26528
rect 34624 26450 34652 26726
rect 34716 26586 34744 27066
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34808 26586 34836 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 34244 26444 34296 26450
rect 34244 26386 34296 26392
rect 34612 26444 34664 26450
rect 34612 26386 34664 26392
rect 35360 26296 35388 27066
rect 35440 26308 35492 26314
rect 35360 26268 35440 26296
rect 34336 26240 34388 26246
rect 34336 26182 34388 26188
rect 33968 26036 34020 26042
rect 33968 25978 34020 25984
rect 34348 25838 34376 26182
rect 35360 25974 35388 26268
rect 35440 26250 35492 26256
rect 36544 26308 36596 26314
rect 36544 26250 36596 26256
rect 35348 25968 35400 25974
rect 35348 25910 35400 25916
rect 33784 25832 33836 25838
rect 33784 25774 33836 25780
rect 34336 25832 34388 25838
rect 34336 25774 34388 25780
rect 34612 25832 34664 25838
rect 34612 25774 34664 25780
rect 34624 25498 34652 25774
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34612 25492 34664 25498
rect 34612 25434 34664 25440
rect 33876 24948 33928 24954
rect 33876 24890 33928 24896
rect 33888 24206 33916 24890
rect 35348 24608 35400 24614
rect 35348 24550 35400 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34244 24268 34296 24274
rect 34244 24210 34296 24216
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 33888 23322 33916 24142
rect 33980 23662 34008 24142
rect 33968 23656 34020 23662
rect 33968 23598 34020 23604
rect 33876 23316 33928 23322
rect 33876 23258 33928 23264
rect 33980 23118 34008 23598
rect 34256 23526 34284 24210
rect 35072 24132 35124 24138
rect 35072 24074 35124 24080
rect 34520 24064 34572 24070
rect 34520 24006 34572 24012
rect 34704 24064 34756 24070
rect 34704 24006 34756 24012
rect 34532 23866 34560 24006
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34244 23520 34296 23526
rect 34244 23462 34296 23468
rect 34612 23520 34664 23526
rect 34612 23462 34664 23468
rect 34256 23254 34284 23462
rect 34244 23248 34296 23254
rect 34244 23190 34296 23196
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 33600 22976 33652 22982
rect 34624 22930 34652 23462
rect 33600 22918 33652 22924
rect 34440 22902 34652 22930
rect 34152 22636 34204 22642
rect 34152 22578 34204 22584
rect 33508 22500 33560 22506
rect 33508 22442 33560 22448
rect 33520 22098 33548 22442
rect 33508 22092 33560 22098
rect 33508 22034 33560 22040
rect 33876 21956 33928 21962
rect 33876 21898 33928 21904
rect 33324 21480 33376 21486
rect 33324 21422 33376 21428
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 33244 19514 33272 19654
rect 33232 19508 33284 19514
rect 33232 19450 33284 19456
rect 33336 19394 33364 21422
rect 33888 20398 33916 21898
rect 34164 21894 34192 22578
rect 34244 22432 34296 22438
rect 34244 22374 34296 22380
rect 34152 21888 34204 21894
rect 34152 21830 34204 21836
rect 34164 21690 34192 21830
rect 34152 21684 34204 21690
rect 34152 21626 34204 21632
rect 34060 21548 34112 21554
rect 34256 21536 34284 22374
rect 34440 22148 34468 22902
rect 34716 22778 34744 24006
rect 35084 23662 35112 24074
rect 35360 23866 35388 24550
rect 35348 23860 35400 23866
rect 35348 23802 35400 23808
rect 35072 23656 35124 23662
rect 35072 23598 35124 23604
rect 34796 23588 34848 23594
rect 34796 23530 34848 23536
rect 34704 22772 34756 22778
rect 34624 22732 34704 22760
rect 34624 22250 34652 22732
rect 34704 22714 34756 22720
rect 34808 22710 34836 23530
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35624 23316 35676 23322
rect 35624 23258 35676 23264
rect 35636 23118 35664 23258
rect 35624 23112 35676 23118
rect 35624 23054 35676 23060
rect 35808 23044 35860 23050
rect 35808 22986 35860 22992
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 34796 22704 34848 22710
rect 34796 22646 34848 22652
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 34716 22386 34744 22578
rect 34716 22358 34836 22386
rect 34624 22222 34744 22250
rect 34440 22120 34560 22148
rect 34532 22114 34560 22120
rect 34532 22098 34652 22114
rect 34532 22092 34664 22098
rect 34532 22086 34612 22092
rect 34612 22034 34664 22040
rect 34336 22024 34388 22030
rect 34336 21966 34388 21972
rect 34348 21690 34376 21966
rect 34336 21684 34388 21690
rect 34336 21626 34388 21632
rect 34716 21554 34744 22222
rect 34808 21894 34836 22358
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34112 21508 34284 21536
rect 34704 21548 34756 21554
rect 34060 21490 34112 21496
rect 34704 21490 34756 21496
rect 34808 21146 34836 21830
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21140 34848 21146
rect 34796 21082 34848 21088
rect 34704 21004 34756 21010
rect 34704 20946 34756 20952
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 33876 20392 33928 20398
rect 33876 20334 33928 20340
rect 33244 19366 33364 19394
rect 33140 17740 33192 17746
rect 33060 17700 33140 17728
rect 33140 17682 33192 17688
rect 32864 17672 32916 17678
rect 32864 17614 32916 17620
rect 32772 17604 32824 17610
rect 32772 17546 32824 17552
rect 33140 17604 33192 17610
rect 33244 17592 33272 19366
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 33192 17564 33272 17592
rect 33140 17546 33192 17552
rect 32680 17536 32732 17542
rect 32680 17478 32732 17484
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32404 15496 32456 15502
rect 32404 15438 32456 15444
rect 31944 13524 31996 13530
rect 31944 13466 31996 13472
rect 32128 13524 32180 13530
rect 32128 13466 32180 13472
rect 31760 13388 31812 13394
rect 31760 13330 31812 13336
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 31484 12980 31536 12986
rect 31484 12922 31536 12928
rect 31496 12850 31524 12922
rect 31484 12844 31536 12850
rect 31484 12786 31536 12792
rect 31760 12776 31812 12782
rect 31760 12718 31812 12724
rect 31298 12472 31354 12481
rect 31298 12407 31354 12416
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31116 11688 31168 11694
rect 31116 11630 31168 11636
rect 31128 11354 31156 11630
rect 31116 11348 31168 11354
rect 31116 11290 31168 11296
rect 31206 9616 31262 9625
rect 31206 9551 31262 9560
rect 31220 9450 31248 9551
rect 31208 9444 31260 9450
rect 31208 9386 31260 9392
rect 31312 7886 31340 12407
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31404 11150 31432 11698
rect 31392 11144 31444 11150
rect 31392 11086 31444 11092
rect 31392 9444 31444 9450
rect 31392 9386 31444 9392
rect 31404 9042 31432 9386
rect 31392 9036 31444 9042
rect 31392 8978 31444 8984
rect 31392 8900 31444 8906
rect 31392 8842 31444 8848
rect 31404 8498 31432 8842
rect 31772 8634 31800 12718
rect 31956 12714 31984 13466
rect 32508 12782 32536 16594
rect 32692 14346 32720 17478
rect 33336 16590 33364 19110
rect 33416 18148 33468 18154
rect 33416 18090 33468 18096
rect 33428 17678 33456 18090
rect 33784 17876 33836 17882
rect 33784 17818 33836 17824
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33796 17610 33824 17818
rect 33784 17604 33836 17610
rect 33784 17546 33836 17552
rect 33324 16584 33376 16590
rect 33324 16526 33376 16532
rect 33980 16114 34008 20538
rect 34428 20392 34480 20398
rect 34428 20334 34480 20340
rect 34244 19712 34296 19718
rect 34244 19654 34296 19660
rect 34256 19378 34284 19654
rect 34440 19514 34468 20334
rect 34532 19718 34560 20878
rect 34716 19990 34744 20946
rect 35164 20936 35216 20942
rect 35360 20924 35388 22918
rect 35820 22710 35848 22986
rect 35900 22976 35952 22982
rect 35900 22918 35952 22924
rect 35912 22778 35940 22918
rect 35900 22772 35952 22778
rect 35900 22714 35952 22720
rect 35808 22704 35860 22710
rect 35808 22646 35860 22652
rect 35440 22160 35492 22166
rect 35440 22102 35492 22108
rect 35216 20896 35388 20924
rect 35164 20878 35216 20884
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 34808 20058 34836 20402
rect 35452 20398 35480 22102
rect 35820 22098 35848 22646
rect 35900 22432 35952 22438
rect 35900 22374 35952 22380
rect 35808 22092 35860 22098
rect 35808 22034 35860 22040
rect 35912 21962 35940 22374
rect 35900 21956 35952 21962
rect 35900 21898 35952 21904
rect 35912 21010 35940 21898
rect 35900 21004 35952 21010
rect 35900 20946 35952 20952
rect 35912 20602 35940 20946
rect 35900 20596 35952 20602
rect 35900 20538 35952 20544
rect 35440 20392 35492 20398
rect 35440 20334 35492 20340
rect 35348 20324 35400 20330
rect 35348 20266 35400 20272
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34796 20052 34848 20058
rect 34796 19994 34848 20000
rect 35360 19990 35388 20266
rect 34704 19984 34756 19990
rect 34704 19926 34756 19932
rect 35348 19984 35400 19990
rect 35348 19926 35400 19932
rect 35072 19848 35124 19854
rect 35072 19790 35124 19796
rect 34520 19712 34572 19718
rect 34520 19654 34572 19660
rect 34428 19508 34480 19514
rect 34428 19450 34480 19456
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34532 19242 34560 19654
rect 35084 19514 35112 19790
rect 35072 19508 35124 19514
rect 35072 19450 35124 19456
rect 34520 19236 34572 19242
rect 34520 19178 34572 19184
rect 35348 19236 35400 19242
rect 35348 19178 35400 19184
rect 34796 19168 34848 19174
rect 34796 19110 34848 19116
rect 34704 18896 34756 18902
rect 34704 18838 34756 18844
rect 34716 18290 34744 18838
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 34808 18222 34836 19110
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18850 35388 19178
rect 35176 18834 35388 18850
rect 35452 18834 35480 20334
rect 35912 19854 35940 20538
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 36188 20058 36216 20402
rect 36176 20052 36228 20058
rect 36176 19994 36228 20000
rect 35900 19848 35952 19854
rect 35900 19790 35952 19796
rect 35716 19168 35768 19174
rect 35716 19110 35768 19116
rect 35532 18896 35584 18902
rect 35532 18838 35584 18844
rect 35164 18828 35388 18834
rect 35216 18822 35388 18828
rect 35440 18828 35492 18834
rect 35164 18770 35216 18776
rect 35440 18770 35492 18776
rect 35176 18426 35204 18770
rect 35544 18426 35572 18838
rect 35728 18698 35756 19110
rect 35716 18692 35768 18698
rect 35716 18634 35768 18640
rect 36280 18630 36308 20402
rect 36268 18624 36320 18630
rect 36268 18566 36320 18572
rect 35164 18420 35216 18426
rect 35164 18362 35216 18368
rect 35532 18420 35584 18426
rect 35532 18362 35584 18368
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34060 17536 34112 17542
rect 34060 17478 34112 17484
rect 34428 17536 34480 17542
rect 34428 17478 34480 17484
rect 34072 17338 34100 17478
rect 34440 17338 34468 17478
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 34428 17332 34480 17338
rect 34428 17274 34480 17280
rect 34520 17264 34572 17270
rect 34348 17212 34520 17218
rect 35532 17264 35584 17270
rect 34348 17206 34572 17212
rect 35530 17232 35532 17241
rect 35584 17232 35586 17241
rect 34348 17190 34560 17206
rect 34348 17134 34376 17190
rect 35530 17167 35586 17176
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34520 17128 34572 17134
rect 34520 17070 34572 17076
rect 34704 17128 34756 17134
rect 34704 17070 34756 17076
rect 34980 17128 35032 17134
rect 34980 17070 35032 17076
rect 34348 16250 34376 17070
rect 34532 16998 34560 17070
rect 34428 16992 34480 16998
rect 34428 16934 34480 16940
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34612 16992 34664 16998
rect 34612 16934 34664 16940
rect 34440 16810 34468 16934
rect 34624 16810 34652 16934
rect 34440 16782 34652 16810
rect 34716 16794 34744 17070
rect 34992 16998 35020 17070
rect 34980 16992 35032 16998
rect 34980 16934 35032 16940
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16794 35388 16934
rect 34704 16788 34756 16794
rect 34704 16730 34756 16736
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 34796 16652 34848 16658
rect 34796 16594 34848 16600
rect 34336 16244 34388 16250
rect 34336 16186 34388 16192
rect 32864 16108 32916 16114
rect 32864 16050 32916 16056
rect 33968 16108 34020 16114
rect 33968 16050 34020 16056
rect 32876 15094 32904 16050
rect 33876 16040 33928 16046
rect 33876 15982 33928 15988
rect 33888 15706 33916 15982
rect 33876 15700 33928 15706
rect 33876 15642 33928 15648
rect 32956 15360 33008 15366
rect 32956 15302 33008 15308
rect 32864 15088 32916 15094
rect 32864 15030 32916 15036
rect 32968 14958 32996 15302
rect 33048 15088 33100 15094
rect 33048 15030 33100 15036
rect 32956 14952 33008 14958
rect 32956 14894 33008 14900
rect 32968 14482 32996 14894
rect 33060 14618 33088 15030
rect 33416 15020 33468 15026
rect 33416 14962 33468 14968
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 32956 14476 33008 14482
rect 32956 14418 33008 14424
rect 32680 14340 32732 14346
rect 32680 14282 32732 14288
rect 33244 13938 33272 14758
rect 33428 14634 33456 14962
rect 33600 14816 33652 14822
rect 33600 14758 33652 14764
rect 33336 14618 33456 14634
rect 33324 14612 33456 14618
rect 33376 14606 33456 14612
rect 33324 14554 33376 14560
rect 33336 14074 33364 14554
rect 33612 14482 33640 14758
rect 33600 14476 33652 14482
rect 33652 14436 33732 14464
rect 33600 14418 33652 14424
rect 33324 14068 33376 14074
rect 33324 14010 33376 14016
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 32588 13864 32640 13870
rect 32588 13806 32640 13812
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 31944 12708 31996 12714
rect 31944 12650 31996 12656
rect 32036 11552 32088 11558
rect 32036 11494 32088 11500
rect 32048 11150 32076 11494
rect 32600 11354 32628 13806
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 32968 13326 32996 13670
rect 32956 13320 33008 13326
rect 32956 13262 33008 13268
rect 33048 13252 33100 13258
rect 33048 13194 33100 13200
rect 33060 12986 33088 13194
rect 33152 12986 33180 13874
rect 33600 13728 33652 13734
rect 33600 13670 33652 13676
rect 33508 13320 33560 13326
rect 33508 13262 33560 13268
rect 33324 13252 33376 13258
rect 33324 13194 33376 13200
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 33140 12980 33192 12986
rect 33140 12922 33192 12928
rect 33336 12918 33364 13194
rect 33520 12986 33548 13262
rect 33612 13190 33640 13670
rect 33704 13530 33732 14436
rect 34060 14408 34112 14414
rect 34060 14350 34112 14356
rect 33876 14000 33928 14006
rect 33876 13942 33928 13948
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 33692 13524 33744 13530
rect 33692 13466 33744 13472
rect 33796 13326 33824 13874
rect 33888 13326 33916 13942
rect 33968 13932 34020 13938
rect 33968 13874 34020 13880
rect 33784 13320 33836 13326
rect 33784 13262 33836 13268
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 33600 13184 33652 13190
rect 33600 13126 33652 13132
rect 33508 12980 33560 12986
rect 33508 12922 33560 12928
rect 33324 12912 33376 12918
rect 33324 12854 33376 12860
rect 32956 12844 33008 12850
rect 32876 12804 32956 12832
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32324 10674 32352 11086
rect 32588 11008 32640 11014
rect 32588 10950 32640 10956
rect 31944 10668 31996 10674
rect 31944 10610 31996 10616
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 31956 9450 31984 10610
rect 32508 10470 32536 10610
rect 32600 10606 32628 10950
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 32508 10062 32536 10406
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32128 9920 32180 9926
rect 32128 9862 32180 9868
rect 32140 9674 32168 9862
rect 32140 9654 32260 9674
rect 32876 9654 32904 12804
rect 32956 12786 33008 12792
rect 32956 11892 33008 11898
rect 32956 11834 33008 11840
rect 32968 11218 32996 11834
rect 33232 11688 33284 11694
rect 33232 11630 33284 11636
rect 33244 11286 33272 11630
rect 33232 11280 33284 11286
rect 33232 11222 33284 11228
rect 32956 11212 33008 11218
rect 32956 11154 33008 11160
rect 33140 11144 33192 11150
rect 33140 11086 33192 11092
rect 33152 10470 33180 11086
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 33244 9926 33272 11222
rect 33232 9920 33284 9926
rect 33232 9862 33284 9868
rect 32140 9648 32272 9654
rect 32140 9646 32220 9648
rect 32220 9590 32272 9596
rect 32864 9648 32916 9654
rect 32864 9590 32916 9596
rect 33140 9648 33192 9654
rect 33140 9590 33192 9596
rect 31944 9444 31996 9450
rect 31944 9386 31996 9392
rect 31956 8974 31984 9386
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 32048 9110 32076 9318
rect 32036 9104 32088 9110
rect 32036 9046 32088 9052
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 31760 8628 31812 8634
rect 31760 8570 31812 8576
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 31760 8424 31812 8430
rect 31760 8366 31812 8372
rect 31668 8016 31720 8022
rect 31668 7958 31720 7964
rect 31300 7880 31352 7886
rect 31220 7828 31300 7834
rect 31220 7822 31352 7828
rect 31220 7806 31340 7822
rect 31680 7818 31708 7958
rect 31772 7954 31800 8366
rect 31864 8090 31892 8910
rect 31852 8084 31904 8090
rect 31852 8026 31904 8032
rect 31760 7948 31812 7954
rect 31760 7890 31812 7896
rect 31668 7812 31720 7818
rect 31024 7472 31076 7478
rect 31024 7414 31076 7420
rect 31220 6866 31248 7806
rect 31668 7754 31720 7760
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 31484 7744 31536 7750
rect 31484 7686 31536 7692
rect 31312 7546 31340 7686
rect 31496 7546 31524 7686
rect 31300 7540 31352 7546
rect 31300 7482 31352 7488
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31312 7002 31340 7278
rect 31772 7206 31800 7890
rect 31864 7410 31892 8026
rect 31852 7404 31904 7410
rect 31852 7346 31904 7352
rect 31760 7200 31812 7206
rect 31760 7142 31812 7148
rect 31300 6996 31352 7002
rect 31300 6938 31352 6944
rect 31208 6860 31260 6866
rect 31208 6802 31260 6808
rect 31944 6792 31996 6798
rect 31944 6734 31996 6740
rect 31116 6656 31168 6662
rect 31116 6598 31168 6604
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 31128 5914 31156 6598
rect 31220 6458 31248 6598
rect 31956 6458 31984 6734
rect 31208 6452 31260 6458
rect 31208 6394 31260 6400
rect 31944 6452 31996 6458
rect 31944 6394 31996 6400
rect 32048 6390 32076 9046
rect 32232 8906 32260 9590
rect 32588 9580 32640 9586
rect 32588 9522 32640 9528
rect 32600 9178 32628 9522
rect 33152 9178 33180 9590
rect 33232 9444 33284 9450
rect 33232 9386 33284 9392
rect 32588 9172 32640 9178
rect 32588 9114 32640 9120
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 32496 8968 32548 8974
rect 32496 8910 32548 8916
rect 32220 8900 32272 8906
rect 32220 8842 32272 8848
rect 32128 7336 32180 7342
rect 32128 7278 32180 7284
rect 32140 6458 32168 7278
rect 32508 6866 32536 8910
rect 32968 8634 32996 8978
rect 33140 8968 33192 8974
rect 33244 8956 33272 9386
rect 33612 9178 33640 13126
rect 33796 11762 33824 13262
rect 33980 12850 34008 13874
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33784 11756 33836 11762
rect 33784 11698 33836 11704
rect 33876 11620 33928 11626
rect 33876 11562 33928 11568
rect 33888 10742 33916 11562
rect 33876 10736 33928 10742
rect 33796 10684 33876 10690
rect 33796 10678 33928 10684
rect 33692 10668 33744 10674
rect 33692 10610 33744 10616
rect 33796 10662 33916 10678
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33192 8928 33364 8956
rect 33140 8910 33192 8916
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 32956 8628 33008 8634
rect 32956 8570 33008 8576
rect 33152 7002 33180 8774
rect 33336 8430 33364 8928
rect 33324 8424 33376 8430
rect 33324 8366 33376 8372
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 33140 6996 33192 7002
rect 33140 6938 33192 6944
rect 32496 6860 32548 6866
rect 32496 6802 32548 6808
rect 33244 6798 33272 8298
rect 33704 7546 33732 10610
rect 33796 8974 33824 10662
rect 33876 10532 33928 10538
rect 33876 10474 33928 10480
rect 33888 10062 33916 10474
rect 34072 10062 34100 14350
rect 34244 13184 34296 13190
rect 34244 13126 34296 13132
rect 34256 12986 34284 13126
rect 34244 12980 34296 12986
rect 34244 12922 34296 12928
rect 34336 12708 34388 12714
rect 34336 12650 34388 12656
rect 33876 10056 33928 10062
rect 33876 9998 33928 10004
rect 33968 10056 34020 10062
rect 33968 9998 34020 10004
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 33980 9722 34008 9998
rect 33968 9716 34020 9722
rect 33968 9658 34020 9664
rect 33784 8968 33836 8974
rect 33784 8910 33836 8916
rect 33796 8498 33824 8910
rect 33784 8492 33836 8498
rect 33784 8434 33836 8440
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 33324 7268 33376 7274
rect 33324 7210 33376 7216
rect 33232 6792 33284 6798
rect 33232 6734 33284 6740
rect 32588 6724 32640 6730
rect 32588 6666 32640 6672
rect 32128 6452 32180 6458
rect 32128 6394 32180 6400
rect 31760 6384 31812 6390
rect 31760 6326 31812 6332
rect 32036 6384 32088 6390
rect 32036 6326 32088 6332
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 30760 5766 30880 5794
rect 30852 5710 30880 5766
rect 30840 5704 30892 5710
rect 30840 5646 30892 5652
rect 30748 5636 30800 5642
rect 30748 5578 30800 5584
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30196 5160 30248 5166
rect 30196 5102 30248 5108
rect 30208 4826 30236 5102
rect 30392 5098 30420 5510
rect 30656 5228 30708 5234
rect 30656 5170 30708 5176
rect 30380 5092 30432 5098
rect 30380 5034 30432 5040
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 30668 4622 30696 5170
rect 30760 4826 30788 5578
rect 30852 5370 30880 5646
rect 30840 5364 30892 5370
rect 30840 5306 30892 5312
rect 31772 5302 31800 6326
rect 32600 6322 32628 6666
rect 33140 6656 33192 6662
rect 33140 6598 33192 6604
rect 33152 6390 33180 6598
rect 33140 6384 33192 6390
rect 33140 6326 33192 6332
rect 32496 6316 32548 6322
rect 32496 6258 32548 6264
rect 32588 6316 32640 6322
rect 32588 6258 32640 6264
rect 32036 6248 32088 6254
rect 32036 6190 32088 6196
rect 32048 5914 32076 6190
rect 32508 5914 32536 6258
rect 33336 6118 33364 7210
rect 34072 7206 34100 9998
rect 34348 9994 34376 12650
rect 34808 11234 34836 16594
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34808 11206 34928 11234
rect 34900 10810 34928 11206
rect 34888 10804 34940 10810
rect 34888 10746 34940 10752
rect 36556 10674 36584 26250
rect 36832 22094 36860 29106
rect 37280 29028 37332 29034
rect 37280 28970 37332 28976
rect 37292 23118 37320 28970
rect 37280 23112 37332 23118
rect 37280 23054 37332 23060
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37384 22778 37412 22918
rect 37372 22772 37424 22778
rect 37372 22714 37424 22720
rect 37830 22536 37886 22545
rect 37830 22471 37832 22480
rect 37884 22471 37886 22480
rect 37832 22442 37884 22448
rect 36740 22066 36860 22094
rect 36740 21593 36768 22066
rect 36726 21584 36782 21593
rect 36726 21519 36782 21528
rect 36740 12434 36768 21519
rect 38384 20732 38436 20738
rect 38384 20674 38436 20680
rect 38396 20505 38424 20674
rect 38382 20496 38438 20505
rect 38382 20431 38438 20440
rect 38384 18012 38436 18018
rect 38384 17954 38436 17960
rect 38396 17785 38424 17954
rect 38382 17776 38438 17785
rect 38382 17711 38438 17720
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37660 16017 37688 16050
rect 37646 16008 37702 16017
rect 37646 15943 37702 15952
rect 37832 15904 37884 15910
rect 37832 15846 37884 15852
rect 37844 15745 37872 15846
rect 37830 15736 37886 15745
rect 37830 15671 37886 15680
rect 36648 12406 36768 12434
rect 36648 10674 36676 12406
rect 37278 11656 37334 11665
rect 37278 11591 37334 11600
rect 37292 11150 37320 11591
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 37924 11076 37976 11082
rect 37924 11018 37976 11024
rect 37936 10985 37964 11018
rect 37922 10976 37978 10985
rect 37922 10911 37978 10920
rect 36544 10668 36596 10674
rect 36544 10610 36596 10616
rect 36636 10668 36688 10674
rect 36636 10610 36688 10616
rect 34612 10600 34664 10606
rect 34612 10542 34664 10548
rect 34624 10266 34652 10542
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34612 10260 34664 10266
rect 34612 10202 34664 10208
rect 34336 9988 34388 9994
rect 34336 9930 34388 9936
rect 34348 9450 34376 9930
rect 36648 9489 36676 10610
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36634 9480 36690 9489
rect 34336 9444 34388 9450
rect 36634 9415 36690 9424
rect 34336 9386 34388 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 36648 9042 36676 9415
rect 36636 9036 36688 9042
rect 36636 8978 36688 8984
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 33324 6112 33376 6118
rect 33324 6054 33376 6060
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 32036 5908 32088 5914
rect 32036 5850 32088 5856
rect 32496 5908 32548 5914
rect 32496 5850 32548 5856
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 31956 5370 31984 5646
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 31760 5296 31812 5302
rect 31760 5238 31812 5244
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 30748 4820 30800 4826
rect 30748 4762 30800 4768
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 30656 4616 30708 4622
rect 30656 4558 30708 4564
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36924 3194 36952 10406
rect 38108 8968 38160 8974
rect 38106 8936 38108 8945
rect 38160 8936 38162 8945
rect 38106 8871 38162 8880
rect 36912 3188 36964 3194
rect 36912 3130 36964 3136
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 37188 2848 37240 2854
rect 37188 2790 37240 2796
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 13004 2446 13032 2790
rect 16224 2446 16252 2790
rect 17420 2446 17448 2790
rect 21928 2446 21956 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 2136 2440 2188 2446
rect 4068 2440 4120 2446
rect 2136 2382 2188 2388
rect 3896 2366 4016 2394
rect 4068 2382 4120 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 32 800 60 2246
rect 1964 800 1992 2246
rect 3896 800 3924 2366
rect 3988 2310 4016 2366
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6472 870 6592 898
rect 6472 800 6500 870
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 6564 762 6592 870
rect 6840 762 6868 2246
rect 8496 1306 8524 2382
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11164 1442 11192 2314
rect 12900 2304 12952 2310
rect 15016 2304 15068 2310
rect 12900 2246 12952 2252
rect 14844 2264 15016 2292
rect 8404 1278 8524 1306
rect 10980 1414 11192 1442
rect 8404 800 8432 1278
rect 10980 800 11008 1414
rect 12912 800 12940 2246
rect 14844 800 14872 2264
rect 15016 2246 15068 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 17420 800 17448 2246
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 26436 800 26464 2246
rect 37200 1465 37228 2790
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 37476 1306 37504 2382
rect 37384 1278 37504 1306
rect 37384 800 37412 1278
rect 6564 734 6868 762
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 34794 0 34850 800
rect 37370 0 37426 800
rect 39302 0 39358 800
<< via2 >>
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 938 36760 994 36816
rect 1582 24948 1638 24984
rect 1582 24928 1584 24948
rect 1584 24928 1636 24948
rect 1636 24928 1638 24948
rect 3054 22636 3110 22672
rect 3054 22616 3056 22636
rect 3056 22616 3108 22636
rect 3108 22616 3110 22636
rect 2410 21548 2466 21584
rect 2410 21528 2412 21548
rect 2412 21528 2464 21548
rect 2464 21528 2466 21548
rect 2226 20576 2282 20632
rect 938 20440 994 20496
rect 938 18400 994 18456
rect 938 15680 994 15736
rect 938 13640 994 13696
rect 938 11600 994 11656
rect 938 8880 994 8936
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 5170 38392 5226 38448
rect 6458 38256 6514 38312
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27240 4122 27296
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4618 23060 4620 23080
rect 4620 23060 4672 23080
rect 4672 23060 4674 23080
rect 4618 23024 4674 23060
rect 4066 22636 4122 22672
rect 4066 22616 4068 22636
rect 4068 22616 4120 22636
rect 4120 22616 4122 22636
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3974 22072 4030 22128
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4066 20460 4122 20496
rect 4066 20440 4068 20460
rect 4068 20440 4120 20460
rect 4120 20440 4122 20460
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3146 18808 3202 18864
rect 4986 21836 4988 21856
rect 4988 21836 5040 21856
rect 5040 21836 5042 21856
rect 4986 21800 5042 21836
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4434 17176 4490 17232
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3238 9560 3294 9616
rect 1490 6840 1546 6896
rect 938 4120 994 4176
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 8492 4122 8528
rect 4066 8472 4068 8492
rect 4068 8472 4120 8492
rect 4120 8472 4122 8492
rect 8298 26288 8354 26344
rect 6642 22480 6698 22536
rect 7102 22480 7158 22536
rect 5538 17992 5594 18048
rect 5446 16496 5502 16552
rect 6366 17176 6422 17232
rect 6642 20440 6698 20496
rect 7838 23024 7894 23080
rect 7838 22616 7894 22672
rect 7010 21392 7066 21448
rect 5446 9580 5502 9616
rect 5446 9560 5448 9580
rect 5448 9560 5500 9580
rect 5500 9560 5502 9580
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 7470 17740 7526 17776
rect 7470 17720 7472 17740
rect 7472 17720 7524 17740
rect 7524 17720 7526 17740
rect 8022 17484 8024 17504
rect 8024 17484 8076 17504
rect 8076 17484 8078 17504
rect 8022 17448 8078 17484
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 8482 22480 8538 22536
rect 8298 22108 8300 22128
rect 8300 22108 8352 22128
rect 8352 22108 8354 22128
rect 8298 22072 8354 22108
rect 9310 22092 9366 22128
rect 9770 30232 9826 30288
rect 9310 22072 9312 22092
rect 9312 22072 9364 22092
rect 9364 22072 9366 22092
rect 9034 20712 9090 20768
rect 8666 19760 8722 19816
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 10966 30268 10968 30288
rect 10968 30268 11020 30288
rect 11020 30268 11022 30288
rect 10966 30232 11022 30268
rect 11702 37868 11758 37904
rect 11702 37848 11704 37868
rect 11704 37848 11756 37868
rect 11756 37848 11758 37868
rect 12990 38664 13046 38720
rect 22098 38664 22154 38720
rect 11702 32020 11758 32056
rect 11702 32000 11704 32020
rect 11704 32000 11756 32020
rect 11756 32000 11758 32020
rect 12346 33768 12402 33824
rect 11978 32816 12034 32872
rect 12990 35980 12992 36000
rect 12992 35980 13044 36000
rect 13044 35980 13046 36000
rect 12990 35944 13046 35980
rect 12070 29552 12126 29608
rect 9034 15972 9090 16008
rect 9034 15952 9036 15972
rect 9036 15952 9088 15972
rect 9088 15952 9090 15972
rect 9034 15136 9090 15192
rect 9954 18944 10010 19000
rect 9862 18264 9918 18320
rect 9586 17484 9588 17504
rect 9588 17484 9640 17504
rect 9640 17484 9642 17504
rect 9586 17448 9642 17484
rect 9678 16360 9734 16416
rect 10322 20712 10378 20768
rect 8206 9596 8208 9616
rect 8208 9596 8260 9616
rect 8260 9596 8262 9616
rect 8206 9560 8262 9596
rect 10414 19080 10470 19136
rect 10414 17992 10470 18048
rect 8942 9560 8998 9616
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10138 10648 10194 10704
rect 10598 18708 10600 18728
rect 10600 18708 10652 18728
rect 10652 18708 10654 18728
rect 10598 18672 10654 18708
rect 10598 18164 10600 18184
rect 10600 18164 10652 18184
rect 10652 18164 10654 18184
rect 10598 18128 10654 18164
rect 12070 25200 12126 25256
rect 11886 21256 11942 21312
rect 11610 20304 11666 20360
rect 10966 18708 10968 18728
rect 10968 18708 11020 18728
rect 11020 18708 11022 18728
rect 10966 18672 11022 18708
rect 11334 18128 11390 18184
rect 11242 17856 11298 17912
rect 10322 10376 10378 10432
rect 11886 19236 11942 19272
rect 11886 19216 11888 19236
rect 11888 19216 11940 19236
rect 11940 19216 11942 19236
rect 11702 17992 11758 18048
rect 13174 32000 13230 32056
rect 12806 27104 12862 27160
rect 12714 24284 12716 24304
rect 12716 24284 12768 24304
rect 12768 24284 12770 24304
rect 12714 24248 12770 24284
rect 12254 21972 12256 21992
rect 12256 21972 12308 21992
rect 12308 21972 12310 21992
rect 12254 21936 12310 21972
rect 12162 20304 12218 20360
rect 12070 17584 12126 17640
rect 12438 18672 12494 18728
rect 12714 19080 12770 19136
rect 12622 17992 12678 18048
rect 12806 17448 12862 17504
rect 13358 29028 13414 29064
rect 13358 29008 13360 29028
rect 13360 29008 13412 29028
rect 13412 29008 13414 29028
rect 13174 24792 13230 24848
rect 13358 23860 13414 23896
rect 13358 23840 13360 23860
rect 13360 23840 13412 23860
rect 13412 23840 13414 23860
rect 14094 33360 14150 33416
rect 13910 29824 13966 29880
rect 14462 37304 14518 37360
rect 15106 36760 15162 36816
rect 14186 29552 14242 29608
rect 15198 31456 15254 31512
rect 15014 30096 15070 30152
rect 14554 27548 14556 27568
rect 14556 27548 14608 27568
rect 14608 27548 14610 27568
rect 14554 27512 14610 27548
rect 14186 27240 14242 27296
rect 13726 25356 13782 25392
rect 13726 25336 13728 25356
rect 13728 25336 13780 25356
rect 13780 25336 13782 25356
rect 14094 24268 14150 24304
rect 14094 24248 14096 24268
rect 14096 24248 14148 24268
rect 14148 24248 14150 24268
rect 13358 21684 13414 21720
rect 13358 21664 13360 21684
rect 13360 21664 13412 21684
rect 13412 21664 13414 21684
rect 12990 19080 13046 19136
rect 13082 18708 13084 18728
rect 13084 18708 13136 18728
rect 13136 18708 13138 18728
rect 13082 18672 13138 18708
rect 13082 17312 13138 17368
rect 12898 16396 12900 16416
rect 12900 16396 12952 16416
rect 12952 16396 12954 16416
rect 12898 16360 12954 16396
rect 13082 15680 13138 15736
rect 13266 11056 13322 11112
rect 13910 23860 13966 23896
rect 13910 23840 13912 23860
rect 13912 23840 13964 23860
rect 13964 23840 13966 23860
rect 13818 19896 13874 19952
rect 13634 19488 13690 19544
rect 13634 19080 13690 19136
rect 13726 16768 13782 16824
rect 14830 26424 14886 26480
rect 15290 30368 15346 30424
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 15566 30504 15622 30560
rect 15382 29960 15438 30016
rect 15566 29280 15622 29336
rect 15474 28464 15530 28520
rect 15382 27940 15438 27976
rect 15382 27920 15384 27940
rect 15384 27920 15436 27940
rect 15436 27920 15438 27940
rect 15382 27104 15438 27160
rect 17774 36252 17776 36272
rect 17776 36252 17828 36272
rect 17828 36252 17830 36272
rect 17774 36216 17830 36252
rect 16486 33360 16542 33416
rect 16578 32136 16634 32192
rect 16486 31864 16542 31920
rect 15842 29960 15898 30016
rect 15566 24792 15622 24848
rect 16210 29180 16212 29200
rect 16212 29180 16264 29200
rect 16264 29180 16266 29200
rect 16210 29144 16266 29180
rect 16118 28076 16174 28112
rect 16118 28056 16120 28076
rect 16120 28056 16172 28076
rect 16172 28056 16174 28076
rect 16854 34040 16910 34096
rect 17406 33396 17408 33416
rect 17408 33396 17460 33416
rect 17460 33396 17462 33416
rect 17406 33360 17462 33396
rect 17866 34040 17922 34096
rect 18326 35672 18382 35728
rect 17590 31864 17646 31920
rect 18142 32816 18198 32872
rect 18234 32000 18290 32056
rect 17774 31320 17830 31376
rect 15934 24792 15990 24848
rect 15566 23704 15622 23760
rect 14002 19080 14058 19136
rect 14278 20032 14334 20088
rect 14922 19216 14978 19272
rect 14922 17992 14978 18048
rect 15842 24112 15898 24168
rect 15842 24012 15844 24032
rect 15844 24012 15896 24032
rect 15896 24012 15898 24032
rect 15842 23976 15898 24012
rect 15842 23568 15898 23624
rect 16578 25200 16634 25256
rect 16486 23432 16542 23488
rect 15566 17856 15622 17912
rect 15842 15816 15898 15872
rect 15842 15544 15898 15600
rect 15842 15136 15898 15192
rect 15750 15020 15806 15056
rect 15750 15000 15752 15020
rect 15752 15000 15804 15020
rect 15804 15000 15806 15020
rect 16578 19508 16634 19544
rect 16578 19488 16580 19508
rect 16580 19488 16632 19508
rect 16632 19488 16634 19508
rect 17682 30912 17738 30968
rect 17866 30504 17922 30560
rect 17406 27512 17462 27568
rect 18602 36252 18604 36272
rect 18604 36252 18656 36272
rect 18656 36252 18658 36272
rect 18602 36216 18658 36252
rect 18786 33768 18842 33824
rect 18326 30776 18382 30832
rect 18050 29028 18106 29064
rect 18050 29008 18052 29028
rect 18052 29008 18104 29028
rect 18104 29008 18106 29028
rect 17130 24384 17186 24440
rect 18418 28736 18474 28792
rect 17866 24656 17922 24712
rect 16854 19624 16910 19680
rect 16302 15272 16358 15328
rect 16854 15816 16910 15872
rect 15014 9696 15070 9752
rect 16762 14048 16818 14104
rect 17866 20032 17922 20088
rect 17866 19624 17922 19680
rect 17774 17312 17830 17368
rect 17958 16516 18014 16552
rect 17958 16496 17960 16516
rect 17960 16496 18012 16516
rect 18012 16496 18014 16516
rect 18694 30776 18750 30832
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19430 35028 19432 35048
rect 19432 35028 19484 35048
rect 19484 35028 19486 35048
rect 19430 34992 19486 35028
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19430 34740 19486 34776
rect 19430 34720 19432 34740
rect 19432 34720 19484 34740
rect 19484 34720 19486 34740
rect 18694 30232 18750 30288
rect 18970 30912 19026 30968
rect 18970 30388 19026 30424
rect 18970 30368 18972 30388
rect 18972 30368 19024 30388
rect 19024 30368 19026 30388
rect 18878 29960 18934 30016
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19614 33224 19670 33280
rect 19154 30776 19210 30832
rect 19154 29960 19210 30016
rect 18878 29280 18934 29336
rect 19062 29144 19118 29200
rect 18786 29008 18842 29064
rect 18602 26152 18658 26208
rect 22558 38292 22560 38312
rect 22560 38292 22612 38312
rect 22612 38292 22614 38312
rect 22558 38256 22614 38292
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19982 31764 19984 31784
rect 19984 31764 20036 31784
rect 20036 31764 20038 31784
rect 19982 31728 20038 31764
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19890 29960 19946 30016
rect 20166 31320 20222 31376
rect 20442 34620 20444 34640
rect 20444 34620 20496 34640
rect 20496 34620 20498 34640
rect 20442 34584 20498 34620
rect 20442 34176 20498 34232
rect 20810 34176 20866 34232
rect 21270 35012 21326 35048
rect 21270 34992 21272 35012
rect 21272 34992 21324 35012
rect 21324 34992 21326 35012
rect 20902 32136 20958 32192
rect 20442 31592 20498 31648
rect 19798 29552 19854 29608
rect 19982 29416 20038 29472
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 20166 29708 20222 29744
rect 20166 29688 20168 29708
rect 20168 29688 20220 29708
rect 20220 29688 20222 29708
rect 20534 31048 20590 31104
rect 20718 30912 20774 30968
rect 21546 34584 21602 34640
rect 21362 31456 21418 31512
rect 22098 36080 22154 36136
rect 22190 35536 22246 35592
rect 22190 35400 22246 35456
rect 22834 35944 22890 36000
rect 22466 34468 22522 34504
rect 21822 33224 21878 33280
rect 21638 31628 21640 31648
rect 21640 31628 21692 31648
rect 21692 31628 21694 31648
rect 21638 31592 21694 31628
rect 20718 30096 20774 30152
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19522 27820 19524 27840
rect 19524 27820 19576 27840
rect 19576 27820 19578 27840
rect 19522 27784 19578 27820
rect 19430 27512 19486 27568
rect 19338 26424 19394 26480
rect 18602 23976 18658 24032
rect 18510 23724 18566 23760
rect 18510 23704 18512 23724
rect 18512 23704 18564 23724
rect 18564 23704 18566 23724
rect 18418 17484 18420 17504
rect 18420 17484 18472 17504
rect 18472 17484 18474 17504
rect 18418 17448 18474 17484
rect 17866 15544 17922 15600
rect 17958 15000 18014 15056
rect 17866 13912 17922 13968
rect 11794 3984 11850 4040
rect 13174 3984 13230 4040
rect 18326 15136 18382 15192
rect 18142 9696 18198 9752
rect 17866 9560 17922 9616
rect 18970 18128 19026 18184
rect 18786 14068 18842 14104
rect 18786 14048 18788 14068
rect 18788 14048 18840 14068
rect 18840 14048 18842 14068
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19706 25764 19762 25800
rect 19706 25744 19708 25764
rect 19708 25744 19760 25764
rect 19760 25744 19762 25764
rect 19706 25472 19762 25528
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 21270 29824 21326 29880
rect 20534 27376 20590 27432
rect 20534 26424 20590 26480
rect 20258 25064 20314 25120
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19246 18128 19302 18184
rect 20994 27648 21050 27704
rect 20810 27512 20866 27568
rect 20902 26424 20958 26480
rect 20810 26188 20812 26208
rect 20812 26188 20864 26208
rect 20864 26188 20866 26208
rect 20810 26152 20866 26188
rect 20534 24928 20590 24984
rect 20442 24792 20498 24848
rect 20626 24520 20682 24576
rect 20626 24112 20682 24168
rect 20718 23704 20774 23760
rect 21178 25472 21234 25528
rect 20442 23160 20498 23216
rect 20994 23568 21050 23624
rect 20902 23160 20958 23216
rect 21086 23432 21142 23488
rect 21454 29960 21510 30016
rect 22466 34448 22468 34468
rect 22468 34448 22520 34468
rect 22520 34448 22522 34468
rect 22098 32544 22154 32600
rect 21914 31592 21970 31648
rect 22374 32680 22430 32736
rect 22190 31764 22192 31784
rect 22192 31764 22244 31784
rect 22244 31764 22246 31784
rect 22190 31728 22246 31764
rect 21822 29824 21878 29880
rect 23018 35672 23074 35728
rect 22926 34720 22982 34776
rect 23110 35400 23166 35456
rect 23110 33088 23166 33144
rect 22650 32408 22706 32464
rect 22098 29552 22154 29608
rect 20534 22208 20590 22264
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20166 19488 20222 19544
rect 19890 18672 19946 18728
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19798 18128 19854 18184
rect 19338 17856 19394 17912
rect 19706 17856 19762 17912
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19798 17040 19854 17096
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 21178 22500 21234 22536
rect 21178 22480 21180 22500
rect 21180 22480 21232 22500
rect 21232 22480 21234 22500
rect 21362 23296 21418 23352
rect 20442 17312 20498 17368
rect 23018 32136 23074 32192
rect 22742 32000 22798 32056
rect 23478 34604 23534 34640
rect 23478 34584 23480 34604
rect 23480 34584 23532 34604
rect 23532 34584 23534 34604
rect 23386 31864 23442 31920
rect 22282 28328 22338 28384
rect 22098 27376 22154 27432
rect 22926 30368 22982 30424
rect 22834 29960 22890 30016
rect 22742 28464 22798 28520
rect 22650 28056 22706 28112
rect 22558 27920 22614 27976
rect 22374 25064 22430 25120
rect 22282 24928 22338 24984
rect 22190 24656 22246 24712
rect 22190 24248 22246 24304
rect 21822 22752 21878 22808
rect 22926 28736 22982 28792
rect 23202 30232 23258 30288
rect 23110 29416 23166 29472
rect 22926 28328 22982 28384
rect 25042 38392 25098 38448
rect 27066 38664 27122 38720
rect 31206 38700 31208 38720
rect 31208 38700 31260 38720
rect 31260 38700 31262 38720
rect 31206 38664 31262 38700
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 37922 38800 37978 38856
rect 24582 36760 24638 36816
rect 23846 32272 23902 32328
rect 23754 32136 23810 32192
rect 23938 32000 23994 32056
rect 22834 24656 22890 24712
rect 22466 24112 22522 24168
rect 22006 22480 22062 22536
rect 22650 23568 22706 23624
rect 23202 25880 23258 25936
rect 23110 24792 23166 24848
rect 23570 27512 23626 27568
rect 23754 28600 23810 28656
rect 22466 22344 22522 22400
rect 22190 19896 22246 19952
rect 20442 16532 20444 16552
rect 20444 16532 20496 16552
rect 20496 16532 20498 16552
rect 20442 16496 20498 16532
rect 20350 15408 20406 15464
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19246 11620 19302 11656
rect 19246 11600 19248 11620
rect 19248 11600 19300 11620
rect 19300 11600 19302 11620
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19614 11756 19670 11792
rect 19614 11736 19616 11756
rect 19616 11736 19668 11756
rect 19668 11736 19670 11756
rect 18602 10920 18658 10976
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19890 10004 19892 10024
rect 19892 10004 19944 10024
rect 19944 10004 19946 10024
rect 19890 9968 19946 10004
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 21178 12144 21234 12200
rect 19798 9444 19854 9480
rect 19798 9424 19800 9444
rect 19800 9424 19852 9444
rect 19852 9424 19854 9444
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19982 8628 20038 8664
rect 19982 8608 19984 8628
rect 19984 8608 20036 8628
rect 20036 8608 20038 8628
rect 18694 6840 18750 6896
rect 21086 10140 21088 10160
rect 21088 10140 21140 10160
rect 21140 10140 21142 10160
rect 21086 10104 21142 10140
rect 21086 9968 21142 10024
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 21822 19080 21878 19136
rect 21914 18964 21970 19000
rect 21914 18944 21916 18964
rect 21916 18944 21968 18964
rect 21968 18944 21970 18964
rect 22190 18708 22192 18728
rect 22192 18708 22244 18728
rect 22244 18708 22246 18728
rect 22190 18672 22246 18708
rect 22558 22208 22614 22264
rect 22650 19252 22652 19272
rect 22652 19252 22704 19272
rect 22704 19252 22706 19272
rect 22650 19216 22706 19252
rect 21822 17856 21878 17912
rect 21914 16496 21970 16552
rect 22098 12824 22154 12880
rect 25410 37868 25466 37904
rect 25410 37848 25412 37868
rect 25412 37848 25464 37868
rect 25464 37848 25466 37868
rect 25318 36236 25374 36272
rect 25318 36216 25320 36236
rect 25320 36216 25372 36236
rect 25372 36216 25374 36236
rect 25226 35944 25282 36000
rect 24490 34484 24492 34504
rect 24492 34484 24544 34504
rect 24544 34484 24546 34504
rect 24490 34448 24546 34484
rect 24674 34448 24730 34504
rect 24490 32272 24546 32328
rect 24674 28600 24730 28656
rect 24122 25780 24124 25800
rect 24124 25780 24176 25800
rect 24176 25780 24178 25800
rect 24122 25744 24178 25780
rect 24398 24404 24454 24440
rect 24398 24384 24400 24404
rect 24400 24384 24452 24404
rect 24452 24384 24454 24404
rect 24766 26152 24822 26208
rect 24582 25356 24638 25392
rect 24582 25336 24584 25356
rect 24584 25336 24636 25356
rect 24636 25336 24638 25356
rect 24582 24928 24638 24984
rect 24766 25200 24822 25256
rect 25502 35944 25558 36000
rect 25502 35556 25558 35592
rect 25502 35536 25504 35556
rect 25504 35536 25556 35556
rect 25556 35536 25558 35556
rect 25410 34720 25466 34776
rect 25502 34176 25558 34232
rect 26054 36252 26056 36272
rect 26056 36252 26108 36272
rect 26108 36252 26110 36272
rect 26054 36216 26110 36252
rect 26054 36100 26110 36136
rect 26054 36080 26056 36100
rect 26056 36080 26108 36100
rect 26108 36080 26110 36100
rect 25962 34992 26018 35048
rect 25318 31592 25374 31648
rect 25410 29824 25466 29880
rect 24858 24520 24914 24576
rect 23110 21936 23166 21992
rect 23018 21664 23074 21720
rect 23386 20324 23442 20360
rect 23386 20304 23388 20324
rect 23388 20304 23440 20324
rect 23440 20304 23442 20324
rect 23018 19216 23074 19272
rect 23202 18944 23258 19000
rect 22834 17992 22890 18048
rect 23018 18264 23074 18320
rect 22926 17720 22982 17776
rect 23110 17856 23166 17912
rect 22926 16496 22982 16552
rect 23938 21528 23994 21584
rect 23938 19352 23994 19408
rect 24214 19488 24270 19544
rect 24122 18808 24178 18864
rect 23846 17312 23902 17368
rect 24306 16496 24362 16552
rect 24306 15680 24362 15736
rect 23202 15444 23204 15464
rect 23204 15444 23256 15464
rect 23256 15444 23258 15464
rect 23202 15408 23258 15444
rect 21454 10376 21510 10432
rect 21914 10104 21970 10160
rect 23110 13252 23166 13288
rect 23110 13232 23112 13252
rect 23112 13232 23164 13252
rect 23164 13232 23166 13252
rect 22926 12044 22928 12064
rect 22928 12044 22980 12064
rect 22980 12044 22982 12064
rect 22926 12008 22982 12044
rect 22190 10376 22246 10432
rect 22466 10004 22468 10024
rect 22468 10004 22520 10024
rect 22520 10004 22522 10024
rect 22466 9968 22522 10004
rect 22466 9288 22522 9344
rect 23662 13368 23718 13424
rect 23662 9968 23718 10024
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 23846 9560 23902 9616
rect 24950 24112 25006 24168
rect 24858 22072 24914 22128
rect 25870 31456 25926 31512
rect 25870 30368 25926 30424
rect 25778 29552 25834 29608
rect 25502 28328 25558 28384
rect 25318 26152 25374 26208
rect 25410 26016 25466 26072
rect 25410 25064 25466 25120
rect 25686 25064 25742 25120
rect 25778 23568 25834 23624
rect 25410 21392 25466 21448
rect 25410 20848 25466 20904
rect 25410 20460 25466 20496
rect 25594 20576 25650 20632
rect 25410 20440 25412 20460
rect 25412 20440 25464 20460
rect 25464 20440 25466 20460
rect 26238 35400 26294 35456
rect 26054 29688 26110 29744
rect 26054 26288 26110 26344
rect 26054 24520 26110 24576
rect 25962 21548 26018 21584
rect 25962 21528 25964 21548
rect 25964 21528 26016 21548
rect 26016 21528 26018 21548
rect 25778 21256 25834 21312
rect 25778 19780 25834 19816
rect 25778 19760 25780 19780
rect 25780 19760 25832 19780
rect 25832 19760 25834 19780
rect 25686 19216 25742 19272
rect 25318 18128 25374 18184
rect 25778 18808 25834 18864
rect 26514 29824 26570 29880
rect 27158 31864 27214 31920
rect 26606 24248 26662 24304
rect 26974 28328 27030 28384
rect 26882 25880 26938 25936
rect 27066 24792 27122 24848
rect 26974 23432 27030 23488
rect 27066 22752 27122 22808
rect 27250 23296 27306 23352
rect 27250 22636 27306 22672
rect 27250 22616 27252 22636
rect 27252 22616 27304 22636
rect 27304 22616 27306 22636
rect 25134 16108 25190 16144
rect 25134 16088 25136 16108
rect 25136 16088 25188 16108
rect 25188 16088 25190 16108
rect 24858 13776 24914 13832
rect 24490 11772 24492 11792
rect 24492 11772 24544 11792
rect 24544 11772 24546 11792
rect 24490 11736 24546 11772
rect 24398 9968 24454 10024
rect 24490 9424 24546 9480
rect 24306 8472 24362 8528
rect 25042 12824 25098 12880
rect 25042 9288 25098 9344
rect 25318 4120 25374 4176
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 28078 31184 28134 31240
rect 28446 34176 28502 34232
rect 28354 31592 28410 31648
rect 27802 26016 27858 26072
rect 26422 17176 26478 17232
rect 25870 13368 25926 13424
rect 25594 11092 25596 11112
rect 25596 11092 25648 11112
rect 25648 11092 25650 11112
rect 25594 11056 25650 11092
rect 26422 12416 26478 12472
rect 25962 12008 26018 12064
rect 26514 11736 26570 11792
rect 25594 9424 25650 9480
rect 25870 9580 25926 9616
rect 25870 9560 25872 9580
rect 25872 9560 25924 9580
rect 25924 9560 25926 9580
rect 25962 9424 26018 9480
rect 28630 31048 28686 31104
rect 28814 31184 28870 31240
rect 29090 28600 29146 28656
rect 28998 28464 29054 28520
rect 28998 28100 29054 28112
rect 28998 28056 29000 28100
rect 29000 28056 29052 28100
rect 29052 28056 29054 28100
rect 28630 25064 28686 25120
rect 30010 28092 30012 28112
rect 30012 28092 30064 28112
rect 30064 28092 30066 28112
rect 30010 28056 30066 28092
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37278 37188 37334 37224
rect 37278 37168 37280 37188
rect 37280 37168 37332 37188
rect 37332 37168 37334 37188
rect 37830 36760 37886 36816
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 27618 17584 27674 17640
rect 30746 26324 30748 26344
rect 30748 26324 30800 26344
rect 30800 26324 30802 26344
rect 30746 26288 30802 26324
rect 28538 18944 28594 19000
rect 28906 19292 28962 19348
rect 28906 19080 28962 19136
rect 29274 18808 29330 18864
rect 28630 17992 28686 18048
rect 27342 14456 27398 14512
rect 26882 12144 26938 12200
rect 27250 11872 27306 11928
rect 29182 17212 29184 17232
rect 29184 17212 29236 17232
rect 29236 17212 29238 17232
rect 28078 11056 28134 11112
rect 28538 13796 28594 13832
rect 28538 13776 28540 13796
rect 28540 13776 28592 13796
rect 28592 13776 28594 13796
rect 28446 13268 28448 13288
rect 28448 13268 28500 13288
rect 28500 13268 28502 13288
rect 28446 13232 28502 13268
rect 29182 17176 29238 17212
rect 28998 13132 29000 13152
rect 29000 13132 29052 13152
rect 29052 13132 29054 13152
rect 28998 13096 29054 13132
rect 28998 12960 29054 13016
rect 28078 4120 28134 4176
rect 29274 13096 29330 13152
rect 29366 12960 29422 13016
rect 31574 29008 31630 29064
rect 31390 28484 31446 28520
rect 31390 28464 31392 28484
rect 31392 28464 31444 28484
rect 31444 28464 31446 28484
rect 30746 14456 30802 14512
rect 31666 22072 31722 22128
rect 33046 29008 33102 29064
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 32678 22108 32680 22128
rect 32680 22108 32732 22128
rect 32732 22108 32734 22128
rect 31022 17992 31078 18048
rect 29550 9444 29606 9480
rect 29550 9424 29552 9444
rect 29552 9424 29604 9444
rect 29604 9424 29606 9444
rect 32678 22072 32734 22108
rect 37922 34040 37978 34096
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 33690 26308 33746 26344
rect 33690 26288 33692 26308
rect 33692 26288 33744 26308
rect 33744 26288 33746 26308
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 31298 12416 31354 12472
rect 31206 9560 31262 9616
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35530 17212 35532 17232
rect 35532 17212 35584 17232
rect 35584 17212 35586 17232
rect 35530 17176 35586 17212
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 37830 22500 37886 22536
rect 37830 22480 37832 22500
rect 37832 22480 37884 22500
rect 37884 22480 37886 22500
rect 36726 21528 36782 21584
rect 38382 20440 38438 20496
rect 38382 17720 38438 17776
rect 37646 15952 37702 16008
rect 37830 15680 37886 15736
rect 37278 11600 37334 11656
rect 37922 10920 37978 10976
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 36634 9424 36690 9480
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38106 8916 38108 8936
rect 38108 8916 38160 8936
rect 38160 8916 38162 8936
rect 38106 8880 38162 8916
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 37186 1400 37242 1456
<< metal3 >>
rect 0 39448 800 39568
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 37917 38858 37983 38861
rect 38618 38858 39418 38888
rect 37917 38856 39418 38858
rect 37917 38800 37922 38856
rect 37978 38800 39418 38856
rect 37917 38798 39418 38800
rect 37917 38795 37983 38798
rect 38618 38768 39418 38798
rect 12198 38660 12204 38724
rect 12268 38722 12274 38724
rect 12985 38722 13051 38725
rect 12268 38720 13051 38722
rect 12268 38664 12990 38720
rect 13046 38664 13051 38720
rect 12268 38662 13051 38664
rect 12268 38660 12274 38662
rect 12985 38659 13051 38662
rect 22093 38722 22159 38725
rect 23422 38722 23428 38724
rect 22093 38720 23428 38722
rect 22093 38664 22098 38720
rect 22154 38664 23428 38720
rect 22093 38662 23428 38664
rect 22093 38659 22159 38662
rect 23422 38660 23428 38662
rect 23492 38660 23498 38724
rect 23974 38660 23980 38724
rect 24044 38722 24050 38724
rect 27061 38722 27127 38725
rect 24044 38720 27127 38722
rect 24044 38664 27066 38720
rect 27122 38664 27127 38720
rect 24044 38662 27127 38664
rect 24044 38660 24050 38662
rect 27061 38659 27127 38662
rect 27470 38660 27476 38724
rect 27540 38722 27546 38724
rect 31201 38722 31267 38725
rect 27540 38720 31267 38722
rect 27540 38664 31206 38720
rect 31262 38664 31267 38720
rect 27540 38662 31267 38664
rect 27540 38660 27546 38662
rect 31201 38659 31267 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 5165 38450 5231 38453
rect 25037 38450 25103 38453
rect 5165 38448 25103 38450
rect 5165 38392 5170 38448
rect 5226 38392 25042 38448
rect 25098 38392 25103 38448
rect 5165 38390 25103 38392
rect 5165 38387 5231 38390
rect 25037 38387 25103 38390
rect 6453 38314 6519 38317
rect 22553 38314 22619 38317
rect 6453 38312 22619 38314
rect 6453 38256 6458 38312
rect 6514 38256 22558 38312
rect 22614 38256 22619 38312
rect 6453 38254 22619 38256
rect 6453 38251 6519 38254
rect 22553 38251 22619 38254
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 11697 37906 11763 37909
rect 25405 37906 25471 37909
rect 11697 37904 25471 37906
rect 11697 37848 11702 37904
rect 11758 37848 25410 37904
rect 25466 37848 25471 37904
rect 11697 37846 25471 37848
rect 11697 37843 11763 37846
rect 25405 37843 25471 37846
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 14222 37300 14228 37364
rect 14292 37362 14298 37364
rect 14457 37362 14523 37365
rect 14292 37360 14523 37362
rect 14292 37304 14462 37360
rect 14518 37304 14523 37360
rect 14292 37302 14523 37304
rect 14292 37300 14298 37302
rect 14457 37299 14523 37302
rect 13486 37164 13492 37228
rect 13556 37226 13562 37228
rect 37273 37226 37339 37229
rect 13556 37224 37339 37226
rect 13556 37168 37278 37224
rect 37334 37168 37339 37224
rect 13556 37166 37339 37168
rect 13556 37164 13562 37166
rect 37273 37163 37339 37166
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 15101 36818 15167 36821
rect 22318 36818 22324 36820
rect 15101 36816 22324 36818
rect 15101 36760 15106 36816
rect 15162 36760 22324 36816
rect 15101 36758 22324 36760
rect 15101 36755 15167 36758
rect 22318 36756 22324 36758
rect 22388 36818 22394 36820
rect 24577 36818 24643 36821
rect 22388 36816 24643 36818
rect 22388 36760 24582 36816
rect 24638 36760 24643 36816
rect 22388 36758 24643 36760
rect 22388 36756 22394 36758
rect 24577 36755 24643 36758
rect 37825 36818 37891 36821
rect 38618 36818 39418 36848
rect 37825 36816 39418 36818
rect 37825 36760 37830 36816
rect 37886 36760 39418 36816
rect 37825 36758 39418 36760
rect 37825 36755 37891 36758
rect 38618 36728 39418 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 17769 36274 17835 36277
rect 18597 36274 18663 36277
rect 17769 36272 18663 36274
rect 17769 36216 17774 36272
rect 17830 36216 18602 36272
rect 18658 36216 18663 36272
rect 17769 36214 18663 36216
rect 17769 36211 17835 36214
rect 18597 36211 18663 36214
rect 25313 36274 25379 36277
rect 26049 36274 26115 36277
rect 25313 36272 26115 36274
rect 25313 36216 25318 36272
rect 25374 36216 26054 36272
rect 26110 36216 26115 36272
rect 25313 36214 26115 36216
rect 25313 36211 25379 36214
rect 26049 36211 26115 36214
rect 22093 36138 22159 36141
rect 26049 36138 26115 36141
rect 22093 36136 26115 36138
rect 22093 36080 22098 36136
rect 22154 36080 26054 36136
rect 26110 36080 26115 36136
rect 22093 36078 26115 36080
rect 22093 36075 22159 36078
rect 26049 36075 26115 36078
rect 12985 36002 13051 36005
rect 13118 36002 13124 36004
rect 12985 36000 13124 36002
rect 12985 35944 12990 36000
rect 13046 35944 13124 36000
rect 12985 35942 13124 35944
rect 12985 35939 13051 35942
rect 13118 35940 13124 35942
rect 13188 35940 13194 36004
rect 22829 36002 22895 36005
rect 23054 36002 23060 36004
rect 22829 36000 23060 36002
rect 22829 35944 22834 36000
rect 22890 35944 23060 36000
rect 22829 35942 23060 35944
rect 22829 35939 22895 35942
rect 23054 35940 23060 35942
rect 23124 35940 23130 36004
rect 25221 36002 25287 36005
rect 25497 36002 25563 36005
rect 25221 36000 25563 36002
rect 25221 35944 25226 36000
rect 25282 35944 25502 36000
rect 25558 35944 25563 36000
rect 25221 35942 25563 35944
rect 25221 35939 25287 35942
rect 25497 35939 25563 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 18321 35730 18387 35733
rect 23013 35730 23079 35733
rect 18321 35728 23079 35730
rect 18321 35672 18326 35728
rect 18382 35672 23018 35728
rect 23074 35672 23079 35728
rect 18321 35670 23079 35672
rect 18321 35667 18387 35670
rect 23013 35667 23079 35670
rect 22185 35594 22251 35597
rect 25497 35594 25563 35597
rect 22185 35592 25563 35594
rect 22185 35536 22190 35592
rect 22246 35536 25502 35592
rect 25558 35536 25563 35592
rect 22185 35534 25563 35536
rect 22185 35531 22251 35534
rect 25497 35531 25563 35534
rect 22185 35458 22251 35461
rect 22318 35458 22324 35460
rect 22185 35456 22324 35458
rect 22185 35400 22190 35456
rect 22246 35400 22324 35456
rect 22185 35398 22324 35400
rect 22185 35395 22251 35398
rect 22318 35396 22324 35398
rect 22388 35396 22394 35460
rect 23105 35458 23171 35461
rect 26233 35458 26299 35461
rect 23105 35456 26299 35458
rect 23105 35400 23110 35456
rect 23166 35400 26238 35456
rect 26294 35400 26299 35456
rect 23105 35398 26299 35400
rect 23105 35395 23171 35398
rect 26233 35395 26299 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19425 35050 19491 35053
rect 19382 35048 19491 35050
rect 19382 34992 19430 35048
rect 19486 34992 19491 35048
rect 19382 34987 19491 34992
rect 21265 35050 21331 35053
rect 25957 35050 26023 35053
rect 21265 35048 26023 35050
rect 21265 34992 21270 35048
rect 21326 34992 25962 35048
rect 26018 34992 26023 35048
rect 21265 34990 26023 34992
rect 21265 34987 21331 34990
rect 25957 34987 26023 34990
rect 0 34688 800 34808
rect 19382 34781 19442 34987
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 19382 34776 19491 34781
rect 19382 34720 19430 34776
rect 19486 34720 19491 34776
rect 19382 34718 19491 34720
rect 19425 34715 19491 34718
rect 22921 34778 22987 34781
rect 24342 34778 24348 34780
rect 22921 34776 24348 34778
rect 22921 34720 22926 34776
rect 22982 34720 24348 34776
rect 22921 34718 24348 34720
rect 22921 34715 22987 34718
rect 24342 34716 24348 34718
rect 24412 34716 24418 34780
rect 25405 34778 25471 34781
rect 25630 34778 25636 34780
rect 25405 34776 25636 34778
rect 25405 34720 25410 34776
rect 25466 34720 25636 34776
rect 25405 34718 25636 34720
rect 25405 34715 25471 34718
rect 25630 34716 25636 34718
rect 25700 34716 25706 34780
rect 20437 34642 20503 34645
rect 21541 34642 21607 34645
rect 23473 34642 23539 34645
rect 20437 34640 23539 34642
rect 20437 34584 20442 34640
rect 20498 34584 21546 34640
rect 21602 34584 23478 34640
rect 23534 34584 23539 34640
rect 20437 34582 23539 34584
rect 20437 34579 20503 34582
rect 21541 34579 21607 34582
rect 23473 34579 23539 34582
rect 22461 34506 22527 34509
rect 24485 34506 24551 34509
rect 22461 34504 24551 34506
rect 22461 34448 22466 34504
rect 22522 34448 24490 34504
rect 24546 34448 24551 34504
rect 22461 34446 24551 34448
rect 22461 34443 22527 34446
rect 24485 34443 24551 34446
rect 24669 34506 24735 34509
rect 25446 34506 25452 34508
rect 24669 34504 25452 34506
rect 24669 34448 24674 34504
rect 24730 34448 25452 34504
rect 24669 34446 25452 34448
rect 24669 34443 24735 34446
rect 25446 34444 25452 34446
rect 25516 34444 25522 34508
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 20437 34234 20503 34237
rect 20805 34234 20871 34237
rect 25497 34234 25563 34237
rect 28441 34234 28507 34237
rect 20437 34232 28507 34234
rect 20437 34176 20442 34232
rect 20498 34176 20810 34232
rect 20866 34176 25502 34232
rect 25558 34176 28446 34232
rect 28502 34176 28507 34232
rect 20437 34174 28507 34176
rect 20437 34171 20503 34174
rect 20805 34171 20871 34174
rect 25497 34171 25563 34174
rect 28441 34171 28507 34174
rect 16849 34098 16915 34101
rect 17861 34098 17927 34101
rect 16849 34096 17927 34098
rect 16849 34040 16854 34096
rect 16910 34040 17866 34096
rect 17922 34040 17927 34096
rect 16849 34038 17927 34040
rect 16849 34035 16915 34038
rect 17861 34035 17927 34038
rect 37917 34098 37983 34101
rect 38618 34098 39418 34128
rect 37917 34096 39418 34098
rect 37917 34040 37922 34096
rect 37978 34040 39418 34096
rect 37917 34038 39418 34040
rect 37917 34035 37983 34038
rect 38618 34008 39418 34038
rect 12341 33826 12407 33829
rect 18781 33826 18847 33829
rect 12341 33824 18847 33826
rect 12341 33768 12346 33824
rect 12402 33768 18786 33824
rect 18842 33768 18847 33824
rect 12341 33766 18847 33768
rect 12341 33763 12407 33766
rect 18781 33763 18847 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 14089 33418 14155 33421
rect 16481 33418 16547 33421
rect 17401 33418 17467 33421
rect 14089 33416 17467 33418
rect 14089 33360 14094 33416
rect 14150 33360 16486 33416
rect 16542 33360 17406 33416
rect 17462 33360 17467 33416
rect 14089 33358 17467 33360
rect 14089 33355 14155 33358
rect 16481 33355 16547 33358
rect 17401 33355 17467 33358
rect 19609 33282 19675 33285
rect 20662 33282 20668 33284
rect 19609 33280 20668 33282
rect 19609 33224 19614 33280
rect 19670 33224 20668 33280
rect 19609 33222 20668 33224
rect 19609 33219 19675 33222
rect 20662 33220 20668 33222
rect 20732 33220 20738 33284
rect 21817 33282 21883 33285
rect 21950 33282 21956 33284
rect 21817 33280 21956 33282
rect 21817 33224 21822 33280
rect 21878 33224 21956 33280
rect 21817 33222 21956 33224
rect 21817 33219 21883 33222
rect 21950 33220 21956 33222
rect 22020 33220 22026 33284
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 23105 33148 23171 33149
rect 23054 33084 23060 33148
rect 23124 33146 23171 33148
rect 23124 33144 23216 33146
rect 23166 33088 23216 33144
rect 23124 33086 23216 33088
rect 23124 33084 23171 33086
rect 23105 33083 23171 33084
rect 11973 32874 12039 32877
rect 18137 32874 18203 32877
rect 11973 32872 18203 32874
rect 11973 32816 11978 32872
rect 12034 32816 18142 32872
rect 18198 32816 18203 32872
rect 11973 32814 18203 32816
rect 11973 32811 12039 32814
rect 18137 32811 18203 32814
rect 22369 32738 22435 32741
rect 22502 32738 22508 32740
rect 22369 32736 22508 32738
rect 22369 32680 22374 32736
rect 22430 32680 22508 32736
rect 22369 32678 22508 32680
rect 22369 32675 22435 32678
rect 22502 32676 22508 32678
rect 22572 32676 22578 32740
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 21582 32540 21588 32604
rect 21652 32602 21658 32604
rect 22093 32602 22159 32605
rect 21652 32600 22159 32602
rect 21652 32544 22098 32600
rect 22154 32544 22159 32600
rect 21652 32542 22159 32544
rect 21652 32540 21658 32542
rect 22093 32539 22159 32542
rect 20478 32404 20484 32468
rect 20548 32466 20554 32468
rect 22645 32466 22711 32469
rect 20548 32464 22711 32466
rect 20548 32408 22650 32464
rect 22706 32408 22711 32464
rect 20548 32406 22711 32408
rect 20548 32404 20554 32406
rect 22645 32403 22711 32406
rect 23841 32330 23907 32333
rect 24485 32330 24551 32333
rect 22050 32328 24551 32330
rect 22050 32272 23846 32328
rect 23902 32272 24490 32328
rect 24546 32272 24551 32328
rect 22050 32270 24551 32272
rect 16573 32194 16639 32197
rect 20897 32194 20963 32197
rect 16573 32192 20963 32194
rect 16573 32136 16578 32192
rect 16634 32136 20902 32192
rect 20958 32136 20963 32192
rect 16573 32134 20963 32136
rect 16573 32131 16639 32134
rect 20897 32131 20963 32134
rect 4210 32128 4526 32129
rect 0 31968 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 11697 32058 11763 32061
rect 13169 32058 13235 32061
rect 11697 32056 13235 32058
rect 11697 32000 11702 32056
rect 11758 32000 13174 32056
rect 13230 32000 13235 32056
rect 11697 31998 13235 32000
rect 11697 31995 11763 31998
rect 13169 31995 13235 31998
rect 18229 32058 18295 32061
rect 18638 32058 18644 32060
rect 18229 32056 18644 32058
rect 18229 32000 18234 32056
rect 18290 32000 18644 32056
rect 18229 31998 18644 32000
rect 18229 31995 18295 31998
rect 18638 31996 18644 31998
rect 18708 31996 18714 32060
rect 16481 31922 16547 31925
rect 17585 31922 17651 31925
rect 22050 31922 22110 32270
rect 23841 32267 23907 32270
rect 24485 32267 24551 32270
rect 23013 32194 23079 32197
rect 23749 32194 23815 32197
rect 23013 32192 23815 32194
rect 23013 32136 23018 32192
rect 23074 32136 23754 32192
rect 23810 32136 23815 32192
rect 23013 32134 23815 32136
rect 23013 32131 23079 32134
rect 23749 32131 23815 32134
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 22737 32058 22803 32061
rect 23933 32058 23999 32061
rect 22737 32056 23999 32058
rect 22737 32000 22742 32056
rect 22798 32000 23938 32056
rect 23994 32000 23999 32056
rect 22737 31998 23999 32000
rect 22737 31995 22803 31998
rect 23933 31995 23999 31998
rect 38618 31968 39418 32088
rect 23381 31922 23447 31925
rect 27153 31924 27219 31925
rect 27102 31922 27108 31924
rect 16481 31920 22110 31922
rect 16481 31864 16486 31920
rect 16542 31864 17590 31920
rect 17646 31864 22110 31920
rect 16481 31862 22110 31864
rect 23246 31920 23447 31922
rect 23246 31864 23386 31920
rect 23442 31864 23447 31920
rect 23246 31862 23447 31864
rect 27062 31862 27108 31922
rect 27172 31920 27219 31924
rect 27214 31864 27219 31920
rect 16481 31859 16547 31862
rect 17585 31859 17651 31862
rect 19977 31786 20043 31789
rect 22185 31786 22251 31789
rect 19977 31784 22251 31786
rect 19977 31728 19982 31784
rect 20038 31728 22190 31784
rect 22246 31728 22251 31784
rect 19977 31726 22251 31728
rect 19977 31723 20043 31726
rect 22185 31723 22251 31726
rect 20437 31650 20503 31653
rect 21633 31650 21699 31653
rect 20437 31648 21699 31650
rect 20437 31592 20442 31648
rect 20498 31592 21638 31648
rect 21694 31592 21699 31648
rect 20437 31590 21699 31592
rect 20437 31587 20503 31590
rect 21633 31587 21699 31590
rect 21909 31650 21975 31653
rect 23246 31650 23306 31862
rect 23381 31859 23447 31862
rect 27102 31860 27108 31862
rect 27172 31860 27219 31864
rect 27153 31859 27219 31860
rect 25313 31650 25379 31653
rect 28349 31650 28415 31653
rect 21909 31648 28415 31650
rect 21909 31592 21914 31648
rect 21970 31592 25318 31648
rect 25374 31592 28354 31648
rect 28410 31592 28415 31648
rect 21909 31590 28415 31592
rect 21909 31587 21975 31590
rect 25313 31587 25379 31590
rect 28349 31587 28415 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 15193 31514 15259 31517
rect 19374 31514 19380 31516
rect 15193 31512 19380 31514
rect 15193 31456 15198 31512
rect 15254 31456 19380 31512
rect 15193 31454 19380 31456
rect 15193 31451 15259 31454
rect 19374 31452 19380 31454
rect 19444 31452 19450 31516
rect 21357 31514 21423 31517
rect 25865 31514 25931 31517
rect 21357 31512 25931 31514
rect 21357 31456 21362 31512
rect 21418 31456 25870 31512
rect 25926 31456 25931 31512
rect 21357 31454 25931 31456
rect 21357 31451 21423 31454
rect 25865 31451 25931 31454
rect 17769 31378 17835 31381
rect 20161 31378 20227 31381
rect 17769 31376 20227 31378
rect 17769 31320 17774 31376
rect 17830 31320 20166 31376
rect 20222 31320 20227 31376
rect 17769 31318 20227 31320
rect 17769 31315 17835 31318
rect 20161 31315 20227 31318
rect 28073 31242 28139 31245
rect 28809 31242 28875 31245
rect 28073 31240 28875 31242
rect 28073 31184 28078 31240
rect 28134 31184 28814 31240
rect 28870 31184 28875 31240
rect 28073 31182 28875 31184
rect 28073 31179 28139 31182
rect 28809 31179 28875 31182
rect 20529 31106 20595 31109
rect 28625 31106 28691 31109
rect 20529 31104 28691 31106
rect 20529 31048 20534 31104
rect 20590 31048 28630 31104
rect 28686 31048 28691 31104
rect 20529 31046 28691 31048
rect 20529 31043 20595 31046
rect 28625 31043 28691 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 17677 30970 17743 30973
rect 18965 30970 19031 30973
rect 17677 30968 19031 30970
rect 17677 30912 17682 30968
rect 17738 30912 18970 30968
rect 19026 30912 19031 30968
rect 17677 30910 19031 30912
rect 17677 30907 17743 30910
rect 18965 30907 19031 30910
rect 19374 30908 19380 30972
rect 19444 30970 19450 30972
rect 20713 30970 20779 30973
rect 19444 30968 20779 30970
rect 19444 30912 20718 30968
rect 20774 30912 20779 30968
rect 19444 30910 20779 30912
rect 19444 30908 19450 30910
rect 20713 30907 20779 30910
rect 18321 30834 18387 30837
rect 18689 30834 18755 30837
rect 18321 30832 18755 30834
rect 18321 30776 18326 30832
rect 18382 30776 18694 30832
rect 18750 30776 18755 30832
rect 18321 30774 18755 30776
rect 18321 30771 18387 30774
rect 18689 30771 18755 30774
rect 19006 30772 19012 30836
rect 19076 30834 19082 30836
rect 19149 30834 19215 30837
rect 19076 30832 19215 30834
rect 19076 30776 19154 30832
rect 19210 30776 19215 30832
rect 19076 30774 19215 30776
rect 19076 30772 19082 30774
rect 19149 30771 19215 30774
rect 15561 30562 15627 30565
rect 17861 30562 17927 30565
rect 15561 30560 17927 30562
rect 15561 30504 15566 30560
rect 15622 30504 17866 30560
rect 17922 30504 17927 30560
rect 15561 30502 17927 30504
rect 15561 30499 15627 30502
rect 17861 30499 17927 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 15285 30426 15351 30429
rect 18965 30426 19031 30429
rect 15285 30424 19031 30426
rect 15285 30368 15290 30424
rect 15346 30368 18970 30424
rect 19026 30368 19031 30424
rect 15285 30366 19031 30368
rect 15285 30363 15351 30366
rect 18965 30363 19031 30366
rect 22921 30426 22987 30429
rect 23606 30426 23612 30428
rect 22921 30424 23612 30426
rect 22921 30368 22926 30424
rect 22982 30368 23612 30424
rect 22921 30366 23612 30368
rect 22921 30363 22987 30366
rect 23606 30364 23612 30366
rect 23676 30364 23682 30428
rect 25865 30426 25931 30429
rect 27286 30426 27292 30428
rect 25865 30424 27292 30426
rect 25865 30368 25870 30424
rect 25926 30368 27292 30424
rect 25865 30366 27292 30368
rect 25865 30363 25931 30366
rect 27286 30364 27292 30366
rect 27356 30364 27362 30428
rect 9765 30290 9831 30293
rect 10961 30290 11027 30293
rect 9765 30288 11027 30290
rect 9765 30232 9770 30288
rect 9826 30232 10966 30288
rect 11022 30232 11027 30288
rect 9765 30230 11027 30232
rect 9765 30227 9831 30230
rect 10961 30227 11027 30230
rect 18689 30290 18755 30293
rect 23197 30290 23263 30293
rect 18689 30288 23263 30290
rect 18689 30232 18694 30288
rect 18750 30232 23202 30288
rect 23258 30232 23263 30288
rect 18689 30230 23263 30232
rect 18689 30227 18755 30230
rect 23197 30227 23263 30230
rect 15009 30154 15075 30157
rect 20713 30154 20779 30157
rect 15009 30152 20779 30154
rect 15009 30096 15014 30152
rect 15070 30096 20718 30152
rect 20774 30096 20779 30152
rect 15009 30094 20779 30096
rect 15009 30091 15075 30094
rect 20713 30091 20779 30094
rect 0 29928 800 30048
rect 15377 30018 15443 30021
rect 15837 30018 15903 30021
rect 18873 30018 18939 30021
rect 19149 30018 19215 30021
rect 19885 30018 19951 30021
rect 21449 30018 21515 30021
rect 22829 30018 22895 30021
rect 15377 30016 18939 30018
rect 15377 29960 15382 30016
rect 15438 29960 15842 30016
rect 15898 29960 18878 30016
rect 18934 29960 18939 30016
rect 15377 29958 18939 29960
rect 15377 29955 15443 29958
rect 15837 29955 15903 29958
rect 18873 29955 18939 29958
rect 19014 30016 22895 30018
rect 19014 29960 19154 30016
rect 19210 29960 19890 30016
rect 19946 29960 21454 30016
rect 21510 29960 22834 30016
rect 22890 29960 22895 30016
rect 19014 29958 22895 29960
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 13905 29882 13971 29885
rect 19014 29882 19074 29958
rect 19149 29955 19215 29958
rect 19885 29955 19951 29958
rect 21449 29955 21515 29958
rect 22829 29955 22895 29958
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 13905 29880 19074 29882
rect 13905 29824 13910 29880
rect 13966 29824 19074 29880
rect 13905 29822 19074 29824
rect 21265 29882 21331 29885
rect 21582 29882 21588 29884
rect 21265 29880 21588 29882
rect 21265 29824 21270 29880
rect 21326 29824 21588 29880
rect 21265 29822 21588 29824
rect 13905 29819 13971 29822
rect 21265 29819 21331 29822
rect 21582 29820 21588 29822
rect 21652 29820 21658 29884
rect 21817 29882 21883 29885
rect 25405 29882 25471 29885
rect 26509 29882 26575 29885
rect 21817 29880 26575 29882
rect 21817 29824 21822 29880
rect 21878 29824 25410 29880
rect 25466 29824 26514 29880
rect 26570 29824 26575 29880
rect 21817 29822 26575 29824
rect 21817 29819 21883 29822
rect 25405 29819 25471 29822
rect 26509 29819 26575 29822
rect 20161 29746 20227 29749
rect 26049 29746 26115 29749
rect 17174 29744 26115 29746
rect 17174 29688 20166 29744
rect 20222 29688 26054 29744
rect 26110 29688 26115 29744
rect 17174 29686 26115 29688
rect 12065 29610 12131 29613
rect 14181 29610 14247 29613
rect 17174 29610 17234 29686
rect 20161 29683 20227 29686
rect 26049 29683 26115 29686
rect 12065 29608 17234 29610
rect 12065 29552 12070 29608
rect 12126 29552 14186 29608
rect 14242 29552 17234 29608
rect 12065 29550 17234 29552
rect 19793 29610 19859 29613
rect 22093 29612 22159 29613
rect 20110 29610 20116 29612
rect 19793 29608 20116 29610
rect 19793 29552 19798 29608
rect 19854 29552 20116 29608
rect 19793 29550 20116 29552
rect 12065 29547 12131 29550
rect 14181 29547 14247 29550
rect 19793 29547 19859 29550
rect 20110 29548 20116 29550
rect 20180 29548 20186 29612
rect 22093 29608 22140 29612
rect 22204 29610 22210 29612
rect 25773 29610 25839 29613
rect 22204 29608 25839 29610
rect 22093 29552 22098 29608
rect 22204 29552 25778 29608
rect 25834 29552 25839 29608
rect 22093 29548 22140 29552
rect 22204 29550 25839 29552
rect 22204 29548 22210 29550
rect 22093 29547 22159 29548
rect 25773 29547 25839 29550
rect 19977 29474 20043 29477
rect 23105 29474 23171 29477
rect 19977 29472 23171 29474
rect 19977 29416 19982 29472
rect 20038 29416 23110 29472
rect 23166 29416 23171 29472
rect 19977 29414 23171 29416
rect 19977 29411 20043 29414
rect 23105 29411 23171 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 15561 29338 15627 29341
rect 18873 29338 18939 29341
rect 15561 29336 18939 29338
rect 15561 29280 15566 29336
rect 15622 29280 18878 29336
rect 18934 29280 18939 29336
rect 15561 29278 18939 29280
rect 15561 29275 15627 29278
rect 18873 29275 18939 29278
rect 38618 29248 39418 29368
rect 16205 29202 16271 29205
rect 19057 29202 19123 29205
rect 16205 29200 19123 29202
rect 16205 29144 16210 29200
rect 16266 29144 19062 29200
rect 19118 29144 19123 29200
rect 16205 29142 19123 29144
rect 16205 29139 16271 29142
rect 19057 29139 19123 29142
rect 13353 29068 13419 29069
rect 13302 29066 13308 29068
rect 13262 29006 13308 29066
rect 13372 29064 13419 29068
rect 13414 29008 13419 29064
rect 13302 29004 13308 29006
rect 13372 29004 13419 29008
rect 13353 29003 13419 29004
rect 18045 29066 18111 29069
rect 18454 29066 18460 29068
rect 18045 29064 18460 29066
rect 18045 29008 18050 29064
rect 18106 29008 18460 29064
rect 18045 29006 18460 29008
rect 18045 29003 18111 29006
rect 18454 29004 18460 29006
rect 18524 29004 18530 29068
rect 18781 29066 18847 29069
rect 19006 29066 19012 29068
rect 18781 29064 19012 29066
rect 18781 29008 18786 29064
rect 18842 29008 19012 29064
rect 18781 29006 19012 29008
rect 18781 29003 18847 29006
rect 19006 29004 19012 29006
rect 19076 29004 19082 29068
rect 31569 29066 31635 29069
rect 33041 29066 33107 29069
rect 31569 29064 33107 29066
rect 31569 29008 31574 29064
rect 31630 29008 33046 29064
rect 33102 29008 33107 29064
rect 31569 29006 33107 29008
rect 31569 29003 31635 29006
rect 33041 29003 33107 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 18413 28794 18479 28797
rect 22921 28794 22987 28797
rect 18413 28792 22987 28794
rect 18413 28736 18418 28792
rect 18474 28736 22926 28792
rect 22982 28736 22987 28792
rect 18413 28734 22987 28736
rect 18413 28731 18479 28734
rect 22921 28731 22987 28734
rect 22502 28596 22508 28660
rect 22572 28658 22578 28660
rect 23749 28658 23815 28661
rect 22572 28656 23815 28658
rect 22572 28600 23754 28656
rect 23810 28600 23815 28656
rect 22572 28598 23815 28600
rect 22572 28596 22578 28598
rect 23749 28595 23815 28598
rect 24669 28658 24735 28661
rect 29085 28658 29151 28661
rect 24669 28656 29151 28658
rect 24669 28600 24674 28656
rect 24730 28600 29090 28656
rect 29146 28600 29151 28656
rect 24669 28598 29151 28600
rect 24669 28595 24735 28598
rect 29085 28595 29151 28598
rect 15469 28522 15535 28525
rect 20294 28522 20300 28524
rect 15469 28520 20300 28522
rect 15469 28464 15474 28520
rect 15530 28464 20300 28520
rect 15469 28462 20300 28464
rect 15469 28459 15535 28462
rect 20294 28460 20300 28462
rect 20364 28522 20370 28524
rect 22737 28522 22803 28525
rect 20364 28520 22803 28522
rect 20364 28464 22742 28520
rect 22798 28464 22803 28520
rect 20364 28462 22803 28464
rect 20364 28460 20370 28462
rect 22737 28459 22803 28462
rect 28993 28522 29059 28525
rect 31385 28522 31451 28525
rect 28993 28520 31451 28522
rect 28993 28464 28998 28520
rect 29054 28464 31390 28520
rect 31446 28464 31451 28520
rect 28993 28462 31451 28464
rect 28993 28459 29059 28462
rect 31385 28459 31451 28462
rect 22277 28386 22343 28389
rect 22921 28386 22987 28389
rect 22277 28384 22987 28386
rect 22277 28328 22282 28384
rect 22338 28328 22926 28384
rect 22982 28328 22987 28384
rect 22277 28326 22987 28328
rect 22277 28323 22343 28326
rect 22921 28323 22987 28326
rect 25497 28386 25563 28389
rect 26969 28386 27035 28389
rect 25497 28384 27035 28386
rect 25497 28328 25502 28384
rect 25558 28328 26974 28384
rect 27030 28328 27035 28384
rect 25497 28326 27035 28328
rect 25497 28323 25563 28326
rect 26969 28323 27035 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 16113 28114 16179 28117
rect 22645 28114 22711 28117
rect 23054 28114 23060 28116
rect 16113 28112 23060 28114
rect 16113 28056 16118 28112
rect 16174 28056 22650 28112
rect 22706 28056 23060 28112
rect 16113 28054 23060 28056
rect 16113 28051 16179 28054
rect 22645 28051 22711 28054
rect 23054 28052 23060 28054
rect 23124 28052 23130 28116
rect 28993 28114 29059 28117
rect 30005 28114 30071 28117
rect 28993 28112 30071 28114
rect 28993 28056 28998 28112
rect 29054 28056 30010 28112
rect 30066 28056 30071 28112
rect 28993 28054 30071 28056
rect 28993 28051 29059 28054
rect 30005 28051 30071 28054
rect 15377 27978 15443 27981
rect 22553 27978 22619 27981
rect 15377 27976 22619 27978
rect 15377 27920 15382 27976
rect 15438 27920 22558 27976
rect 22614 27920 22619 27976
rect 15377 27918 22619 27920
rect 15377 27915 15443 27918
rect 22553 27915 22619 27918
rect 19517 27842 19583 27845
rect 21766 27842 21772 27844
rect 19517 27840 21772 27842
rect 19517 27784 19522 27840
rect 19578 27784 21772 27840
rect 19517 27782 21772 27784
rect 19517 27779 19583 27782
rect 21766 27780 21772 27782
rect 21836 27780 21842 27844
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 20989 27708 21055 27709
rect 20989 27704 21036 27708
rect 21100 27706 21106 27708
rect 20989 27648 20994 27704
rect 20989 27644 21036 27648
rect 21100 27646 21146 27706
rect 21100 27644 21106 27646
rect 20989 27643 21055 27644
rect 14549 27570 14615 27573
rect 17401 27570 17467 27573
rect 14549 27568 17467 27570
rect 14549 27512 14554 27568
rect 14610 27512 17406 27568
rect 17462 27512 17467 27568
rect 14549 27510 17467 27512
rect 14549 27507 14615 27510
rect 17401 27507 17467 27510
rect 19425 27570 19491 27573
rect 20805 27570 20871 27573
rect 23565 27570 23631 27573
rect 19425 27568 23631 27570
rect 19425 27512 19430 27568
rect 19486 27512 20810 27568
rect 20866 27512 23570 27568
rect 23626 27512 23631 27568
rect 19425 27510 23631 27512
rect 19425 27507 19491 27510
rect 20805 27507 20871 27510
rect 23565 27507 23631 27510
rect 20529 27434 20595 27437
rect 22093 27434 22159 27437
rect 20529 27432 22159 27434
rect 20529 27376 20534 27432
rect 20590 27376 22098 27432
rect 22154 27376 22159 27432
rect 20529 27374 22159 27376
rect 20529 27371 20595 27374
rect 22093 27371 22159 27374
rect 0 27298 800 27328
rect 4061 27298 4127 27301
rect 14181 27300 14247 27301
rect 14181 27298 14228 27300
rect 0 27296 4127 27298
rect 0 27240 4066 27296
rect 4122 27240 4127 27296
rect 0 27238 4127 27240
rect 14136 27296 14228 27298
rect 14136 27240 14186 27296
rect 14136 27238 14228 27240
rect 0 27208 800 27238
rect 4061 27235 4127 27238
rect 14181 27236 14228 27238
rect 14292 27236 14298 27300
rect 14181 27235 14247 27236
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 38618 27208 39418 27328
rect 19570 27167 19886 27168
rect 12801 27162 12867 27165
rect 15377 27162 15443 27165
rect 12801 27160 15443 27162
rect 12801 27104 12806 27160
rect 12862 27104 15382 27160
rect 15438 27104 15443 27160
rect 12801 27102 15443 27104
rect 12801 27099 12867 27102
rect 15377 27099 15443 27102
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 14825 26482 14891 26485
rect 19333 26482 19399 26485
rect 20529 26482 20595 26485
rect 14825 26480 20595 26482
rect 14825 26424 14830 26480
rect 14886 26424 19338 26480
rect 19394 26424 20534 26480
rect 20590 26424 20595 26480
rect 14825 26422 20595 26424
rect 14825 26419 14891 26422
rect 19333 26419 19399 26422
rect 20529 26419 20595 26422
rect 20897 26482 20963 26485
rect 22134 26482 22140 26484
rect 20897 26480 22140 26482
rect 20897 26424 20902 26480
rect 20958 26424 22140 26480
rect 20897 26422 22140 26424
rect 20897 26419 20963 26422
rect 22134 26420 22140 26422
rect 22204 26420 22210 26484
rect 8293 26346 8359 26349
rect 26049 26346 26115 26349
rect 8293 26344 26115 26346
rect 8293 26288 8298 26344
rect 8354 26288 26054 26344
rect 26110 26288 26115 26344
rect 8293 26286 26115 26288
rect 8293 26283 8359 26286
rect 26049 26283 26115 26286
rect 30741 26346 30807 26349
rect 33685 26346 33751 26349
rect 30741 26344 33751 26346
rect 30741 26288 30746 26344
rect 30802 26288 33690 26344
rect 33746 26288 33751 26344
rect 30741 26286 33751 26288
rect 30741 26283 30807 26286
rect 33685 26283 33751 26286
rect 18597 26210 18663 26213
rect 19374 26210 19380 26212
rect 18597 26208 19380 26210
rect 18597 26152 18602 26208
rect 18658 26152 19380 26208
rect 18597 26150 19380 26152
rect 18597 26147 18663 26150
rect 19374 26148 19380 26150
rect 19444 26148 19450 26212
rect 20805 26210 20871 26213
rect 24761 26210 24827 26213
rect 20805 26208 24827 26210
rect 20805 26152 20810 26208
rect 20866 26152 24766 26208
rect 24822 26152 24827 26208
rect 20805 26150 24827 26152
rect 20805 26147 20871 26150
rect 24761 26147 24827 26150
rect 25313 26210 25379 26213
rect 25446 26210 25452 26212
rect 25313 26208 25452 26210
rect 25313 26152 25318 26208
rect 25374 26152 25452 26208
rect 25313 26150 25452 26152
rect 25313 26147 25379 26150
rect 25446 26148 25452 26150
rect 25516 26148 25522 26212
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 25405 26074 25471 26077
rect 27797 26074 27863 26077
rect 25405 26072 27863 26074
rect 25405 26016 25410 26072
rect 25466 26016 27802 26072
rect 27858 26016 27863 26072
rect 25405 26014 27863 26016
rect 25405 26011 25471 26014
rect 27797 26011 27863 26014
rect 23197 25938 23263 25941
rect 26877 25938 26943 25941
rect 23197 25936 26943 25938
rect 23197 25880 23202 25936
rect 23258 25880 26882 25936
rect 26938 25880 26943 25936
rect 23197 25878 26943 25880
rect 23197 25875 23263 25878
rect 26877 25875 26943 25878
rect 19701 25802 19767 25805
rect 24117 25802 24183 25805
rect 19701 25800 24183 25802
rect 19701 25744 19706 25800
rect 19762 25744 24122 25800
rect 24178 25744 24183 25800
rect 19701 25742 24183 25744
rect 19701 25739 19767 25742
rect 24117 25739 24183 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19701 25530 19767 25533
rect 21173 25530 21239 25533
rect 19701 25528 21239 25530
rect 19701 25472 19706 25528
rect 19762 25472 21178 25528
rect 21234 25472 21239 25528
rect 19701 25470 21239 25472
rect 19701 25467 19767 25470
rect 21173 25467 21239 25470
rect 13721 25394 13787 25397
rect 24577 25394 24643 25397
rect 13721 25392 24643 25394
rect 13721 25336 13726 25392
rect 13782 25336 24582 25392
rect 24638 25336 24643 25392
rect 13721 25334 24643 25336
rect 13721 25331 13787 25334
rect 24577 25331 24643 25334
rect 0 25258 800 25288
rect 0 25168 858 25258
rect 11830 25196 11836 25260
rect 11900 25258 11906 25260
rect 12065 25258 12131 25261
rect 11900 25256 12131 25258
rect 11900 25200 12070 25256
rect 12126 25200 12131 25256
rect 11900 25198 12131 25200
rect 11900 25196 11906 25198
rect 12065 25195 12131 25198
rect 16573 25258 16639 25261
rect 24761 25258 24827 25261
rect 16573 25256 24827 25258
rect 16573 25200 16578 25256
rect 16634 25200 24766 25256
rect 24822 25200 24827 25256
rect 16573 25198 24827 25200
rect 16573 25195 16639 25198
rect 24761 25195 24827 25198
rect 38618 25168 39418 25288
rect 798 24986 858 25168
rect 20253 25124 20319 25125
rect 20253 25122 20300 25124
rect 20208 25120 20300 25122
rect 20208 25064 20258 25120
rect 20208 25062 20300 25064
rect 20253 25060 20300 25062
rect 20364 25060 20370 25124
rect 22369 25122 22435 25125
rect 25405 25122 25471 25125
rect 22369 25120 25471 25122
rect 22369 25064 22374 25120
rect 22430 25064 25410 25120
rect 25466 25064 25471 25120
rect 22369 25062 25471 25064
rect 20253 25059 20319 25060
rect 22369 25059 22435 25062
rect 25405 25059 25471 25062
rect 25681 25122 25747 25125
rect 28625 25122 28691 25125
rect 25681 25120 28691 25122
rect 25681 25064 25686 25120
rect 25742 25064 28630 25120
rect 28686 25064 28691 25120
rect 25681 25062 28691 25064
rect 25681 25059 25747 25062
rect 28625 25059 28691 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 1577 24986 1643 24989
rect 20529 24986 20595 24989
rect 798 24984 1643 24986
rect 798 24928 1582 24984
rect 1638 24928 1643 24984
rect 798 24926 1643 24928
rect 1577 24923 1643 24926
rect 20302 24984 20595 24986
rect 20302 24928 20534 24984
rect 20590 24928 20595 24984
rect 20302 24926 20595 24928
rect 13169 24850 13235 24853
rect 15561 24850 15627 24853
rect 13169 24848 15627 24850
rect 13169 24792 13174 24848
rect 13230 24792 15566 24848
rect 15622 24792 15627 24848
rect 13169 24790 15627 24792
rect 13169 24787 13235 24790
rect 15561 24787 15627 24790
rect 15929 24850 15995 24853
rect 20302 24850 20362 24926
rect 20529 24923 20595 24926
rect 22277 24986 22343 24989
rect 24577 24986 24643 24989
rect 22277 24984 24643 24986
rect 22277 24928 22282 24984
rect 22338 24928 24582 24984
rect 24638 24928 24643 24984
rect 22277 24926 24643 24928
rect 22277 24923 22343 24926
rect 24577 24923 24643 24926
rect 15929 24848 20362 24850
rect 15929 24792 15934 24848
rect 15990 24792 20362 24848
rect 15929 24790 20362 24792
rect 20437 24850 20503 24853
rect 23105 24850 23171 24853
rect 27061 24852 27127 24853
rect 27061 24850 27108 24852
rect 20437 24848 23171 24850
rect 20437 24792 20442 24848
rect 20498 24792 23110 24848
rect 23166 24792 23171 24848
rect 20437 24790 23171 24792
rect 27016 24848 27108 24850
rect 27016 24792 27066 24848
rect 27016 24790 27108 24792
rect 15929 24787 15995 24790
rect 20437 24787 20503 24790
rect 23105 24787 23171 24790
rect 27061 24788 27108 24790
rect 27172 24788 27178 24852
rect 27061 24787 27127 24788
rect 17861 24714 17927 24717
rect 22185 24714 22251 24717
rect 22829 24714 22895 24717
rect 17861 24712 22895 24714
rect 17861 24656 17866 24712
rect 17922 24656 22190 24712
rect 22246 24656 22834 24712
rect 22890 24656 22895 24712
rect 17861 24654 22895 24656
rect 17861 24651 17927 24654
rect 22185 24651 22251 24654
rect 22829 24651 22895 24654
rect 20621 24578 20687 24581
rect 24853 24578 24919 24581
rect 26049 24578 26115 24581
rect 20621 24576 26115 24578
rect 20621 24520 20626 24576
rect 20682 24520 24858 24576
rect 24914 24520 26054 24576
rect 26110 24520 26115 24576
rect 20621 24518 26115 24520
rect 20621 24515 20687 24518
rect 24853 24515 24919 24518
rect 26049 24515 26115 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 17125 24442 17191 24445
rect 24393 24442 24459 24445
rect 17125 24440 24459 24442
rect 17125 24384 17130 24440
rect 17186 24384 24398 24440
rect 24454 24384 24459 24440
rect 17125 24382 24459 24384
rect 17125 24379 17191 24382
rect 24393 24379 24459 24382
rect 12709 24306 12775 24309
rect 14089 24306 14155 24309
rect 12709 24304 14155 24306
rect 12709 24248 12714 24304
rect 12770 24248 14094 24304
rect 14150 24248 14155 24304
rect 12709 24246 14155 24248
rect 12709 24243 12775 24246
rect 14089 24243 14155 24246
rect 22185 24306 22251 24309
rect 26601 24306 26667 24309
rect 22185 24304 26667 24306
rect 22185 24248 22190 24304
rect 22246 24248 26606 24304
rect 26662 24248 26667 24304
rect 22185 24246 26667 24248
rect 22185 24243 22251 24246
rect 26601 24243 26667 24246
rect 15837 24170 15903 24173
rect 20621 24170 20687 24173
rect 15837 24168 20687 24170
rect 15837 24112 15842 24168
rect 15898 24112 20626 24168
rect 20682 24112 20687 24168
rect 15837 24110 20687 24112
rect 15837 24107 15903 24110
rect 20621 24107 20687 24110
rect 22461 24170 22527 24173
rect 24945 24170 25011 24173
rect 22461 24168 25011 24170
rect 22461 24112 22466 24168
rect 22522 24112 24950 24168
rect 25006 24112 25011 24168
rect 22461 24110 25011 24112
rect 22461 24107 22527 24110
rect 24945 24107 25011 24110
rect 15837 24034 15903 24037
rect 18597 24034 18663 24037
rect 15837 24032 18663 24034
rect 15837 23976 15842 24032
rect 15898 23976 18602 24032
rect 18658 23976 18663 24032
rect 15837 23974 18663 23976
rect 15837 23971 15903 23974
rect 18597 23971 18663 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 13353 23898 13419 23901
rect 13905 23898 13971 23901
rect 13353 23896 13971 23898
rect 13353 23840 13358 23896
rect 13414 23840 13910 23896
rect 13966 23840 13971 23896
rect 13353 23838 13971 23840
rect 13353 23835 13419 23838
rect 13905 23835 13971 23838
rect 15561 23762 15627 23765
rect 18505 23762 18571 23765
rect 15561 23760 18571 23762
rect 15561 23704 15566 23760
rect 15622 23704 18510 23760
rect 18566 23704 18571 23760
rect 15561 23702 18571 23704
rect 15561 23699 15627 23702
rect 18505 23699 18571 23702
rect 20713 23762 20779 23765
rect 20713 23760 22708 23762
rect 20713 23704 20718 23760
rect 20774 23704 22708 23760
rect 20713 23702 22708 23704
rect 20713 23699 20779 23702
rect 22648 23629 22708 23702
rect 15837 23626 15903 23629
rect 20989 23626 21055 23629
rect 15837 23624 21055 23626
rect 15837 23568 15842 23624
rect 15898 23568 20994 23624
rect 21050 23568 21055 23624
rect 15837 23566 21055 23568
rect 15837 23563 15903 23566
rect 20989 23563 21055 23566
rect 22645 23624 22711 23629
rect 22645 23568 22650 23624
rect 22706 23568 22711 23624
rect 22645 23563 22711 23568
rect 25773 23626 25839 23629
rect 27470 23626 27476 23628
rect 25773 23624 27476 23626
rect 25773 23568 25778 23624
rect 25834 23568 27476 23624
rect 25773 23566 27476 23568
rect 25773 23563 25839 23566
rect 27470 23564 27476 23566
rect 27540 23564 27546 23628
rect 16481 23492 16547 23493
rect 16430 23490 16436 23492
rect 16390 23430 16436 23490
rect 16500 23488 16547 23492
rect 16542 23432 16547 23488
rect 16430 23428 16436 23430
rect 16500 23428 16547 23432
rect 16481 23427 16547 23428
rect 21081 23490 21147 23493
rect 26969 23490 27035 23493
rect 21081 23488 27035 23490
rect 21081 23432 21086 23488
rect 21142 23432 26974 23488
rect 27030 23432 27035 23488
rect 21081 23430 27035 23432
rect 21081 23427 21147 23430
rect 26969 23427 27035 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 21357 23354 21423 23357
rect 27245 23354 27311 23357
rect 21357 23352 27311 23354
rect 21357 23296 21362 23352
rect 21418 23296 27250 23352
rect 27306 23296 27311 23352
rect 21357 23294 27311 23296
rect 21357 23291 21423 23294
rect 27245 23291 27311 23294
rect 0 23128 800 23248
rect 20437 23218 20503 23221
rect 20897 23218 20963 23221
rect 20437 23216 20963 23218
rect 20437 23160 20442 23216
rect 20498 23160 20902 23216
rect 20958 23160 20963 23216
rect 20437 23158 20963 23160
rect 20437 23155 20503 23158
rect 20897 23155 20963 23158
rect 4613 23082 4679 23085
rect 7833 23082 7899 23085
rect 4613 23080 7899 23082
rect 4613 23024 4618 23080
rect 4674 23024 7838 23080
rect 7894 23024 7899 23080
rect 4613 23022 7899 23024
rect 4613 23019 4679 23022
rect 7833 23019 7899 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 21817 22810 21883 22813
rect 27061 22810 27127 22813
rect 21817 22808 27127 22810
rect 21817 22752 21822 22808
rect 21878 22752 27066 22808
rect 27122 22752 27127 22808
rect 21817 22750 27127 22752
rect 21817 22747 21883 22750
rect 27061 22747 27127 22750
rect 3049 22674 3115 22677
rect 4061 22674 4127 22677
rect 3049 22672 4127 22674
rect 3049 22616 3054 22672
rect 3110 22616 4066 22672
rect 4122 22616 4127 22672
rect 3049 22614 4127 22616
rect 3049 22611 3115 22614
rect 4061 22611 4127 22614
rect 7833 22674 7899 22677
rect 27245 22674 27311 22677
rect 7833 22672 27311 22674
rect 7833 22616 7838 22672
rect 7894 22616 27250 22672
rect 27306 22616 27311 22672
rect 7833 22614 27311 22616
rect 7833 22611 7899 22614
rect 27245 22611 27311 22614
rect 6637 22538 6703 22541
rect 7097 22538 7163 22541
rect 8477 22538 8543 22541
rect 6637 22536 8543 22538
rect 6637 22480 6642 22536
rect 6698 22480 7102 22536
rect 7158 22480 8482 22536
rect 8538 22480 8543 22536
rect 6637 22478 8543 22480
rect 6637 22475 6703 22478
rect 7097 22475 7163 22478
rect 8477 22475 8543 22478
rect 21173 22538 21239 22541
rect 22001 22538 22067 22541
rect 21173 22536 22067 22538
rect 21173 22480 21178 22536
rect 21234 22480 22006 22536
rect 22062 22480 22067 22536
rect 21173 22478 22067 22480
rect 21173 22475 21239 22478
rect 22001 22475 22067 22478
rect 23974 22476 23980 22540
rect 24044 22476 24050 22540
rect 37825 22538 37891 22541
rect 38618 22538 39418 22568
rect 37825 22536 39418 22538
rect 37825 22480 37830 22536
rect 37886 22480 39418 22536
rect 37825 22478 39418 22480
rect 22461 22402 22527 22405
rect 23982 22402 24042 22476
rect 37825 22475 37891 22478
rect 38618 22448 39418 22478
rect 22461 22400 24042 22402
rect 22461 22344 22466 22400
rect 22522 22344 24042 22400
rect 22461 22342 24042 22344
rect 22461 22339 22527 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 20529 22266 20595 22269
rect 22553 22266 22619 22269
rect 20529 22264 22619 22266
rect 20529 22208 20534 22264
rect 20590 22208 22558 22264
rect 22614 22208 22619 22264
rect 20529 22206 22619 22208
rect 20529 22203 20595 22206
rect 22553 22203 22619 22206
rect 3969 22130 4035 22133
rect 8293 22130 8359 22133
rect 3969 22128 8359 22130
rect 3969 22072 3974 22128
rect 4030 22072 8298 22128
rect 8354 22072 8359 22128
rect 3969 22070 8359 22072
rect 3969 22067 4035 22070
rect 8293 22067 8359 22070
rect 9305 22130 9371 22133
rect 24853 22130 24919 22133
rect 9305 22128 24919 22130
rect 9305 22072 9310 22128
rect 9366 22072 24858 22128
rect 24914 22072 24919 22128
rect 9305 22070 24919 22072
rect 9305 22067 9371 22070
rect 24853 22067 24919 22070
rect 31661 22130 31727 22133
rect 32673 22130 32739 22133
rect 31661 22128 32739 22130
rect 31661 22072 31666 22128
rect 31722 22072 32678 22128
rect 32734 22072 32739 22128
rect 31661 22070 32739 22072
rect 31661 22067 31727 22070
rect 32673 22067 32739 22070
rect 12249 21996 12315 21997
rect 12198 21932 12204 21996
rect 12268 21994 12315 21996
rect 23105 21994 23171 21997
rect 12268 21992 12360 21994
rect 12310 21936 12360 21992
rect 12268 21934 12360 21936
rect 17174 21992 23171 21994
rect 17174 21936 23110 21992
rect 23166 21936 23171 21992
rect 17174 21934 23171 21936
rect 12268 21932 12315 21934
rect 12249 21931 12315 21932
rect 4981 21858 5047 21861
rect 17174 21858 17234 21934
rect 23105 21931 23171 21934
rect 4981 21856 17234 21858
rect 4981 21800 4986 21856
rect 5042 21800 17234 21856
rect 4981 21798 17234 21800
rect 4981 21795 5047 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 13353 21722 13419 21725
rect 13486 21722 13492 21724
rect 13353 21720 13492 21722
rect 13353 21664 13358 21720
rect 13414 21664 13492 21720
rect 13353 21662 13492 21664
rect 13353 21659 13419 21662
rect 13486 21660 13492 21662
rect 13556 21660 13562 21724
rect 23013 21722 23079 21725
rect 23422 21722 23428 21724
rect 23013 21720 23428 21722
rect 23013 21664 23018 21720
rect 23074 21664 23428 21720
rect 23013 21662 23428 21664
rect 23013 21659 23079 21662
rect 23422 21660 23428 21662
rect 23492 21660 23498 21724
rect 2405 21586 2471 21589
rect 23933 21586 23999 21589
rect 2405 21584 23999 21586
rect 2405 21528 2410 21584
rect 2466 21528 23938 21584
rect 23994 21528 23999 21584
rect 2405 21526 23999 21528
rect 2405 21523 2471 21526
rect 23933 21523 23999 21526
rect 25957 21586 26023 21589
rect 36721 21586 36787 21589
rect 25957 21584 36787 21586
rect 25957 21528 25962 21584
rect 26018 21528 36726 21584
rect 36782 21528 36787 21584
rect 25957 21526 36787 21528
rect 25957 21523 26023 21526
rect 36721 21523 36787 21526
rect 7005 21450 7071 21453
rect 25405 21450 25471 21453
rect 7005 21448 25471 21450
rect 7005 21392 7010 21448
rect 7066 21392 25410 21448
rect 25466 21392 25471 21448
rect 7005 21390 25471 21392
rect 7005 21387 7071 21390
rect 25405 21387 25471 21390
rect 11881 21314 11947 21317
rect 25773 21314 25839 21317
rect 11881 21312 25839 21314
rect 11881 21256 11886 21312
rect 11942 21256 25778 21312
rect 25834 21256 25839 21312
rect 11881 21254 25839 21256
rect 11881 21251 11947 21254
rect 25773 21251 25839 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 25405 20906 25471 20909
rect 9814 20904 25471 20906
rect 9814 20848 25410 20904
rect 25466 20848 25471 20904
rect 9814 20846 25471 20848
rect 9029 20772 9095 20773
rect 9029 20770 9076 20772
rect 8984 20768 9076 20770
rect 8984 20712 9034 20768
rect 8984 20710 9076 20712
rect 9029 20708 9076 20710
rect 9140 20708 9146 20772
rect 9029 20707 9095 20708
rect 2221 20634 2287 20637
rect 9814 20634 9874 20846
rect 25405 20843 25471 20846
rect 10317 20772 10383 20773
rect 10317 20770 10364 20772
rect 10272 20768 10364 20770
rect 10272 20712 10322 20768
rect 10272 20710 10364 20712
rect 10317 20708 10364 20710
rect 10428 20708 10434 20772
rect 10317 20707 10383 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 25589 20636 25655 20637
rect 25589 20634 25636 20636
rect 2221 20632 9874 20634
rect 2221 20576 2226 20632
rect 2282 20576 9874 20632
rect 2221 20574 9874 20576
rect 25544 20632 25636 20634
rect 25544 20576 25594 20632
rect 25544 20574 25636 20576
rect 2221 20571 2287 20574
rect 25589 20572 25636 20574
rect 25700 20572 25706 20636
rect 25589 20571 25655 20572
rect 0 20498 800 20528
rect 933 20498 999 20501
rect 0 20496 999 20498
rect 0 20440 938 20496
rect 994 20440 999 20496
rect 0 20438 999 20440
rect 0 20408 800 20438
rect 933 20435 999 20438
rect 4061 20498 4127 20501
rect 6637 20498 6703 20501
rect 25405 20498 25471 20501
rect 4061 20496 25471 20498
rect 4061 20440 4066 20496
rect 4122 20440 6642 20496
rect 6698 20440 25410 20496
rect 25466 20440 25471 20496
rect 4061 20438 25471 20440
rect 4061 20435 4127 20438
rect 6637 20435 6703 20438
rect 25405 20435 25471 20438
rect 38377 20498 38443 20501
rect 38618 20498 39418 20528
rect 38377 20496 39418 20498
rect 38377 20440 38382 20496
rect 38438 20440 39418 20496
rect 38377 20438 39418 20440
rect 38377 20435 38443 20438
rect 38618 20408 39418 20438
rect 11605 20362 11671 20365
rect 12157 20362 12223 20365
rect 23381 20362 23447 20365
rect 11605 20360 23447 20362
rect 11605 20304 11610 20360
rect 11666 20304 12162 20360
rect 12218 20304 23386 20360
rect 23442 20304 23447 20360
rect 11605 20302 23447 20304
rect 11605 20299 11671 20302
rect 12157 20299 12223 20302
rect 23381 20299 23447 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 14273 20090 14339 20093
rect 17861 20090 17927 20093
rect 14273 20088 17927 20090
rect 14273 20032 14278 20088
rect 14334 20032 17866 20088
rect 17922 20032 17927 20088
rect 14273 20030 17927 20032
rect 14273 20027 14339 20030
rect 17861 20027 17927 20030
rect 13813 19954 13879 19957
rect 20478 19954 20484 19956
rect 13813 19952 20484 19954
rect 13813 19896 13818 19952
rect 13874 19896 20484 19952
rect 13813 19894 20484 19896
rect 13813 19891 13879 19894
rect 20478 19892 20484 19894
rect 20548 19954 20554 19956
rect 22185 19954 22251 19957
rect 20548 19952 22251 19954
rect 20548 19896 22190 19952
rect 22246 19896 22251 19952
rect 20548 19894 22251 19896
rect 20548 19892 20554 19894
rect 22185 19891 22251 19894
rect 8661 19818 8727 19821
rect 25773 19818 25839 19821
rect 8661 19816 25839 19818
rect 8661 19760 8666 19816
rect 8722 19760 25778 19816
rect 25834 19760 25839 19816
rect 8661 19758 25839 19760
rect 8661 19755 8727 19758
rect 25773 19755 25839 19758
rect 16849 19682 16915 19685
rect 17861 19682 17927 19685
rect 16849 19680 17927 19682
rect 16849 19624 16854 19680
rect 16910 19624 17866 19680
rect 17922 19624 17927 19680
rect 16849 19622 17927 19624
rect 16849 19619 16915 19622
rect 17861 19619 17927 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 13629 19546 13695 19549
rect 16573 19546 16639 19549
rect 13629 19544 16639 19546
rect 13629 19488 13634 19544
rect 13690 19488 16578 19544
rect 16634 19488 16639 19544
rect 13629 19486 16639 19488
rect 13629 19483 13695 19486
rect 16573 19483 16639 19486
rect 20161 19546 20227 19549
rect 24209 19546 24275 19549
rect 20161 19544 24275 19546
rect 20161 19488 20166 19544
rect 20222 19488 24214 19544
rect 24270 19488 24275 19544
rect 20161 19486 24275 19488
rect 20161 19483 20227 19486
rect 24209 19483 24275 19486
rect 23933 19410 23999 19413
rect 12390 19408 23999 19410
rect 12390 19352 23938 19408
rect 23994 19352 23999 19408
rect 12390 19350 23999 19352
rect 11881 19274 11947 19277
rect 12390 19274 12450 19350
rect 23933 19347 23999 19350
rect 28901 19350 28967 19353
rect 28901 19348 29010 19350
rect 28901 19292 28906 19348
rect 28962 19292 29010 19348
rect 28901 19287 29010 19292
rect 11881 19272 12450 19274
rect 11881 19216 11886 19272
rect 11942 19216 12450 19272
rect 11881 19214 12450 19216
rect 14917 19274 14983 19277
rect 22645 19274 22711 19277
rect 14917 19272 22711 19274
rect 14917 19216 14922 19272
rect 14978 19216 22650 19272
rect 22706 19216 22711 19272
rect 14917 19214 22711 19216
rect 11881 19211 11947 19214
rect 14917 19211 14983 19214
rect 22645 19211 22711 19214
rect 23013 19274 23079 19277
rect 25681 19274 25747 19277
rect 23013 19272 25747 19274
rect 23013 19216 23018 19272
rect 23074 19216 25686 19272
rect 25742 19216 25747 19272
rect 23013 19214 25747 19216
rect 23013 19211 23079 19214
rect 25681 19211 25747 19214
rect 28950 19141 29010 19287
rect 10409 19138 10475 19141
rect 12709 19138 12775 19141
rect 10409 19136 12775 19138
rect 10409 19080 10414 19136
rect 10470 19080 12714 19136
rect 12770 19080 12775 19136
rect 10409 19078 12775 19080
rect 10409 19075 10475 19078
rect 12709 19075 12775 19078
rect 12985 19138 13051 19141
rect 13629 19138 13695 19141
rect 12985 19136 13695 19138
rect 12985 19080 12990 19136
rect 13046 19080 13634 19136
rect 13690 19080 13695 19136
rect 12985 19078 13695 19080
rect 12985 19075 13051 19078
rect 13629 19075 13695 19078
rect 13997 19138 14063 19141
rect 21817 19138 21883 19141
rect 13997 19136 21883 19138
rect 13997 19080 14002 19136
rect 14058 19080 21822 19136
rect 21878 19080 21883 19136
rect 13997 19078 21883 19080
rect 13997 19075 14063 19078
rect 21817 19075 21883 19078
rect 28901 19136 29010 19141
rect 28901 19080 28906 19136
rect 28962 19080 29010 19136
rect 28901 19078 29010 19080
rect 28901 19075 28967 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 9949 19002 10015 19005
rect 21909 19002 21975 19005
rect 9949 19000 21975 19002
rect 9949 18944 9954 19000
rect 10010 18944 21914 19000
rect 21970 18944 21975 19000
rect 9949 18942 21975 18944
rect 9949 18939 10015 18942
rect 21909 18939 21975 18942
rect 23197 19002 23263 19005
rect 28533 19002 28599 19005
rect 23197 19000 28599 19002
rect 23197 18944 23202 19000
rect 23258 18944 28538 19000
rect 28594 18944 28599 19000
rect 23197 18942 28599 18944
rect 23197 18939 23263 18942
rect 28533 18939 28599 18942
rect 3141 18866 3207 18869
rect 24117 18866 24183 18869
rect 3141 18864 24183 18866
rect 3141 18808 3146 18864
rect 3202 18808 24122 18864
rect 24178 18808 24183 18864
rect 3141 18806 24183 18808
rect 3141 18803 3207 18806
rect 24117 18803 24183 18806
rect 25773 18866 25839 18869
rect 29269 18866 29335 18869
rect 25773 18864 29335 18866
rect 25773 18808 25778 18864
rect 25834 18808 29274 18864
rect 29330 18808 29335 18864
rect 25773 18806 29335 18808
rect 25773 18803 25839 18806
rect 29269 18803 29335 18806
rect 10593 18730 10659 18733
rect 10961 18730 11027 18733
rect 10593 18728 11027 18730
rect 10593 18672 10598 18728
rect 10654 18672 10966 18728
rect 11022 18672 11027 18728
rect 10593 18670 11027 18672
rect 10593 18667 10659 18670
rect 10961 18667 11027 18670
rect 12433 18730 12499 18733
rect 13077 18730 13143 18733
rect 12433 18728 13143 18730
rect 12433 18672 12438 18728
rect 12494 18672 13082 18728
rect 13138 18672 13143 18728
rect 12433 18670 13143 18672
rect 12433 18667 12499 18670
rect 13077 18667 13143 18670
rect 19885 18730 19951 18733
rect 22185 18730 22251 18733
rect 19885 18728 22251 18730
rect 19885 18672 19890 18728
rect 19946 18672 22190 18728
rect 22246 18672 22251 18728
rect 19885 18670 22251 18672
rect 19885 18667 19951 18670
rect 22185 18667 22251 18670
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 9857 18322 9923 18325
rect 23013 18322 23079 18325
rect 9857 18320 23079 18322
rect 9857 18264 9862 18320
rect 9918 18264 23018 18320
rect 23074 18264 23079 18320
rect 9857 18262 23079 18264
rect 9857 18259 9923 18262
rect 23013 18259 23079 18262
rect 10593 18186 10659 18189
rect 11329 18186 11395 18189
rect 10593 18184 11395 18186
rect 10593 18128 10598 18184
rect 10654 18128 11334 18184
rect 11390 18128 11395 18184
rect 10593 18126 11395 18128
rect 10593 18123 10659 18126
rect 11329 18123 11395 18126
rect 18965 18186 19031 18189
rect 19241 18186 19307 18189
rect 18965 18184 19307 18186
rect 18965 18128 18970 18184
rect 19026 18128 19246 18184
rect 19302 18128 19307 18184
rect 18965 18126 19307 18128
rect 18965 18123 19031 18126
rect 19241 18123 19307 18126
rect 19793 18186 19859 18189
rect 25313 18186 25379 18189
rect 19793 18184 25379 18186
rect 19793 18128 19798 18184
rect 19854 18128 25318 18184
rect 25374 18128 25379 18184
rect 19793 18126 25379 18128
rect 19793 18123 19859 18126
rect 25313 18123 25379 18126
rect 5533 18050 5599 18053
rect 9622 18050 9628 18052
rect 5533 18048 9628 18050
rect 5533 17992 5538 18048
rect 5594 17992 9628 18048
rect 5533 17990 9628 17992
rect 5533 17987 5599 17990
rect 9622 17988 9628 17990
rect 9692 17988 9698 18052
rect 10409 18050 10475 18053
rect 11697 18050 11763 18053
rect 12617 18050 12683 18053
rect 10409 18048 12683 18050
rect 10409 17992 10414 18048
rect 10470 17992 11702 18048
rect 11758 17992 12622 18048
rect 12678 17992 12683 18048
rect 10409 17990 12683 17992
rect 10409 17987 10475 17990
rect 11697 17987 11763 17990
rect 12617 17987 12683 17990
rect 14917 18050 14983 18053
rect 20478 18050 20484 18052
rect 14917 18048 20484 18050
rect 14917 17992 14922 18048
rect 14978 17992 20484 18048
rect 14917 17990 20484 17992
rect 14917 17987 14983 17990
rect 20478 17988 20484 17990
rect 20548 18050 20554 18052
rect 22829 18050 22895 18053
rect 20548 18048 22895 18050
rect 20548 17992 22834 18048
rect 22890 17992 22895 18048
rect 20548 17990 22895 17992
rect 20548 17988 20554 17990
rect 22829 17987 22895 17990
rect 28625 18050 28691 18053
rect 31017 18050 31083 18053
rect 28625 18048 31083 18050
rect 28625 17992 28630 18048
rect 28686 17992 31022 18048
rect 31078 17992 31083 18048
rect 28625 17990 31083 17992
rect 28625 17987 28691 17990
rect 31017 17987 31083 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 11237 17914 11303 17917
rect 15561 17914 15627 17917
rect 19333 17916 19399 17917
rect 19333 17914 19380 17916
rect 11237 17912 15627 17914
rect 11237 17856 11242 17912
rect 11298 17856 15566 17912
rect 15622 17856 15627 17912
rect 11237 17854 15627 17856
rect 19288 17912 19380 17914
rect 19288 17856 19338 17912
rect 19288 17854 19380 17856
rect 11237 17851 11303 17854
rect 15561 17851 15627 17854
rect 19333 17852 19380 17854
rect 19444 17852 19450 17916
rect 19701 17914 19767 17917
rect 21817 17914 21883 17917
rect 19701 17912 21883 17914
rect 19701 17856 19706 17912
rect 19762 17856 21822 17912
rect 21878 17856 21883 17912
rect 19701 17854 21883 17856
rect 19333 17851 19399 17852
rect 19701 17851 19767 17854
rect 21817 17851 21883 17854
rect 21950 17852 21956 17916
rect 22020 17914 22026 17916
rect 23105 17914 23171 17917
rect 22020 17912 23171 17914
rect 22020 17856 23110 17912
rect 23166 17856 23171 17912
rect 22020 17854 23171 17856
rect 22020 17852 22026 17854
rect 23105 17851 23171 17854
rect 7465 17778 7531 17781
rect 22921 17778 22987 17781
rect 7465 17776 22987 17778
rect 7465 17720 7470 17776
rect 7526 17720 22926 17776
rect 22982 17720 22987 17776
rect 7465 17718 22987 17720
rect 7465 17715 7531 17718
rect 22921 17715 22987 17718
rect 38377 17778 38443 17781
rect 38618 17778 39418 17808
rect 38377 17776 39418 17778
rect 38377 17720 38382 17776
rect 38438 17720 39418 17776
rect 38377 17718 39418 17720
rect 38377 17715 38443 17718
rect 38618 17688 39418 17718
rect 12065 17642 12131 17645
rect 27613 17642 27679 17645
rect 12065 17640 27679 17642
rect 12065 17584 12070 17640
rect 12126 17584 27618 17640
rect 27674 17584 27679 17640
rect 12065 17582 27679 17584
rect 12065 17579 12131 17582
rect 27613 17579 27679 17582
rect 8017 17506 8083 17509
rect 9581 17506 9647 17509
rect 8017 17504 9647 17506
rect 8017 17448 8022 17504
rect 8078 17448 9586 17504
rect 9642 17448 9647 17504
rect 8017 17446 9647 17448
rect 8017 17443 8083 17446
rect 9581 17443 9647 17446
rect 12801 17506 12867 17509
rect 18413 17506 18479 17509
rect 12801 17504 18479 17506
rect 12801 17448 12806 17504
rect 12862 17448 18418 17504
rect 18474 17448 18479 17504
rect 12801 17446 18479 17448
rect 12801 17443 12867 17446
rect 18413 17443 18479 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 13077 17370 13143 17373
rect 17769 17370 17835 17373
rect 13077 17368 17835 17370
rect 13077 17312 13082 17368
rect 13138 17312 17774 17368
rect 17830 17312 17835 17368
rect 13077 17310 17835 17312
rect 13077 17307 13143 17310
rect 17769 17307 17835 17310
rect 20294 17308 20300 17372
rect 20364 17370 20370 17372
rect 20437 17370 20503 17373
rect 20364 17368 20503 17370
rect 20364 17312 20442 17368
rect 20498 17312 20503 17368
rect 20364 17310 20503 17312
rect 20364 17308 20370 17310
rect 20437 17307 20503 17310
rect 23841 17370 23907 17373
rect 23974 17370 23980 17372
rect 23841 17368 23980 17370
rect 23841 17312 23846 17368
rect 23902 17312 23980 17368
rect 23841 17310 23980 17312
rect 23841 17307 23907 17310
rect 23974 17308 23980 17310
rect 24044 17308 24050 17372
rect 4429 17234 4495 17237
rect 6361 17234 6427 17237
rect 26417 17234 26483 17237
rect 4429 17232 26483 17234
rect 4429 17176 4434 17232
rect 4490 17176 6366 17232
rect 6422 17176 26422 17232
rect 26478 17176 26483 17232
rect 4429 17174 26483 17176
rect 4429 17171 4495 17174
rect 6361 17171 6427 17174
rect 26417 17171 26483 17174
rect 29177 17234 29243 17237
rect 35525 17234 35591 17237
rect 29177 17232 35591 17234
rect 29177 17176 29182 17232
rect 29238 17176 35530 17232
rect 35586 17176 35591 17232
rect 29177 17174 35591 17176
rect 29177 17171 29243 17174
rect 35525 17171 35591 17174
rect 19793 17098 19859 17101
rect 20110 17098 20116 17100
rect 19793 17096 20116 17098
rect 19793 17040 19798 17096
rect 19854 17040 20116 17096
rect 19793 17038 20116 17040
rect 19793 17035 19859 17038
rect 20110 17036 20116 17038
rect 20180 17036 20186 17100
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 13118 16764 13124 16828
rect 13188 16826 13194 16828
rect 13721 16826 13787 16829
rect 13188 16824 17050 16826
rect 13188 16768 13726 16824
rect 13782 16768 17050 16824
rect 13188 16766 17050 16768
rect 13188 16764 13194 16766
rect 13721 16763 13787 16766
rect 16990 16692 17050 16766
rect 16982 16628 16988 16692
rect 17052 16628 17058 16692
rect 5441 16554 5507 16557
rect 17953 16554 18019 16557
rect 20437 16554 20503 16557
rect 5441 16552 18019 16554
rect 5441 16496 5446 16552
rect 5502 16496 17958 16552
rect 18014 16496 18019 16552
rect 5441 16494 18019 16496
rect 5441 16491 5507 16494
rect 17953 16491 18019 16494
rect 18094 16552 20503 16554
rect 18094 16496 20442 16552
rect 20498 16496 20503 16552
rect 18094 16494 20503 16496
rect 9673 16420 9739 16421
rect 9622 16356 9628 16420
rect 9692 16418 9739 16420
rect 12893 16418 12959 16421
rect 18094 16418 18154 16494
rect 20437 16491 20503 16494
rect 21766 16492 21772 16556
rect 21836 16554 21842 16556
rect 21909 16554 21975 16557
rect 21836 16552 21975 16554
rect 21836 16496 21914 16552
rect 21970 16496 21975 16552
rect 21836 16494 21975 16496
rect 21836 16492 21842 16494
rect 21909 16491 21975 16494
rect 22921 16554 22987 16557
rect 24301 16556 24367 16557
rect 23606 16554 23612 16556
rect 22921 16552 23612 16554
rect 22921 16496 22926 16552
rect 22982 16496 23612 16552
rect 22921 16494 23612 16496
rect 22921 16491 22987 16494
rect 23606 16492 23612 16494
rect 23676 16492 23682 16556
rect 24301 16554 24348 16556
rect 24256 16552 24348 16554
rect 24256 16496 24306 16552
rect 24256 16494 24348 16496
rect 24301 16492 24348 16494
rect 24412 16492 24418 16556
rect 24301 16491 24367 16492
rect 9692 16416 9784 16418
rect 9734 16360 9784 16416
rect 9692 16358 9784 16360
rect 12893 16416 18154 16418
rect 12893 16360 12898 16416
rect 12954 16360 18154 16416
rect 12893 16358 18154 16360
rect 9692 16356 9739 16358
rect 9673 16355 9739 16356
rect 12893 16355 12959 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 16982 16084 16988 16148
rect 17052 16146 17058 16148
rect 25129 16146 25195 16149
rect 17052 16144 25195 16146
rect 17052 16088 25134 16144
rect 25190 16088 25195 16144
rect 17052 16086 25195 16088
rect 17052 16084 17058 16086
rect 25129 16083 25195 16086
rect 9029 16010 9095 16013
rect 37641 16010 37707 16013
rect 9029 16008 37707 16010
rect 9029 15952 9034 16008
rect 9090 15952 37646 16008
rect 37702 15952 37707 16008
rect 9029 15950 37707 15952
rect 9029 15947 9095 15950
rect 37641 15947 37707 15950
rect 15837 15874 15903 15877
rect 16849 15874 16915 15877
rect 15837 15872 16915 15874
rect 15837 15816 15842 15872
rect 15898 15816 16854 15872
rect 16910 15816 16915 15872
rect 15837 15814 16915 15816
rect 15837 15811 15903 15814
rect 16849 15811 16915 15814
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 13077 15738 13143 15741
rect 24301 15738 24367 15741
rect 13077 15736 24367 15738
rect 13077 15680 13082 15736
rect 13138 15680 24306 15736
rect 24362 15680 24367 15736
rect 13077 15678 24367 15680
rect 13077 15675 13143 15678
rect 24301 15675 24367 15678
rect 37825 15738 37891 15741
rect 38618 15738 39418 15768
rect 37825 15736 39418 15738
rect 37825 15680 37830 15736
rect 37886 15680 39418 15736
rect 37825 15678 39418 15680
rect 37825 15675 37891 15678
rect 38618 15648 39418 15678
rect 15837 15602 15903 15605
rect 17861 15602 17927 15605
rect 15837 15600 17927 15602
rect 15837 15544 15842 15600
rect 15898 15544 17866 15600
rect 17922 15544 17927 15600
rect 15837 15542 17927 15544
rect 15837 15539 15903 15542
rect 16254 15333 16314 15542
rect 17861 15539 17927 15542
rect 20345 15466 20411 15469
rect 21030 15466 21036 15468
rect 20345 15464 21036 15466
rect 20345 15408 20350 15464
rect 20406 15408 21036 15464
rect 20345 15406 21036 15408
rect 20345 15403 20411 15406
rect 21030 15404 21036 15406
rect 21100 15466 21106 15468
rect 23197 15466 23263 15469
rect 21100 15464 23263 15466
rect 21100 15408 23202 15464
rect 23258 15408 23263 15464
rect 21100 15406 23263 15408
rect 21100 15404 21106 15406
rect 23197 15403 23263 15406
rect 16254 15328 16363 15333
rect 16254 15272 16302 15328
rect 16358 15272 16363 15328
rect 16254 15270 16363 15272
rect 16297 15267 16363 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 9029 15196 9095 15197
rect 9029 15192 9076 15196
rect 9140 15194 9146 15196
rect 15837 15194 15903 15197
rect 18321 15194 18387 15197
rect 9029 15136 9034 15192
rect 9029 15132 9076 15136
rect 9140 15134 9186 15194
rect 15837 15192 18387 15194
rect 15837 15136 15842 15192
rect 15898 15136 18326 15192
rect 18382 15136 18387 15192
rect 15837 15134 18387 15136
rect 9140 15132 9146 15134
rect 9029 15131 9095 15132
rect 15837 15131 15903 15134
rect 18321 15131 18387 15134
rect 15745 15058 15811 15061
rect 17953 15058 18019 15061
rect 15745 15056 18019 15058
rect 15745 15000 15750 15056
rect 15806 15000 17958 15056
rect 18014 15000 18019 15056
rect 15745 14998 18019 15000
rect 15745 14995 15811 14998
rect 17953 14995 18019 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 27337 14514 27403 14517
rect 30741 14514 30807 14517
rect 27337 14512 30807 14514
rect 27337 14456 27342 14512
rect 27398 14456 30746 14512
rect 30802 14456 30807 14512
rect 27337 14454 30807 14456
rect 27337 14451 27403 14454
rect 30741 14451 30807 14454
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 16757 14106 16823 14109
rect 18781 14106 18847 14109
rect 16757 14104 18847 14106
rect 16757 14048 16762 14104
rect 16818 14048 18786 14104
rect 18842 14048 18847 14104
rect 16757 14046 18847 14048
rect 16757 14043 16823 14046
rect 18781 14043 18847 14046
rect 16430 13908 16436 13972
rect 16500 13970 16506 13972
rect 17861 13970 17927 13973
rect 16500 13968 17927 13970
rect 16500 13912 17866 13968
rect 17922 13912 17927 13968
rect 16500 13910 17927 13912
rect 16500 13908 16506 13910
rect 17861 13907 17927 13910
rect 24853 13834 24919 13837
rect 28533 13834 28599 13837
rect 24853 13832 28599 13834
rect 24853 13776 24858 13832
rect 24914 13776 28538 13832
rect 28594 13776 28599 13832
rect 24853 13774 28599 13776
rect 24853 13771 24919 13774
rect 28533 13771 28599 13774
rect 0 13698 800 13728
rect 933 13698 999 13701
rect 0 13696 999 13698
rect 0 13640 938 13696
rect 994 13640 999 13696
rect 0 13638 999 13640
rect 0 13608 800 13638
rect 933 13635 999 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 38618 13608 39418 13728
rect 34930 13567 35246 13568
rect 23657 13426 23723 13429
rect 25865 13426 25931 13429
rect 23657 13424 25931 13426
rect 23657 13368 23662 13424
rect 23718 13368 25870 13424
rect 25926 13368 25931 13424
rect 23657 13366 25931 13368
rect 23657 13363 23723 13366
rect 25865 13363 25931 13366
rect 23105 13290 23171 13293
rect 28441 13290 28507 13293
rect 23105 13288 28507 13290
rect 23105 13232 23110 13288
rect 23166 13232 28446 13288
rect 28502 13232 28507 13288
rect 23105 13230 28507 13232
rect 23105 13227 23171 13230
rect 28441 13227 28507 13230
rect 28993 13154 29059 13157
rect 29269 13154 29335 13157
rect 28993 13152 29335 13154
rect 28993 13096 28998 13152
rect 29054 13096 29274 13152
rect 29330 13096 29335 13152
rect 28993 13094 29335 13096
rect 28993 13091 29059 13094
rect 29269 13091 29335 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 28993 13018 29059 13021
rect 29361 13018 29427 13021
rect 28993 13016 29427 13018
rect 28993 12960 28998 13016
rect 29054 12960 29366 13016
rect 29422 12960 29427 13016
rect 28993 12958 29427 12960
rect 28993 12955 29059 12958
rect 29361 12955 29427 12958
rect 22093 12882 22159 12885
rect 25037 12882 25103 12885
rect 22093 12880 25103 12882
rect 22093 12824 22098 12880
rect 22154 12824 25042 12880
rect 25098 12824 25103 12880
rect 22093 12822 25103 12824
rect 22093 12819 22159 12822
rect 25037 12819 25103 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 26417 12474 26483 12477
rect 31293 12474 31359 12477
rect 26417 12472 31359 12474
rect 26417 12416 26422 12472
rect 26478 12416 31298 12472
rect 31354 12416 31359 12472
rect 26417 12414 31359 12416
rect 26417 12411 26483 12414
rect 31293 12411 31359 12414
rect 21173 12202 21239 12205
rect 26877 12202 26943 12205
rect 21173 12200 26943 12202
rect 21173 12144 21178 12200
rect 21234 12144 26882 12200
rect 26938 12144 26943 12200
rect 21173 12142 26943 12144
rect 21173 12139 21239 12142
rect 26877 12139 26943 12142
rect 22921 12066 22987 12069
rect 25957 12066 26023 12069
rect 22921 12064 26023 12066
rect 22921 12008 22926 12064
rect 22982 12008 25962 12064
rect 26018 12008 26023 12064
rect 22921 12006 26023 12008
rect 22921 12003 22987 12006
rect 25957 12003 26023 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 27245 11932 27311 11933
rect 27245 11930 27292 11932
rect 27200 11928 27292 11930
rect 27200 11872 27250 11928
rect 27200 11870 27292 11872
rect 27245 11868 27292 11870
rect 27356 11868 27362 11932
rect 27245 11867 27311 11868
rect 19609 11794 19675 11797
rect 20478 11794 20484 11796
rect 19609 11792 20484 11794
rect 19609 11736 19614 11792
rect 19670 11736 20484 11792
rect 19609 11734 20484 11736
rect 19609 11731 19675 11734
rect 20478 11732 20484 11734
rect 20548 11732 20554 11796
rect 24485 11794 24551 11797
rect 26509 11794 26575 11797
rect 24485 11792 26575 11794
rect 24485 11736 24490 11792
rect 24546 11736 26514 11792
rect 26570 11736 26575 11792
rect 24485 11734 26575 11736
rect 24485 11731 24551 11734
rect 26509 11731 26575 11734
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 19241 11658 19307 11661
rect 37273 11658 37339 11661
rect 19241 11656 37339 11658
rect 19241 11600 19246 11656
rect 19302 11600 37278 11656
rect 37334 11600 37339 11656
rect 19241 11598 37339 11600
rect 19241 11595 19307 11598
rect 37273 11595 37339 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 13261 11114 13327 11117
rect 25589 11114 25655 11117
rect 13261 11112 25655 11114
rect 13261 11056 13266 11112
rect 13322 11056 25594 11112
rect 25650 11056 25655 11112
rect 13261 11054 25655 11056
rect 13261 11051 13327 11054
rect 25589 11051 25655 11054
rect 28073 11114 28139 11117
rect 29678 11114 29684 11116
rect 28073 11112 29684 11114
rect 28073 11056 28078 11112
rect 28134 11056 29684 11112
rect 28073 11054 29684 11056
rect 28073 11051 28139 11054
rect 29678 11052 29684 11054
rect 29748 11052 29754 11116
rect 18454 10916 18460 10980
rect 18524 10978 18530 10980
rect 18597 10978 18663 10981
rect 18524 10976 18663 10978
rect 18524 10920 18602 10976
rect 18658 10920 18663 10976
rect 18524 10918 18663 10920
rect 18524 10916 18530 10918
rect 18597 10915 18663 10918
rect 37917 10978 37983 10981
rect 38618 10978 39418 11008
rect 37917 10976 39418 10978
rect 37917 10920 37922 10976
rect 37978 10920 39418 10976
rect 37917 10918 39418 10920
rect 37917 10915 37983 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 38618 10888 39418 10918
rect 19570 10847 19886 10848
rect 10133 10706 10199 10709
rect 10358 10706 10364 10708
rect 10133 10704 10364 10706
rect 10133 10648 10138 10704
rect 10194 10648 10364 10704
rect 10133 10646 10364 10648
rect 10133 10643 10199 10646
rect 10358 10644 10364 10646
rect 10428 10644 10434 10708
rect 10317 10434 10383 10437
rect 21449 10434 21515 10437
rect 22185 10434 22251 10437
rect 10317 10432 22251 10434
rect 10317 10376 10322 10432
rect 10378 10376 21454 10432
rect 21510 10376 22190 10432
rect 22246 10376 22251 10432
rect 10317 10374 22251 10376
rect 10317 10371 10383 10374
rect 21449 10371 21515 10374
rect 22185 10371 22251 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 21081 10162 21147 10165
rect 21909 10162 21975 10165
rect 21081 10160 21975 10162
rect 21081 10104 21086 10160
rect 21142 10104 21914 10160
rect 21970 10104 21975 10160
rect 21081 10102 21975 10104
rect 21081 10099 21147 10102
rect 21909 10099 21975 10102
rect 19885 10026 19951 10029
rect 21081 10026 21147 10029
rect 19885 10024 21147 10026
rect 19885 9968 19890 10024
rect 19946 9968 21086 10024
rect 21142 9968 21147 10024
rect 19885 9966 21147 9968
rect 19885 9963 19951 9966
rect 21081 9963 21147 9966
rect 22461 10026 22527 10029
rect 23657 10026 23723 10029
rect 24393 10026 24459 10029
rect 22461 10024 24459 10026
rect 22461 9968 22466 10024
rect 22522 9968 23662 10024
rect 23718 9968 24398 10024
rect 24454 9968 24459 10024
rect 22461 9966 24459 9968
rect 22461 9963 22527 9966
rect 23657 9963 23723 9966
rect 24393 9963 24459 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 15009 9754 15075 9757
rect 18137 9754 18203 9757
rect 15009 9752 18203 9754
rect 15009 9696 15014 9752
rect 15070 9696 18142 9752
rect 18198 9696 18203 9752
rect 15009 9694 18203 9696
rect 15009 9691 15075 9694
rect 18137 9691 18203 9694
rect 3233 9618 3299 9621
rect 5441 9618 5507 9621
rect 3233 9616 5507 9618
rect 3233 9560 3238 9616
rect 3294 9560 5446 9616
rect 5502 9560 5507 9616
rect 3233 9558 5507 9560
rect 3233 9555 3299 9558
rect 5441 9555 5507 9558
rect 8201 9618 8267 9621
rect 8937 9618 9003 9621
rect 8201 9616 9003 9618
rect 8201 9560 8206 9616
rect 8262 9560 8942 9616
rect 8998 9560 9003 9616
rect 8201 9558 9003 9560
rect 8201 9555 8267 9558
rect 8937 9555 9003 9558
rect 17861 9618 17927 9621
rect 20294 9618 20300 9620
rect 17861 9616 20300 9618
rect 17861 9560 17866 9616
rect 17922 9560 20300 9616
rect 17861 9558 20300 9560
rect 17861 9555 17927 9558
rect 20294 9556 20300 9558
rect 20364 9556 20370 9620
rect 23841 9618 23907 9621
rect 25865 9618 25931 9621
rect 23841 9616 25931 9618
rect 23841 9560 23846 9616
rect 23902 9560 25870 9616
rect 25926 9560 25931 9616
rect 23841 9558 25931 9560
rect 23841 9555 23907 9558
rect 25865 9555 25931 9558
rect 29678 9556 29684 9620
rect 29748 9618 29754 9620
rect 31201 9618 31267 9621
rect 29748 9616 31267 9618
rect 29748 9560 31206 9616
rect 31262 9560 31267 9616
rect 29748 9558 31267 9560
rect 29748 9556 29754 9558
rect 31201 9555 31267 9558
rect 19793 9482 19859 9485
rect 24485 9482 24551 9485
rect 19793 9480 24551 9482
rect 19793 9424 19798 9480
rect 19854 9424 24490 9480
rect 24546 9424 24551 9480
rect 19793 9422 24551 9424
rect 19793 9419 19859 9422
rect 24485 9419 24551 9422
rect 25589 9482 25655 9485
rect 25957 9482 26023 9485
rect 25589 9480 26023 9482
rect 25589 9424 25594 9480
rect 25650 9424 25962 9480
rect 26018 9424 26023 9480
rect 25589 9422 26023 9424
rect 25589 9419 25655 9422
rect 25957 9419 26023 9422
rect 29545 9482 29611 9485
rect 36629 9482 36695 9485
rect 29545 9480 36695 9482
rect 29545 9424 29550 9480
rect 29606 9424 36634 9480
rect 36690 9424 36695 9480
rect 29545 9422 36695 9424
rect 29545 9419 29611 9422
rect 36629 9419 36695 9422
rect 22461 9346 22527 9349
rect 25037 9346 25103 9349
rect 22461 9344 25103 9346
rect 22461 9288 22466 9344
rect 22522 9288 25042 9344
rect 25098 9288 25103 9344
rect 22461 9286 25103 9288
rect 22461 9283 22527 9286
rect 25037 9283 25103 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 38101 8938 38167 8941
rect 38618 8938 39418 8968
rect 38101 8936 39418 8938
rect 38101 8880 38106 8936
rect 38162 8880 39418 8936
rect 38101 8878 39418 8880
rect 38101 8875 38167 8878
rect 38618 8848 39418 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 19977 8666 20043 8669
rect 20662 8666 20668 8668
rect 19977 8664 20668 8666
rect 19977 8608 19982 8664
rect 20038 8608 20668 8664
rect 19977 8606 20668 8608
rect 19977 8603 20043 8606
rect 20662 8604 20668 8606
rect 20732 8604 20738 8668
rect 4061 8530 4127 8533
rect 23974 8530 23980 8532
rect 4061 8528 23980 8530
rect 4061 8472 4066 8528
rect 4122 8472 23980 8528
rect 4061 8470 23980 8472
rect 4061 8467 4127 8470
rect 23974 8468 23980 8470
rect 24044 8530 24050 8532
rect 24301 8530 24367 8533
rect 24044 8528 24367 8530
rect 24044 8472 24306 8528
rect 24362 8472 24367 8528
rect 24044 8470 24367 8472
rect 24044 8468 24050 8470
rect 24301 8467 24367 8470
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 18689 6900 18755 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 18638 6836 18644 6900
rect 18708 6898 18755 6900
rect 18708 6896 18800 6898
rect 18750 6840 18800 6896
rect 18708 6838 18800 6840
rect 18708 6836 18755 6838
rect 18689 6835 18755 6836
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 38618 6128 39418 6248
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 25313 4178 25379 4181
rect 28073 4178 28139 4181
rect 25313 4176 28139 4178
rect 25313 4120 25318 4176
rect 25374 4120 28078 4176
rect 28134 4120 28139 4176
rect 25313 4118 28139 4120
rect 25313 4115 25379 4118
rect 28073 4115 28139 4118
rect 38618 4088 39418 4208
rect 11789 4044 11855 4045
rect 11789 4040 11836 4044
rect 11900 4042 11906 4044
rect 13169 4042 13235 4045
rect 13302 4042 13308 4044
rect 11789 3984 11794 4040
rect 11789 3980 11836 3984
rect 11900 3982 11946 4042
rect 13169 4040 13308 4042
rect 13169 3984 13174 4040
rect 13230 3984 13308 4040
rect 13169 3982 13308 3984
rect 11900 3980 11906 3982
rect 11789 3979 11855 3980
rect 13169 3979 13235 3982
rect 13302 3980 13308 3982
rect 13372 3980 13378 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 0 2048 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 37181 1458 37247 1461
rect 38618 1458 39418 1488
rect 37181 1456 39418 1458
rect 37181 1400 37186 1456
rect 37242 1400 39418 1456
rect 37181 1398 39418 1400
rect 37181 1395 37247 1398
rect 38618 1368 39418 1398
<< via3 >>
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 12204 38660 12268 38724
rect 23428 38660 23492 38724
rect 23980 38660 24044 38724
rect 27476 38660 27540 38724
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 14228 37300 14292 37364
rect 13492 37164 13556 37228
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 22324 36756 22388 36820
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 13124 35940 13188 36004
rect 23060 35940 23124 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 22324 35396 22388 35460
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 24348 34716 24412 34780
rect 25636 34716 25700 34780
rect 25452 34444 25516 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 20668 33220 20732 33284
rect 21956 33220 22020 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 23060 33144 23124 33148
rect 23060 33088 23110 33144
rect 23110 33088 23124 33144
rect 23060 33084 23124 33088
rect 22508 32676 22572 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 21588 32540 21652 32604
rect 20484 32404 20548 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 18644 31996 18708 32060
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 27108 31920 27172 31924
rect 27108 31864 27158 31920
rect 27158 31864 27172 31920
rect 27108 31860 27172 31864
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 19380 31452 19444 31516
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19380 30908 19444 30972
rect 19012 30772 19076 30836
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 23612 30364 23676 30428
rect 27292 30364 27356 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 21588 29820 21652 29884
rect 20116 29548 20180 29612
rect 22140 29608 22204 29612
rect 22140 29552 22154 29608
rect 22154 29552 22204 29608
rect 22140 29548 22204 29552
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 13308 29064 13372 29068
rect 13308 29008 13358 29064
rect 13358 29008 13372 29064
rect 13308 29004 13372 29008
rect 18460 29004 18524 29068
rect 19012 29004 19076 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 22508 28596 22572 28660
rect 20300 28460 20364 28524
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 23060 28052 23124 28116
rect 21772 27780 21836 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 21036 27704 21100 27708
rect 21036 27648 21050 27704
rect 21050 27648 21100 27704
rect 21036 27644 21100 27648
rect 14228 27296 14292 27300
rect 14228 27240 14242 27296
rect 14242 27240 14292 27296
rect 14228 27236 14292 27240
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 22140 26420 22204 26484
rect 19380 26148 19444 26212
rect 25452 26148 25516 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 11836 25196 11900 25260
rect 20300 25120 20364 25124
rect 20300 25064 20314 25120
rect 20314 25064 20364 25120
rect 20300 25060 20364 25064
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 27108 24848 27172 24852
rect 27108 24792 27122 24848
rect 27122 24792 27172 24848
rect 27108 24788 27172 24792
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 27476 23564 27540 23628
rect 16436 23488 16500 23492
rect 16436 23432 16486 23488
rect 16486 23432 16500 23488
rect 16436 23428 16500 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 23980 22476 24044 22540
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 12204 21992 12268 21996
rect 12204 21936 12254 21992
rect 12254 21936 12268 21992
rect 12204 21932 12268 21936
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 13492 21660 13556 21724
rect 23428 21660 23492 21724
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 9076 20768 9140 20772
rect 9076 20712 9090 20768
rect 9090 20712 9140 20768
rect 9076 20708 9140 20712
rect 10364 20768 10428 20772
rect 10364 20712 10378 20768
rect 10378 20712 10428 20768
rect 10364 20708 10428 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 25636 20632 25700 20636
rect 25636 20576 25650 20632
rect 25650 20576 25700 20632
rect 25636 20572 25700 20576
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 20484 19892 20548 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 9628 17988 9692 18052
rect 20484 17988 20548 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19380 17912 19444 17916
rect 19380 17856 19394 17912
rect 19394 17856 19444 17912
rect 19380 17852 19444 17856
rect 21956 17852 22020 17916
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 20300 17308 20364 17372
rect 23980 17308 24044 17372
rect 20116 17036 20180 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 13124 16764 13188 16828
rect 16988 16628 17052 16692
rect 9628 16416 9692 16420
rect 21772 16492 21836 16556
rect 23612 16492 23676 16556
rect 24348 16552 24412 16556
rect 24348 16496 24362 16552
rect 24362 16496 24412 16552
rect 24348 16492 24412 16496
rect 9628 16360 9678 16416
rect 9678 16360 9692 16416
rect 9628 16356 9692 16360
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 16988 16084 17052 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 21036 15404 21100 15468
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 9076 15192 9140 15196
rect 9076 15136 9090 15192
rect 9090 15136 9140 15192
rect 9076 15132 9140 15136
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 16436 13908 16500 13972
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 27292 11928 27356 11932
rect 27292 11872 27306 11928
rect 27306 11872 27356 11928
rect 27292 11868 27356 11872
rect 20484 11732 20548 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 29684 11052 29748 11116
rect 18460 10916 18524 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 10364 10644 10428 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 20300 9556 20364 9620
rect 29684 9556 29748 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 20668 8604 20732 8668
rect 23980 8468 24044 8532
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 18644 6896 18708 6900
rect 18644 6840 18694 6896
rect 18694 6840 18708 6896
rect 18644 6836 18708 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 11836 4040 11900 4044
rect 11836 3984 11850 4040
rect 11850 3984 11900 4040
rect 11836 3980 11900 3984
rect 13308 3980 13372 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 38656 4528 39216
rect 19568 39200 19888 39216
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 12203 38724 12269 38725
rect 12203 38660 12204 38724
rect 12268 38660 12269 38724
rect 12203 38659 12269 38660
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 11835 25260 11901 25261
rect 11835 25196 11836 25260
rect 11900 25196 11901 25260
rect 11835 25195 11901 25196
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 9075 20772 9141 20773
rect 9075 20708 9076 20772
rect 9140 20708 9141 20772
rect 9075 20707 9141 20708
rect 10363 20772 10429 20773
rect 10363 20708 10364 20772
rect 10428 20708 10429 20772
rect 10363 20707 10429 20708
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 9078 15197 9138 20707
rect 9627 18052 9693 18053
rect 9627 17988 9628 18052
rect 9692 17988 9693 18052
rect 9627 17987 9693 17988
rect 9630 16421 9690 17987
rect 9627 16420 9693 16421
rect 9627 16356 9628 16420
rect 9692 16356 9693 16420
rect 9627 16355 9693 16356
rect 9075 15196 9141 15197
rect 9075 15132 9076 15196
rect 9140 15132 9141 15196
rect 9075 15131 9141 15132
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 10366 10709 10426 20707
rect 10363 10708 10429 10709
rect 10363 10644 10364 10708
rect 10428 10644 10429 10708
rect 10363 10643 10429 10644
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 11838 4045 11898 25195
rect 12206 21997 12266 38659
rect 19568 38112 19888 39136
rect 23427 38724 23493 38725
rect 23427 38660 23428 38724
rect 23492 38660 23493 38724
rect 23427 38659 23493 38660
rect 23979 38724 24045 38725
rect 23979 38660 23980 38724
rect 24044 38660 24045 38724
rect 23979 38659 24045 38660
rect 27475 38724 27541 38725
rect 27475 38660 27476 38724
rect 27540 38660 27541 38724
rect 27475 38659 27541 38660
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 14227 37364 14293 37365
rect 14227 37300 14228 37364
rect 14292 37300 14293 37364
rect 14227 37299 14293 37300
rect 13491 37228 13557 37229
rect 13491 37164 13492 37228
rect 13556 37164 13557 37228
rect 13491 37163 13557 37164
rect 13123 36004 13189 36005
rect 13123 35940 13124 36004
rect 13188 35940 13189 36004
rect 13123 35939 13189 35940
rect 12203 21996 12269 21997
rect 12203 21932 12204 21996
rect 12268 21932 12269 21996
rect 12203 21931 12269 21932
rect 13126 16829 13186 35939
rect 13307 29068 13373 29069
rect 13307 29004 13308 29068
rect 13372 29004 13373 29068
rect 13307 29003 13373 29004
rect 13123 16828 13189 16829
rect 13123 16764 13124 16828
rect 13188 16764 13189 16828
rect 13123 16763 13189 16764
rect 13310 4045 13370 29003
rect 13494 21725 13554 37163
rect 14230 27301 14290 37299
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 22323 36820 22389 36821
rect 22323 36756 22324 36820
rect 22388 36756 22389 36820
rect 22323 36755 22389 36756
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 22326 35461 22386 36755
rect 23059 36004 23125 36005
rect 23059 35940 23060 36004
rect 23124 35940 23125 36004
rect 23059 35939 23125 35940
rect 22323 35460 22389 35461
rect 22323 35396 22324 35460
rect 22388 35396 22389 35460
rect 22323 35395 22389 35396
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 20667 33284 20733 33285
rect 20667 33220 20668 33284
rect 20732 33220 20733 33284
rect 20667 33219 20733 33220
rect 21955 33284 22021 33285
rect 21955 33220 21956 33284
rect 22020 33220 22021 33284
rect 21955 33219 22021 33220
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 18643 32060 18709 32061
rect 18643 31996 18644 32060
rect 18708 31996 18709 32060
rect 18643 31995 18709 31996
rect 18459 29068 18525 29069
rect 18459 29004 18460 29068
rect 18524 29004 18525 29068
rect 18459 29003 18525 29004
rect 14227 27300 14293 27301
rect 14227 27236 14228 27300
rect 14292 27236 14293 27300
rect 14227 27235 14293 27236
rect 16435 23492 16501 23493
rect 16435 23428 16436 23492
rect 16500 23428 16501 23492
rect 16435 23427 16501 23428
rect 13491 21724 13557 21725
rect 13491 21660 13492 21724
rect 13556 21660 13557 21724
rect 13491 21659 13557 21660
rect 16438 13973 16498 23427
rect 16987 16692 17053 16693
rect 16987 16628 16988 16692
rect 17052 16628 17053 16692
rect 16987 16627 17053 16628
rect 16990 16149 17050 16627
rect 16987 16148 17053 16149
rect 16987 16084 16988 16148
rect 17052 16084 17053 16148
rect 16987 16083 17053 16084
rect 16435 13972 16501 13973
rect 16435 13908 16436 13972
rect 16500 13908 16501 13972
rect 16435 13907 16501 13908
rect 18462 10981 18522 29003
rect 18459 10980 18525 10981
rect 18459 10916 18460 10980
rect 18524 10916 18525 10980
rect 18459 10915 18525 10916
rect 18646 6901 18706 31995
rect 19568 31584 19888 32608
rect 20483 32468 20549 32469
rect 20483 32404 20484 32468
rect 20548 32404 20549 32468
rect 20483 32403 20549 32404
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19379 31516 19445 31517
rect 19379 31452 19380 31516
rect 19444 31452 19445 31516
rect 19379 31451 19445 31452
rect 19382 30973 19442 31451
rect 19379 30972 19445 30973
rect 19379 30908 19380 30972
rect 19444 30908 19445 30972
rect 19379 30907 19445 30908
rect 19011 30836 19077 30837
rect 19011 30772 19012 30836
rect 19076 30772 19077 30836
rect 19011 30771 19077 30772
rect 19014 29069 19074 30771
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 20115 29612 20181 29613
rect 20115 29548 20116 29612
rect 20180 29548 20181 29612
rect 20115 29547 20181 29548
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19011 29068 19077 29069
rect 19011 29004 19012 29068
rect 19076 29004 19077 29068
rect 19011 29003 19077 29004
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19379 26212 19445 26213
rect 19379 26148 19380 26212
rect 19444 26148 19445 26212
rect 19379 26147 19445 26148
rect 19382 17917 19442 26147
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19379 17916 19445 17917
rect 19379 17852 19380 17916
rect 19444 17852 19445 17916
rect 19379 17851 19445 17852
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 20118 17101 20178 29547
rect 20299 28524 20365 28525
rect 20299 28460 20300 28524
rect 20364 28460 20365 28524
rect 20299 28459 20365 28460
rect 20302 25125 20362 28459
rect 20299 25124 20365 25125
rect 20299 25060 20300 25124
rect 20364 25060 20365 25124
rect 20299 25059 20365 25060
rect 20486 19957 20546 32403
rect 20483 19956 20549 19957
rect 20483 19892 20484 19956
rect 20548 19892 20549 19956
rect 20483 19891 20549 19892
rect 20483 18052 20549 18053
rect 20483 17988 20484 18052
rect 20548 17988 20549 18052
rect 20483 17987 20549 17988
rect 20299 17372 20365 17373
rect 20299 17308 20300 17372
rect 20364 17308 20365 17372
rect 20299 17307 20365 17308
rect 20115 17100 20181 17101
rect 20115 17036 20116 17100
rect 20180 17036 20181 17100
rect 20115 17035 20181 17036
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 20302 9621 20362 17307
rect 20486 11797 20546 17987
rect 20483 11796 20549 11797
rect 20483 11732 20484 11796
rect 20548 11732 20549 11796
rect 20483 11731 20549 11732
rect 20299 9620 20365 9621
rect 20299 9556 20300 9620
rect 20364 9556 20365 9620
rect 20299 9555 20365 9556
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 20670 8669 20730 33219
rect 21587 32604 21653 32605
rect 21587 32540 21588 32604
rect 21652 32540 21653 32604
rect 21587 32539 21653 32540
rect 21590 29885 21650 32539
rect 21587 29884 21653 29885
rect 21587 29820 21588 29884
rect 21652 29820 21653 29884
rect 21587 29819 21653 29820
rect 21771 27844 21837 27845
rect 21771 27780 21772 27844
rect 21836 27780 21837 27844
rect 21771 27779 21837 27780
rect 21035 27708 21101 27709
rect 21035 27644 21036 27708
rect 21100 27644 21101 27708
rect 21035 27643 21101 27644
rect 21038 15469 21098 27643
rect 21774 16557 21834 27779
rect 21958 17917 22018 33219
rect 23062 33149 23122 35939
rect 23059 33148 23125 33149
rect 23059 33084 23060 33148
rect 23124 33084 23125 33148
rect 23059 33083 23125 33084
rect 22507 32740 22573 32741
rect 22507 32676 22508 32740
rect 22572 32676 22573 32740
rect 22507 32675 22573 32676
rect 22139 29612 22205 29613
rect 22139 29548 22140 29612
rect 22204 29548 22205 29612
rect 22139 29547 22205 29548
rect 22142 26485 22202 29547
rect 22510 28661 22570 32675
rect 22507 28660 22573 28661
rect 22507 28596 22508 28660
rect 22572 28596 22573 28660
rect 22507 28595 22573 28596
rect 23062 28117 23122 33083
rect 23059 28116 23125 28117
rect 23059 28052 23060 28116
rect 23124 28052 23125 28116
rect 23059 28051 23125 28052
rect 22139 26484 22205 26485
rect 22139 26420 22140 26484
rect 22204 26420 22205 26484
rect 22139 26419 22205 26420
rect 23430 21725 23490 38659
rect 23611 30428 23677 30429
rect 23611 30364 23612 30428
rect 23676 30364 23677 30428
rect 23611 30363 23677 30364
rect 23427 21724 23493 21725
rect 23427 21660 23428 21724
rect 23492 21660 23493 21724
rect 23427 21659 23493 21660
rect 21955 17916 22021 17917
rect 21955 17852 21956 17916
rect 22020 17852 22021 17916
rect 21955 17851 22021 17852
rect 23614 16557 23674 30363
rect 23982 22541 24042 38659
rect 24347 34780 24413 34781
rect 24347 34716 24348 34780
rect 24412 34716 24413 34780
rect 24347 34715 24413 34716
rect 25635 34780 25701 34781
rect 25635 34716 25636 34780
rect 25700 34716 25701 34780
rect 25635 34715 25701 34716
rect 23979 22540 24045 22541
rect 23979 22476 23980 22540
rect 24044 22476 24045 22540
rect 23979 22475 24045 22476
rect 23979 17372 24045 17373
rect 23979 17308 23980 17372
rect 24044 17308 24045 17372
rect 23979 17307 24045 17308
rect 21771 16556 21837 16557
rect 21771 16492 21772 16556
rect 21836 16492 21837 16556
rect 21771 16491 21837 16492
rect 23611 16556 23677 16557
rect 23611 16492 23612 16556
rect 23676 16492 23677 16556
rect 23611 16491 23677 16492
rect 21035 15468 21101 15469
rect 21035 15404 21036 15468
rect 21100 15404 21101 15468
rect 21035 15403 21101 15404
rect 20667 8668 20733 8669
rect 20667 8604 20668 8668
rect 20732 8604 20733 8668
rect 20667 8603 20733 8604
rect 23982 8533 24042 17307
rect 24350 16557 24410 34715
rect 25451 34508 25517 34509
rect 25451 34444 25452 34508
rect 25516 34444 25517 34508
rect 25451 34443 25517 34444
rect 25454 26213 25514 34443
rect 25451 26212 25517 26213
rect 25451 26148 25452 26212
rect 25516 26148 25517 26212
rect 25451 26147 25517 26148
rect 25638 20637 25698 34715
rect 27107 31924 27173 31925
rect 27107 31860 27108 31924
rect 27172 31860 27173 31924
rect 27107 31859 27173 31860
rect 27110 24853 27170 31859
rect 27291 30428 27357 30429
rect 27291 30364 27292 30428
rect 27356 30364 27357 30428
rect 27291 30363 27357 30364
rect 27107 24852 27173 24853
rect 27107 24788 27108 24852
rect 27172 24788 27173 24852
rect 27107 24787 27173 24788
rect 25635 20636 25701 20637
rect 25635 20572 25636 20636
rect 25700 20572 25701 20636
rect 25635 20571 25701 20572
rect 24347 16556 24413 16557
rect 24347 16492 24348 16556
rect 24412 16492 24413 16556
rect 24347 16491 24413 16492
rect 27294 11933 27354 30363
rect 27478 23629 27538 38659
rect 34928 38656 35248 39216
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 27475 23628 27541 23629
rect 27475 23564 27476 23628
rect 27540 23564 27541 23628
rect 27475 23563 27541 23564
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 27291 11932 27357 11933
rect 27291 11868 27292 11932
rect 27356 11868 27357 11932
rect 27291 11867 27357 11868
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 29683 11116 29749 11117
rect 29683 11052 29684 11116
rect 29748 11052 29749 11116
rect 29683 11051 29749 11052
rect 29686 9621 29746 11051
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 29683 9620 29749 9621
rect 29683 9556 29684 9620
rect 29748 9556 29749 9620
rect 29683 9555 29749 9556
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 23979 8532 24045 8533
rect 23979 8468 23980 8532
rect 24044 8468 24045 8532
rect 23979 8467 24045 8468
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 18643 6900 18709 6901
rect 18643 6836 18644 6900
rect 18708 6836 18709 6900
rect 18643 6835 18709 6836
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 11835 4044 11901 4045
rect 11835 3980 11836 4044
rect 11900 3980 11901 4044
rect 11835 3979 11901 3980
rect 13307 4044 13373 4045
rect 13307 3980 13308 4044
rect 13372 3980 13373 4044
rect 13307 3979 13373 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _1275_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1276_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1688980957
transform 1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1278_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1279_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1280_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1281_
timestamp 1688980957
transform 1 0 18492 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _1282_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1283_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1285_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _1286_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14444 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  _1287_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_2  _1288_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20424 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _1289_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__a21boi_1  _1290_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1688980957
transform 1 0 17204 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__nand3b_2  _1293_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1294_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _1296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1297_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1298_
timestamp 1688980957
transform 1 0 19412 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_4  _1299_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_1  _1300_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_4  _1301_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  _1302_
timestamp 1688980957
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__a221oi_2  _1303_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1305_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1307_
timestamp 1688980957
transform 1 0 21068 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1308_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1309_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23736 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1311_
timestamp 1688980957
transform 1 0 15456 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _1312_
timestamp 1688980957
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 1688980957
transform 1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1314_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1315_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1316_
timestamp 1688980957
transform 1 0 11592 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1317_
timestamp 1688980957
transform 1 0 16560 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1318_
timestamp 1688980957
transform 1 0 15640 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1319_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1320_
timestamp 1688980957
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _1321_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_1  _1322_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1323_
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1324_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _1325_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1326_
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1688980957
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1328_
timestamp 1688980957
transform 1 0 16100 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1329_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1330_
timestamp 1688980957
transform 1 0 16928 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1331_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_8  _1332_
timestamp 1688980957
transform 1 0 17940 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _1333_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1334_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_8  _1335_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__or3_4  _1336_
timestamp 1688980957
transform 1 0 18032 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1337_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_4  _1338_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18676 0 -1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_1  _1339_
timestamp 1688980957
transform 1 0 13892 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1340_
timestamp 1688980957
transform 1 0 14260 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__o2bb2a_2  _1341_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1342_
timestamp 1688980957
transform 1 0 17940 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1343_
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1344_
timestamp 1688980957
transform 1 0 18584 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__a221o_1  _1345_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26312 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1346_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27140 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1347_
timestamp 1688980957
transform 1 0 27600 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1688980957
transform 1 0 28980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1349_
timestamp 1688980957
transform 1 0 17388 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1350_
timestamp 1688980957
transform 1 0 18400 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_2  _1351_
timestamp 1688980957
transform 1 0 16008 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 1688980957
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1353_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _1355_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_4  _1356_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1357_
timestamp 1688980957
transform 1 0 18124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1359_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16100 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1360_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_8  _1361_
timestamp 1688980957
transform 1 0 19136 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _1362_
timestamp 1688980957
transform 1 0 16928 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__o22ai_4  _1363_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _1364_
timestamp 1688980957
transform 1 0 16468 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_4  _1365_
timestamp 1688980957
transform 1 0 16192 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _1366_
timestamp 1688980957
transform 1 0 18584 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1367_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25576 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1368_
timestamp 1688980957
transform 1 0 19964 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__a211o_1  _1369_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24932 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1370_
timestamp 1688980957
transform 1 0 24656 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1371_
timestamp 1688980957
transform 1 0 25116 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1372_
timestamp 1688980957
transform 1 0 28980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1373_
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1374_
timestamp 1688980957
transform 1 0 28704 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1375_
timestamp 1688980957
transform 1 0 29256 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1376_
timestamp 1688980957
transform 1 0 29716 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1377_
timestamp 1688980957
transform 1 0 31004 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1378_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30452 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 1688980957
transform 1 0 25300 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1380_
timestamp 1688980957
transform 1 0 25300 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1381_
timestamp 1688980957
transform 1 0 25024 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1382_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1688980957
transform 1 0 28612 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1385_
timestamp 1688980957
transform 1 0 29900 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1386_
timestamp 1688980957
transform 1 0 30544 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1387_
timestamp 1688980957
transform 1 0 25576 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1388_
timestamp 1688980957
transform 1 0 25760 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1389_
timestamp 1688980957
transform 1 0 26312 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1390_
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1391_
timestamp 1688980957
transform 1 0 36248 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1688980957
transform 1 0 35512 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1393_
timestamp 1688980957
transform 1 0 35512 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1394_
timestamp 1688980957
transform 1 0 35512 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1395_
timestamp 1688980957
transform 1 0 29072 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1396_
timestamp 1688980957
transform 1 0 29808 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29624 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1398_
timestamp 1688980957
transform 1 0 24380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1399_
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp 1688980957
transform 1 0 25208 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1401_
timestamp 1688980957
transform 1 0 24564 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1402_
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1403_
timestamp 1688980957
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1404_
timestamp 1688980957
transform 1 0 25760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1405_
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1406_
timestamp 1688980957
transform 1 0 29992 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1688980957
transform 1 0 25484 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1408_
timestamp 1688980957
transform 1 0 26036 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1409_
timestamp 1688980957
transform 1 0 25300 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1410_
timestamp 1688980957
transform 1 0 26128 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1411_
timestamp 1688980957
transform 1 0 31004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp 1688980957
transform 1 0 31280 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1413_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1414_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1415_
timestamp 1688980957
transform 1 0 20148 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1416_
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1417_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20516 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_4  _1419_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_2  _1420_
timestamp 1688980957
transform 1 0 23000 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1421_
timestamp 1688980957
transform 1 0 22724 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1422_
timestamp 1688980957
transform 1 0 22264 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1423_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1424_
timestamp 1688980957
transform 1 0 21988 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1425_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1426_
timestamp 1688980957
transform 1 0 22908 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1427_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_4  _1428_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22264 0 1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__nor4_1  _1429_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21896 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1430_
timestamp 1688980957
transform 1 0 22172 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1431_
timestamp 1688980957
transform 1 0 21344 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _1432_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22816 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1433_
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1688980957
transform 1 0 12328 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1435_
timestamp 1688980957
transform 1 0 13156 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1437_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__o211ai_4  _1438_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1439_
timestamp 1688980957
transform 1 0 25392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1440_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1441_
timestamp 1688980957
transform 1 0 18032 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _1442_
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1443_
timestamp 1688980957
transform 1 0 16744 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1444_
timestamp 1688980957
transform 1 0 23644 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1445_
timestamp 1688980957
transform 1 0 17480 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1446_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16468 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1688980957
transform 1 0 22172 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1448_
timestamp 1688980957
transform 1 0 22632 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1449_
timestamp 1688980957
transform 1 0 18124 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1450_
timestamp 1688980957
transform 1 0 20424 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1451_
timestamp 1688980957
transform 1 0 18400 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1452_
timestamp 1688980957
transform 1 0 21252 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1453_
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1454_
timestamp 1688980957
transform 1 0 25208 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1455_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23552 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1688980957
transform 1 0 20608 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1457_
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1458_
timestamp 1688980957
transform 1 0 20700 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1459_
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1460_
timestamp 1688980957
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1461_
timestamp 1688980957
transform 1 0 32844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1462_
timestamp 1688980957
transform 1 0 33120 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1463_
timestamp 1688980957
transform 1 0 33580 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1464_
timestamp 1688980957
transform 1 0 14536 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1465_
timestamp 1688980957
transform 1 0 14168 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1466_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1467_
timestamp 1688980957
transform 1 0 18124 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1688980957
transform 1 0 15732 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1469_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1470_
timestamp 1688980957
transform 1 0 12880 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1471_
timestamp 1688980957
transform 1 0 13064 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1472_
timestamp 1688980957
transform 1 0 13984 0 -1 27200
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_8  _1473_
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__and3_2  _1474_
timestamp 1688980957
transform 1 0 20424 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1475_
timestamp 1688980957
transform 1 0 16192 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1476_
timestamp 1688980957
transform 1 0 17020 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1477_
timestamp 1688980957
transform 1 0 17204 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1478_
timestamp 1688980957
transform 1 0 18768 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1479_
timestamp 1688980957
transform 1 0 17112 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1480_
timestamp 1688980957
transform 1 0 17756 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1481_
timestamp 1688980957
transform 1 0 18216 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1482_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1483_
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1484_
timestamp 1688980957
transform 1 0 17572 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1485_
timestamp 1688980957
transform 1 0 18584 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1487_
timestamp 1688980957
transform 1 0 17848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_4  _1488_
timestamp 1688980957
transform 1 0 17112 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _1489_
timestamp 1688980957
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1490_
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1491_
timestamp 1688980957
transform 1 0 16928 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1492_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1493_
timestamp 1688980957
transform 1 0 17572 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1494_
timestamp 1688980957
transform 1 0 17112 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1495_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1496_
timestamp 1688980957
transform 1 0 18768 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1497_
timestamp 1688980957
transform 1 0 16100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1498_
timestamp 1688980957
transform 1 0 16652 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1499_
timestamp 1688980957
transform 1 0 17940 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1500_
timestamp 1688980957
transform 1 0 18032 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _1501_
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1502_
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1503_
timestamp 1688980957
transform 1 0 14352 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1504_
timestamp 1688980957
transform 1 0 14536 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp 1688980957
transform 1 0 15640 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1506_
timestamp 1688980957
transform 1 0 18216 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1507_
timestamp 1688980957
transform 1 0 14628 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1508_
timestamp 1688980957
transform 1 0 12236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1509_
timestamp 1688980957
transform 1 0 12420 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1510_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1511_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1512_
timestamp 1688980957
transform 1 0 19412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1513_
timestamp 1688980957
transform 1 0 30176 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1514_
timestamp 1688980957
transform 1 0 14168 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1515_
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1516_
timestamp 1688980957
transform 1 0 14444 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1517_
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1518_
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1688980957
transform 1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1521_
timestamp 1688980957
transform 1 0 12144 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1522_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12328 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1523_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19688 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_4  _1524_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1525_
timestamp 1688980957
transform 1 0 19044 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1526_
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1527_
timestamp 1688980957
transform 1 0 18032 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1528_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1529_
timestamp 1688980957
transform 1 0 17388 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1530_
timestamp 1688980957
transform 1 0 16836 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1531_
timestamp 1688980957
transform 1 0 16100 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _1532_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1533_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1534_
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1535_
timestamp 1688980957
transform 1 0 17112 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1536_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _1537_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18124 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1538_
timestamp 1688980957
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1539_
timestamp 1688980957
transform 1 0 19872 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1540_
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1542_
timestamp 1688980957
transform 1 0 17296 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1688980957
transform 1 0 22816 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1544_
timestamp 1688980957
transform 1 0 20976 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1545_
timestamp 1688980957
transform 1 0 22080 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1546_
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1548_
timestamp 1688980957
transform 1 0 22632 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1549_
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1550_
timestamp 1688980957
transform 1 0 19780 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1551_
timestamp 1688980957
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1552_
timestamp 1688980957
transform 1 0 20424 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1553_
timestamp 1688980957
transform 1 0 20424 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _1554_
timestamp 1688980957
transform 1 0 19596 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1555_
timestamp 1688980957
transform 1 0 20240 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _1556_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1557_
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1558_
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1559_
timestamp 1688980957
transform 1 0 20608 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1560_
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1561_
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1688980957
transform 1 0 15824 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1563_
timestamp 1688980957
transform 1 0 16100 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1564_
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1565_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1566_
timestamp 1688980957
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1567_
timestamp 1688980957
transform 1 0 19780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1568_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1569_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1570_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1571_
timestamp 1688980957
transform 1 0 22816 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1572_
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1573_
timestamp 1688980957
transform 1 0 22632 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1574_
timestamp 1688980957
transform 1 0 23368 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1575_
timestamp 1688980957
transform 1 0 23000 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1576_
timestamp 1688980957
transform 1 0 20148 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1688980957
transform 1 0 20516 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1578_
timestamp 1688980957
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1579_
timestamp 1688980957
transform 1 0 25576 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1580_
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1581_
timestamp 1688980957
transform 1 0 23644 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1688980957
transform 1 0 22264 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1583_
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 1688980957
transform 1 0 22264 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1585_
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1586_
timestamp 1688980957
transform 1 0 23460 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1688980957
transform 1 0 19044 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1588_
timestamp 1688980957
transform 1 0 19412 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1589_
timestamp 1688980957
transform 1 0 20056 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1590_
timestamp 1688980957
transform 1 0 19504 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1591_
timestamp 1688980957
transform 1 0 21988 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1592_
timestamp 1688980957
transform 1 0 28980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1593_
timestamp 1688980957
transform 1 0 28888 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1594_
timestamp 1688980957
transform 1 0 31924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1595_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1596_
timestamp 1688980957
transform 1 0 22080 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1597_
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1598_
timestamp 1688980957
transform 1 0 22540 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1599_
timestamp 1688980957
transform 1 0 22724 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1600_
timestamp 1688980957
transform 1 0 23092 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1601_
timestamp 1688980957
transform 1 0 22172 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 1688980957
transform 1 0 23460 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1603_
timestamp 1688980957
transform 1 0 22724 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1604_
timestamp 1688980957
transform 1 0 24288 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1605_
timestamp 1688980957
transform 1 0 23736 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1606_
timestamp 1688980957
transform 1 0 22724 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1688980957
transform 1 0 22540 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1608_
timestamp 1688980957
transform 1 0 21252 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1688980957
transform 1 0 21896 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1610_
timestamp 1688980957
transform 1 0 22908 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1611_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23552 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1612_
timestamp 1688980957
transform 1 0 22908 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1613_
timestamp 1688980957
transform 1 0 20424 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1614_
timestamp 1688980957
transform 1 0 20976 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1615_
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _1616_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _1617_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__a22oi_1  _1618_
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1619_
timestamp 1688980957
transform 1 0 14352 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1620_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15548 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1621_
timestamp 1688980957
transform 1 0 19688 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1688980957
transform 1 0 14720 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1623_
timestamp 1688980957
transform 1 0 14904 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1624_
timestamp 1688980957
transform 1 0 12880 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _1626_
timestamp 1688980957
transform 1 0 12880 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _1627_
timestamp 1688980957
transform 1 0 25852 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1628_
timestamp 1688980957
transform 1 0 19872 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1629_
timestamp 1688980957
transform 1 0 19412 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1630_
timestamp 1688980957
transform 1 0 17296 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1631_
timestamp 1688980957
transform 1 0 18216 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1688980957
transform 1 0 18768 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1633_
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1634_
timestamp 1688980957
transform 1 0 19412 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1635_
timestamp 1688980957
transform 1 0 19780 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1637_
timestamp 1688980957
transform 1 0 18400 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1638_
timestamp 1688980957
transform 1 0 19320 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_4  _1639_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_2  _1640_
timestamp 1688980957
transform 1 0 29072 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1641_
timestamp 1688980957
transform 1 0 30544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1642_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31832 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1643_
timestamp 1688980957
transform 1 0 26312 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1644_
timestamp 1688980957
transform 1 0 26036 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1645_
timestamp 1688980957
transform 1 0 26496 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1646_
timestamp 1688980957
transform 1 0 30636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1647_
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 1688980957
transform 1 0 33120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1688980957
transform 1 0 31556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1650_
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1651_
timestamp 1688980957
transform 1 0 32384 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1652_
timestamp 1688980957
transform 1 0 35972 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1688980957
transform 1 0 35236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1654_
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1655_
timestamp 1688980957
transform 1 0 34776 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1656_
timestamp 1688980957
transform 1 0 35144 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1657_
timestamp 1688980957
transform 1 0 34408 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1658_
timestamp 1688980957
transform 1 0 29624 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1659_
timestamp 1688980957
transform 1 0 30360 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1660_
timestamp 1688980957
transform 1 0 30912 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1688980957
transform 1 0 25392 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1662_
timestamp 1688980957
transform 1 0 25576 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1663_
timestamp 1688980957
transform 1 0 25300 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1664_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1665_
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1688980957
transform 1 0 33120 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1667_
timestamp 1688980957
transform 1 0 32384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1668_
timestamp 1688980957
transform 1 0 32660 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1669_
timestamp 1688980957
transform 1 0 29624 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1670_
timestamp 1688980957
transform 1 0 30360 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _1671_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30544 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1688980957
transform 1 0 25392 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1673_
timestamp 1688980957
transform 1 0 26036 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1674_
timestamp 1688980957
transform 1 0 25760 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1688980957
transform 1 0 26680 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1676_
timestamp 1688980957
transform 1 0 30728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1677_
timestamp 1688980957
transform 1 0 31648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1678_
timestamp 1688980957
transform 1 0 31004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1679_
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1680_
timestamp 1688980957
transform 1 0 32292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1681_
timestamp 1688980957
transform 1 0 31832 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1682_
timestamp 1688980957
transform 1 0 31372 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1683_
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1684_
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1685_
timestamp 1688980957
transform 1 0 29256 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1686_
timestamp 1688980957
transform 1 0 28612 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1687_
timestamp 1688980957
transform 1 0 25208 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1688_
timestamp 1688980957
transform 1 0 25208 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1689_
timestamp 1688980957
transform 1 0 25392 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1690_
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1691_
timestamp 1688980957
transform 1 0 28336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1692_
timestamp 1688980957
transform 1 0 27784 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1688980957
transform 1 0 29072 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1694_
timestamp 1688980957
transform 1 0 28612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1695_
timestamp 1688980957
transform 1 0 29440 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1696_
timestamp 1688980957
transform 1 0 20792 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1697_
timestamp 1688980957
transform 1 0 19596 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1698_
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1699_
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1700_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_2  _1701_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1702_
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1703_
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1704_
timestamp 1688980957
transform 1 0 20516 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_4  _1705_
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_8  _1706_
timestamp 1688980957
transform 1 0 22356 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _1707_
timestamp 1688980957
transform 1 0 27140 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1708_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1688980957
transform 1 0 34684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1688980957
transform 1 0 33856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1711_
timestamp 1688980957
transform 1 0 34960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1712_
timestamp 1688980957
transform 1 0 32844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1713_
timestamp 1688980957
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1714_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1715_
timestamp 1688980957
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1716_
timestamp 1688980957
transform 1 0 20700 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _1717_
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1718_
timestamp 1688980957
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1719_
timestamp 1688980957
transform 1 0 25944 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1720_
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1721_
timestamp 1688980957
transform 1 0 28796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1722_
timestamp 1688980957
transform 1 0 29716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1723_
timestamp 1688980957
transform 1 0 24564 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1724_
timestamp 1688980957
transform 1 0 25484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1725_
timestamp 1688980957
transform 1 0 25392 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1726_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1727_
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1728_
timestamp 1688980957
transform 1 0 27048 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _1729_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22632 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1731_
timestamp 1688980957
transform 1 0 27600 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1732_
timestamp 1688980957
transform 1 0 25760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1733_
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1734_
timestamp 1688980957
transform 1 0 26864 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1735_
timestamp 1688980957
transform 1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1736_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1737_
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1738_
timestamp 1688980957
transform 1 0 33764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1739_
timestamp 1688980957
transform 1 0 34408 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1740_
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1741_
timestamp 1688980957
transform 1 0 34592 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1742_
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1743_
timestamp 1688980957
transform 1 0 31280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1744_
timestamp 1688980957
transform 1 0 32476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1745_
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1746_
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1747_
timestamp 1688980957
transform 1 0 28704 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1748_
timestamp 1688980957
transform 1 0 21896 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1749_
timestamp 1688980957
transform 1 0 23276 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1750_
timestamp 1688980957
transform 1 0 25300 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_4  _1751_
timestamp 1688980957
transform 1 0 29440 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1752_
timestamp 1688980957
transform 1 0 29624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1753_
timestamp 1688980957
transform 1 0 30268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp 1688980957
transform 1 0 30544 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1755_
timestamp 1688980957
transform 1 0 31188 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1756_
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1757_
timestamp 1688980957
transform 1 0 29716 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1758_
timestamp 1688980957
transform 1 0 33488 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1759_
timestamp 1688980957
transform 1 0 33856 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1760_
timestamp 1688980957
transform 1 0 33764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1761_
timestamp 1688980957
transform 1 0 29624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1762_
timestamp 1688980957
transform 1 0 31556 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1688980957
transform 1 0 25576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1764_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1765_
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1766_
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1767_
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1768_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19136 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1769_
timestamp 1688980957
transform 1 0 25392 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1770_
timestamp 1688980957
transform 1 0 29992 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1771_
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1772_
timestamp 1688980957
transform 1 0 31004 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1773_
timestamp 1688980957
transform 1 0 31924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1774_
timestamp 1688980957
transform 1 0 32844 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1775_
timestamp 1688980957
transform 1 0 33120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1776_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33212 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1777_
timestamp 1688980957
transform 1 0 33396 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1778_
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _1779_
timestamp 1688980957
transform 1 0 20240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1780_
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1781_
timestamp 1688980957
transform 1 0 28888 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1782_
timestamp 1688980957
transform 1 0 33488 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1783_
timestamp 1688980957
transform 1 0 33028 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1784_
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1785_
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1786_
timestamp 1688980957
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1787_
timestamp 1688980957
transform 1 0 28612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1788_
timestamp 1688980957
transform 1 0 30544 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1789_
timestamp 1688980957
transform 1 0 33120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1790_
timestamp 1688980957
transform 1 0 29624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1791_
timestamp 1688980957
transform 1 0 31096 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1792_
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1793_
timestamp 1688980957
transform 1 0 29900 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1794_
timestamp 1688980957
transform 1 0 22172 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1795_
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1796_
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1797_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1798_
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1799_
timestamp 1688980957
transform 1 0 22172 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1800_
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1801_
timestamp 1688980957
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1802_
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1803_
timestamp 1688980957
transform 1 0 28244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1804_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1805_
timestamp 1688980957
transform 1 0 31280 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1806_
timestamp 1688980957
transform 1 0 29256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1807_
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1808_
timestamp 1688980957
transform 1 0 21344 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a2111oi_1  _1809_
timestamp 1688980957
transform 1 0 28244 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1810_
timestamp 1688980957
transform 1 0 28612 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1811_
timestamp 1688980957
transform 1 0 30728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1812_
timestamp 1688980957
transform 1 0 32568 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1813_
timestamp 1688980957
transform 1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1814_
timestamp 1688980957
transform 1 0 28152 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1815_
timestamp 1688980957
transform 1 0 27324 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1816_
timestamp 1688980957
transform 1 0 20976 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1817_
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1818_
timestamp 1688980957
transform 1 0 23276 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1819_
timestamp 1688980957
transform 1 0 22448 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1820_
timestamp 1688980957
transform 1 0 20240 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1821_
timestamp 1688980957
transform 1 0 23092 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1822_
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1823_
timestamp 1688980957
transform 1 0 32936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1824_
timestamp 1688980957
transform 1 0 23092 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _1825_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1826_
timestamp 1688980957
transform 1 0 25576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1827_
timestamp 1688980957
transform 1 0 24656 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1828_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1829_
timestamp 1688980957
transform 1 0 21160 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1830_
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1831_
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1832_
timestamp 1688980957
transform 1 0 22632 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1833_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25024 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1834_
timestamp 1688980957
transform 1 0 25024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1835_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1836_
timestamp 1688980957
transform 1 0 25024 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1837_
timestamp 1688980957
transform 1 0 27324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1838_
timestamp 1688980957
transform 1 0 28428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1839_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1840_
timestamp 1688980957
transform 1 0 25668 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1841_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1842_
timestamp 1688980957
transform 1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1843_
timestamp 1688980957
transform 1 0 14904 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1844_
timestamp 1688980957
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _1845_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1846_
timestamp 1688980957
transform 1 0 15548 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1847_
timestamp 1688980957
transform 1 0 14628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1848_
timestamp 1688980957
transform 1 0 13800 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1849_
timestamp 1688980957
transform 1 0 14720 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1850_
timestamp 1688980957
transform 1 0 14628 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1851_
timestamp 1688980957
transform 1 0 14904 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1852_
timestamp 1688980957
transform 1 0 16376 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1853_
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1854_
timestamp 1688980957
transform 1 0 15456 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1855_
timestamp 1688980957
transform 1 0 15364 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1856_
timestamp 1688980957
transform 1 0 15088 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1857_
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1858_
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_4  _1859_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_4  _1860_
timestamp 1688980957
transform 1 0 14996 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1861_
timestamp 1688980957
transform 1 0 33396 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1862_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34224 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1863_
timestamp 1688980957
transform 1 0 33120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1864_
timestamp 1688980957
transform 1 0 32660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1865_
timestamp 1688980957
transform 1 0 28428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1867_
timestamp 1688980957
transform 1 0 31556 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1868_
timestamp 1688980957
transform 1 0 24564 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1869_
timestamp 1688980957
transform 1 0 30820 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1870_
timestamp 1688980957
transform 1 0 30728 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1871_
timestamp 1688980957
transform 1 0 23828 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _1872_
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1873_
timestamp 1688980957
transform 1 0 25668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1874_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26036 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1875_
timestamp 1688980957
transform 1 0 26220 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1876_
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1877_
timestamp 1688980957
transform 1 0 30452 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1878_
timestamp 1688980957
transform 1 0 31556 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1879_
timestamp 1688980957
transform 1 0 31188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1880_
timestamp 1688980957
transform 1 0 29992 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1881_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29440 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1882_
timestamp 1688980957
transform 1 0 29808 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1883_
timestamp 1688980957
transform 1 0 26680 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1884_
timestamp 1688980957
transform 1 0 26036 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1885_
timestamp 1688980957
transform 1 0 26404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1886_
timestamp 1688980957
transform 1 0 31556 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1887_
timestamp 1688980957
transform 1 0 31188 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1888_
timestamp 1688980957
transform 1 0 32476 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1889_
timestamp 1688980957
transform 1 0 25668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1890_
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1891_
timestamp 1688980957
transform 1 0 26220 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1892_
timestamp 1688980957
transform 1 0 26680 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1893_
timestamp 1688980957
transform 1 0 30176 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1894_
timestamp 1688980957
transform 1 0 32660 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1895_
timestamp 1688980957
transform 1 0 28520 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1896_
timestamp 1688980957
transform 1 0 32476 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1897_
timestamp 1688980957
transform 1 0 32568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1898_
timestamp 1688980957
transform 1 0 30452 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1899_
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1900_
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1901_
timestamp 1688980957
transform 1 0 31188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1902_
timestamp 1688980957
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1903_
timestamp 1688980957
transform 1 0 32016 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1904_
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1905_
timestamp 1688980957
transform 1 0 30912 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1906_
timestamp 1688980957
transform 1 0 27508 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1907_
timestamp 1688980957
transform 1 0 31188 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1908_
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1909_
timestamp 1688980957
transform 1 0 31004 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1910_
timestamp 1688980957
transform 1 0 29440 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1911_
timestamp 1688980957
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1912_
timestamp 1688980957
transform 1 0 30728 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1914_
timestamp 1688980957
transform 1 0 23368 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1915_
timestamp 1688980957
transform 1 0 21620 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1916_
timestamp 1688980957
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1917_
timestamp 1688980957
transform 1 0 26036 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1918_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1919_
timestamp 1688980957
transform 1 0 26864 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1920_
timestamp 1688980957
transform 1 0 24472 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1921_
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1922_
timestamp 1688980957
transform 1 0 28152 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _1923_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1924_
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1925_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30728 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _1926_
timestamp 1688980957
transform 1 0 33120 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1927_
timestamp 1688980957
transform 1 0 32752 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1928_
timestamp 1688980957
transform 1 0 32384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1929_
timestamp 1688980957
transform 1 0 28152 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1930_
timestamp 1688980957
transform 1 0 33488 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1931_
timestamp 1688980957
transform 1 0 34040 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1932_
timestamp 1688980957
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 1688980957
transform 1 0 27416 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1934_
timestamp 1688980957
transform 1 0 27784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1935_
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1936_
timestamp 1688980957
transform 1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1937_
timestamp 1688980957
transform 1 0 28152 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _1938_
timestamp 1688980957
transform 1 0 25300 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1939_
timestamp 1688980957
transform 1 0 25944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1940_
timestamp 1688980957
transform 1 0 26772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1941_
timestamp 1688980957
transform 1 0 27140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1942_
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1943_
timestamp 1688980957
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1944_
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1945_
timestamp 1688980957
transform 1 0 28428 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1946_
timestamp 1688980957
transform 1 0 35512 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1947_
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1948_
timestamp 1688980957
transform 1 0 34132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1949_
timestamp 1688980957
transform 1 0 33856 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1950_
timestamp 1688980957
transform 1 0 27324 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1951_
timestamp 1688980957
transform 1 0 33764 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1952_
timestamp 1688980957
transform 1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1953_
timestamp 1688980957
transform 1 0 22816 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1954_
timestamp 1688980957
transform 1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1955_
timestamp 1688980957
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1956_
timestamp 1688980957
transform 1 0 24748 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1957_
timestamp 1688980957
transform 1 0 20148 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1958_
timestamp 1688980957
transform 1 0 21252 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1959_
timestamp 1688980957
transform 1 0 25760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1960_
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1961_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1962_
timestamp 1688980957
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1963_
timestamp 1688980957
transform 1 0 24748 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1964_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1965_
timestamp 1688980957
transform 1 0 24656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1966_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_4  _1967_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23000 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1968_
timestamp 1688980957
transform 1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1969_
timestamp 1688980957
transform 1 0 34776 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1970_
timestamp 1688980957
transform 1 0 35144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1971_
timestamp 1688980957
transform 1 0 35604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1972_
timestamp 1688980957
transform 1 0 24104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1973_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1974_
timestamp 1688980957
transform 1 0 33304 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1975_
timestamp 1688980957
transform 1 0 34132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1976_
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1977_
timestamp 1688980957
transform 1 0 21988 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1978_
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1979_
timestamp 1688980957
transform 1 0 20056 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1980_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1981_
timestamp 1688980957
transform 1 0 19504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1982_
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1983_
timestamp 1688980957
transform 1 0 22172 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1984_
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1985_
timestamp 1688980957
transform 1 0 23000 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1986_
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1987_
timestamp 1688980957
transform 1 0 22448 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_4  _1988_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22448 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_1  _1989_
timestamp 1688980957
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1990_
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1991_
timestamp 1688980957
transform 1 0 35512 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1992_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1993_
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1994_
timestamp 1688980957
transform 1 0 26036 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1995_
timestamp 1688980957
transform 1 0 26036 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1996_
timestamp 1688980957
transform 1 0 26404 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1997_
timestamp 1688980957
transform 1 0 20608 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1998_
timestamp 1688980957
transform 1 0 20608 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1999_
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2000_
timestamp 1688980957
transform 1 0 21160 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2001_
timestamp 1688980957
transform 1 0 21068 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2002_
timestamp 1688980957
transform 1 0 22816 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2003_
timestamp 1688980957
transform 1 0 22724 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2004_
timestamp 1688980957
transform 1 0 22448 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2005_
timestamp 1688980957
transform 1 0 24380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2006_
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2007_
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _2008_
timestamp 1688980957
transform 1 0 22080 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2009_
timestamp 1688980957
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2010_
timestamp 1688980957
transform 1 0 31188 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2011_
timestamp 1688980957
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2012_
timestamp 1688980957
transform 1 0 31372 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2013_
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2014_
timestamp 1688980957
transform 1 0 23736 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2015_
timestamp 1688980957
transform 1 0 28336 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2016_
timestamp 1688980957
transform 1 0 28796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2017_
timestamp 1688980957
transform 1 0 13984 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2018_
timestamp 1688980957
transform 1 0 26956 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2019_
timestamp 1688980957
transform 1 0 28796 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2020_
timestamp 1688980957
transform 1 0 29624 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2021_
timestamp 1688980957
transform 1 0 27048 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2022_
timestamp 1688980957
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2023_
timestamp 1688980957
transform 1 0 28152 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2024_
timestamp 1688980957
transform 1 0 27876 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2025_
timestamp 1688980957
transform 1 0 28704 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2026_
timestamp 1688980957
transform 1 0 28980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2027_
timestamp 1688980957
transform 1 0 28336 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2028_
timestamp 1688980957
transform 1 0 28612 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2029_
timestamp 1688980957
transform 1 0 27508 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2030_
timestamp 1688980957
transform 1 0 27416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2031_
timestamp 1688980957
transform 1 0 26956 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2032_
timestamp 1688980957
transform 1 0 26312 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2033_
timestamp 1688980957
transform 1 0 28244 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2034_
timestamp 1688980957
transform 1 0 28428 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2035_
timestamp 1688980957
transform 1 0 14812 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _2036_
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and4_2  _2037_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _2038_
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2039_
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2040_
timestamp 1688980957
transform 1 0 13432 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2041_
timestamp 1688980957
transform 1 0 13984 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2042_
timestamp 1688980957
transform 1 0 12880 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _2043_
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_4  _2044_
timestamp 1688980957
transform 1 0 12696 0 -1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2045_
timestamp 1688980957
transform 1 0 9476 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2046_
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2047_
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2048_
timestamp 1688980957
transform 1 0 10580 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2049_
timestamp 1688980957
transform 1 0 10304 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2050_
timestamp 1688980957
transform 1 0 9016 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2051_
timestamp 1688980957
transform 1 0 7820 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2052_
timestamp 1688980957
transform 1 0 7544 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2053_
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2054_
timestamp 1688980957
transform 1 0 7636 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2055_
timestamp 1688980957
transform 1 0 7176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2056_
timestamp 1688980957
transform 1 0 9568 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2057_
timestamp 1688980957
transform 1 0 10580 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2058_
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2059_
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2060_
timestamp 1688980957
transform 1 0 11592 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2061_
timestamp 1688980957
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2062_
timestamp 1688980957
transform 1 0 9016 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2063_
timestamp 1688980957
transform 1 0 7820 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2064_
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2065_
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2066_
timestamp 1688980957
transform 1 0 9752 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2067_
timestamp 1688980957
transform 1 0 8372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2068_
timestamp 1688980957
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _2069_
timestamp 1688980957
transform 1 0 12604 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2070_
timestamp 1688980957
transform 1 0 12788 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2071_
timestamp 1688980957
transform 1 0 13156 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2072_
timestamp 1688980957
transform 1 0 30728 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2073_
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2074_
timestamp 1688980957
transform 1 0 25760 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2075_
timestamp 1688980957
transform 1 0 25484 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2076_
timestamp 1688980957
transform 1 0 32936 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2077_
timestamp 1688980957
transform 1 0 34040 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2078_
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2079_
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2080_
timestamp 1688980957
transform 1 0 34040 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2081_
timestamp 1688980957
transform 1 0 34132 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2082_
timestamp 1688980957
transform 1 0 27140 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2083_
timestamp 1688980957
transform 1 0 27048 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2084_
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2085_
timestamp 1688980957
transform 1 0 30728 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2086_
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2087_
timestamp 1688980957
transform 1 0 24472 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2088_
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2089_
timestamp 1688980957
transform 1 0 20424 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2090_
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2091_
timestamp 1688980957
transform 1 0 12236 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2092_
timestamp 1688980957
transform 1 0 12512 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2093_
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2094_
timestamp 1688980957
transform 1 0 4876 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2095_
timestamp 1688980957
transform 1 0 5428 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2096_
timestamp 1688980957
transform 1 0 4692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2097_
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2098_
timestamp 1688980957
transform 1 0 7728 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2099_
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2100_
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2101_
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2102_
timestamp 1688980957
transform 1 0 5520 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2103_
timestamp 1688980957
transform 1 0 6440 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2104_
timestamp 1688980957
transform 1 0 5704 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2105_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2106_
timestamp 1688980957
transform 1 0 13984 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2107_
timestamp 1688980957
transform 1 0 32752 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2108_
timestamp 1688980957
transform 1 0 32752 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2109_
timestamp 1688980957
transform 1 0 27232 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2110_
timestamp 1688980957
transform 1 0 27232 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2111_
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2112_
timestamp 1688980957
transform 1 0 33672 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2113_
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2114_
timestamp 1688980957
transform 1 0 31740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2115_
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2116_
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2117_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2118_
timestamp 1688980957
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2119_
timestamp 1688980957
transform 1 0 30912 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2120_
timestamp 1688980957
transform 1 0 30636 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2121_
timestamp 1688980957
transform 1 0 24472 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2122_
timestamp 1688980957
transform 1 0 24656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2123_
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2124_
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2125_
timestamp 1688980957
transform 1 0 10580 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2126_
timestamp 1688980957
transform 1 0 9752 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2127_
timestamp 1688980957
transform 1 0 9292 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2128_
timestamp 1688980957
transform 1 0 5704 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2129_
timestamp 1688980957
transform 1 0 5152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2130_
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2131_
timestamp 1688980957
transform 1 0 4968 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2132_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2133_
timestamp 1688980957
transform 1 0 10672 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2134_
timestamp 1688980957
transform 1 0 9936 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2135_
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2136_
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2137_
timestamp 1688980957
transform 1 0 5336 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2138_
timestamp 1688980957
transform 1 0 7176 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2139_
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2140_
timestamp 1688980957
transform 1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2141_
timestamp 1688980957
transform 1 0 24380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2142_
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2143_
timestamp 1688980957
transform 1 0 16008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2144_
timestamp 1688980957
transform 1 0 15824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2145_
timestamp 1688980957
transform 1 0 15364 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2146_
timestamp 1688980957
transform 1 0 14720 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2147_
timestamp 1688980957
transform 1 0 14168 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_4  _2148_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__a31o_2  _2149_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2150_
timestamp 1688980957
transform 1 0 9292 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2151_
timestamp 1688980957
transform 1 0 8372 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2152_
timestamp 1688980957
transform 1 0 10028 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2153_
timestamp 1688980957
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2154_
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2155_
timestamp 1688980957
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2156_
timestamp 1688980957
transform 1 0 21896 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2157_
timestamp 1688980957
transform 1 0 23184 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _2158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2159_
timestamp 1688980957
transform 1 0 10672 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2160_
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2161_
timestamp 1688980957
transform 1 0 10120 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2162_
timestamp 1688980957
transform 1 0 7452 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2163_
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2164_
timestamp 1688980957
transform 1 0 8280 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2165_
timestamp 1688980957
transform 1 0 30912 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2166_
timestamp 1688980957
transform 1 0 29808 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2167_
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2168_
timestamp 1688980957
transform 1 0 30176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2169_
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2170_
timestamp 1688980957
transform 1 0 24564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2171_
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2172_
timestamp 1688980957
transform 1 0 24196 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2173_
timestamp 1688980957
transform 1 0 24932 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2174_
timestamp 1688980957
transform 1 0 33120 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2175_
timestamp 1688980957
transform 1 0 33488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2176_
timestamp 1688980957
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2177_
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2178_
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2179_
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2180_
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2181_
timestamp 1688980957
transform 1 0 32108 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2182_
timestamp 1688980957
transform 1 0 32752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2183_
timestamp 1688980957
transform 1 0 33120 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2184_
timestamp 1688980957
transform 1 0 33672 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2185_
timestamp 1688980957
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2186_
timestamp 1688980957
transform 1 0 28244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2187_
timestamp 1688980957
transform 1 0 30452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2188_
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2189_
timestamp 1688980957
transform 1 0 31924 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2190_
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2191_
timestamp 1688980957
transform 1 0 33764 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2192_
timestamp 1688980957
transform 1 0 33948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2193_
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2194_
timestamp 1688980957
transform 1 0 34776 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2195_
timestamp 1688980957
transform 1 0 35236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_4  _2196_
timestamp 1688980957
transform 1 0 28336 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _2197_
timestamp 1688980957
transform 1 0 27968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2198_
timestamp 1688980957
transform 1 0 29072 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2199_
timestamp 1688980957
transform 1 0 23000 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2200_
timestamp 1688980957
transform 1 0 23644 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2201_
timestamp 1688980957
transform 1 0 23552 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2202_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2203_
timestamp 1688980957
transform 1 0 25208 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2204_
timestamp 1688980957
transform 1 0 25852 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2205_
timestamp 1688980957
transform 1 0 26496 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2206_
timestamp 1688980957
transform 1 0 27232 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_4  _2207_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2208_
timestamp 1688980957
transform 1 0 11224 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2209_
timestamp 1688980957
transform 1 0 11592 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2210_
timestamp 1688980957
transform 1 0 10212 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2211_
timestamp 1688980957
transform 1 0 10396 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2212_
timestamp 1688980957
transform 1 0 9752 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2213_
timestamp 1688980957
transform 1 0 30360 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2214_
timestamp 1688980957
transform 1 0 29992 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2215_
timestamp 1688980957
transform 1 0 29072 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2216_
timestamp 1688980957
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2217_
timestamp 1688980957
transform 1 0 22632 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2218_
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _2219_
timestamp 1688980957
transform 1 0 28612 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2220_
timestamp 1688980957
transform 1 0 28336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2221_
timestamp 1688980957
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2222_
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2223_
timestamp 1688980957
transform 1 0 28612 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2224_
timestamp 1688980957
transform 1 0 28336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _2225_
timestamp 1688980957
transform 1 0 28336 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2226_
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2227_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2228_
timestamp 1688980957
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2229_
timestamp 1688980957
transform 1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2230_
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2231_
timestamp 1688980957
transform 1 0 11592 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2232_
timestamp 1688980957
transform 1 0 12144 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2233_
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2234_
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2235_
timestamp 1688980957
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _2236_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2237_
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2238_
timestamp 1688980957
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2239_
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2240_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2241_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _2242_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2243_
timestamp 1688980957
transform 1 0 12328 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2244_
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2245_
timestamp 1688980957
transform 1 0 9108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2246_
timestamp 1688980957
transform 1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2247_
timestamp 1688980957
transform 1 0 9108 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2248_
timestamp 1688980957
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2249_
timestamp 1688980957
transform 1 0 9568 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2250_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2251_
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2252_
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2253_
timestamp 1688980957
transform 1 0 8464 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2254_
timestamp 1688980957
transform 1 0 10212 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2255_
timestamp 1688980957
transform 1 0 8188 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2256_
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _2257_
timestamp 1688980957
transform 1 0 7912 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _2258_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8648 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _2259_
timestamp 1688980957
transform 1 0 7820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2260_
timestamp 1688980957
transform 1 0 10304 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2261_
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2262_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2263_
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2264_
timestamp 1688980957
transform 1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2265_
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2266_
timestamp 1688980957
transform 1 0 13248 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2267_
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _2268_
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_4  _2269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2270_
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2271_
timestamp 1688980957
transform 1 0 15272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2272_
timestamp 1688980957
transform 1 0 14352 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2273_
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  _2274_
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2275_
timestamp 1688980957
transform 1 0 17756 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2276_
timestamp 1688980957
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2277_
timestamp 1688980957
transform 1 0 29900 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2278_
timestamp 1688980957
transform 1 0 37352 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2279_
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2280_
timestamp 1688980957
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2281_
timestamp 1688980957
transform 1 0 12144 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2282_
timestamp 1688980957
transform 1 0 9292 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2283_
timestamp 1688980957
transform 1 0 11684 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2284_
timestamp 1688980957
transform 1 0 11592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2285_
timestamp 1688980957
transform 1 0 12972 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2286_
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2287_
timestamp 1688980957
transform 1 0 12236 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2288_
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2289_
timestamp 1688980957
transform 1 0 36616 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2290_
timestamp 1688980957
transform 1 0 37352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _2291_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2292_
timestamp 1688980957
transform 1 0 1932 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2293_
timestamp 1688980957
transform 1 0 1748 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2294_
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2295_
timestamp 1688980957
transform 1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2296_
timestamp 1688980957
transform 1 0 9568 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2297_
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2298_
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2299_
timestamp 1688980957
transform 1 0 3128 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2300_
timestamp 1688980957
transform 1 0 2576 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2301_
timestamp 1688980957
transform 1 0 5704 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2302_
timestamp 1688980957
transform 1 0 19228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2303_
timestamp 1688980957
transform 1 0 2300 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2304_
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2305_
timestamp 1688980957
transform 1 0 4324 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2306_
timestamp 1688980957
transform 1 0 9016 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2307_
timestamp 1688980957
transform 1 0 3220 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2308_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2309_
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2310_
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2311_
timestamp 1688980957
transform 1 0 17572 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2312_
timestamp 1688980957
transform 1 0 17296 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2313_
timestamp 1688980957
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2314_
timestamp 1688980957
transform 1 0 2668 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2315_
timestamp 1688980957
transform 1 0 2024 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2316_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2317_
timestamp 1688980957
transform 1 0 2208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2318_
timestamp 1688980957
transform 1 0 2116 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2319_
timestamp 1688980957
transform 1 0 4600 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2320_
timestamp 1688980957
transform 1 0 22632 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2321_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2322_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2323_
timestamp 1688980957
transform 1 0 7728 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2324_
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2325_
timestamp 1688980957
transform 1 0 5152 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2326_
timestamp 1688980957
transform 1 0 5244 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2327_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2328_
timestamp 1688980957
transform 1 0 2392 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2329_
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2330_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2331_
timestamp 1688980957
transform 1 0 26036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2332_
timestamp 1688980957
transform 1 0 24748 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2333_
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2334_
timestamp 1688980957
transform 1 0 25024 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2335_
timestamp 1688980957
transform 1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2336_
timestamp 1688980957
transform 1 0 26864 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2337_
timestamp 1688980957
transform 1 0 37168 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2338_
timestamp 1688980957
transform 1 0 24840 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2339_
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2340_
timestamp 1688980957
transform 1 0 26956 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2341_
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2342_
timestamp 1688980957
transform 1 0 27876 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2343_
timestamp 1688980957
transform 1 0 32108 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2344_
timestamp 1688980957
transform 1 0 24564 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2345_
timestamp 1688980957
transform 1 0 4968 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2346_
timestamp 1688980957
transform 1 0 25024 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2347_
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2348_
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2349_
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2350_
timestamp 1688980957
transform 1 0 7268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2351_
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2352_
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2353_
timestamp 1688980957
transform 1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2354_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2355_
timestamp 1688980957
transform 1 0 5244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2356_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2357_
timestamp 1688980957
transform 1 0 5704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2358_
timestamp 1688980957
transform 1 0 6624 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2359_
timestamp 1688980957
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2360_
timestamp 1688980957
transform 1 0 8924 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2361_
timestamp 1688980957
transform 1 0 7728 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2362_
timestamp 1688980957
transform 1 0 7360 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2363_
timestamp 1688980957
transform 1 0 8004 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2364_
timestamp 1688980957
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2365_
timestamp 1688980957
transform 1 0 6900 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2366_
timestamp 1688980957
transform 1 0 6532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2367_
timestamp 1688980957
transform 1 0 6440 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2368_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2369_
timestamp 1688980957
transform 1 0 7636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2370_
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2371_
timestamp 1688980957
transform 1 0 11500 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2372_
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2373_
timestamp 1688980957
transform 1 0 14536 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2374_
timestamp 1688980957
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2375_
timestamp 1688980957
transform 1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2376_
timestamp 1688980957
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2377_
timestamp 1688980957
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2378_
timestamp 1688980957
transform 1 0 16192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2379_
timestamp 1688980957
transform 1 0 10580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2380_
timestamp 1688980957
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2381_
timestamp 1688980957
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2382_
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2383_
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2384_
timestamp 1688980957
transform 1 0 12880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2385_
timestamp 1688980957
transform 1 0 12696 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2386_
timestamp 1688980957
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2387_
timestamp 1688980957
transform 1 0 11592 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2388_
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2389_
timestamp 1688980957
transform 1 0 13892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2390_
timestamp 1688980957
transform 1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2391_
timestamp 1688980957
transform 1 0 14904 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2392_
timestamp 1688980957
transform 1 0 14996 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2393_
timestamp 1688980957
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2394_
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2395_
timestamp 1688980957
transform 1 0 10580 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2396_
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2397_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2398_
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 1688980957
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2400_
timestamp 1688980957
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2401_
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2402_
timestamp 1688980957
transform 1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2403_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2404_
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2405_
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2406_
timestamp 1688980957
transform 1 0 30452 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2407__8
timestamp 1688980957
transform 1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2408__9
timestamp 1688980957
transform 1 0 10120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2409__10
timestamp 1688980957
transform 1 0 9384 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2410__11
timestamp 1688980957
transform 1 0 6440 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2411__12
timestamp 1688980957
transform 1 0 7544 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2412__13
timestamp 1688980957
transform 1 0 5888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2413__14
timestamp 1688980957
transform 1 0 9568 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2414__15
timestamp 1688980957
transform 1 0 7912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2415__16
timestamp 1688980957
transform 1 0 4968 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2416__17
timestamp 1688980957
transform 1 0 4416 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2417__18
timestamp 1688980957
transform 1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2418__19
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2419__20
timestamp 1688980957
transform 1 0 4416 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2420__21
timestamp 1688980957
transform 1 0 4416 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2421__22
timestamp 1688980957
transform 1 0 9016 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2422__23
timestamp 1688980957
transform 1 0 9936 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2423__24
timestamp 1688980957
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2424__25
timestamp 1688980957
transform 1 0 30728 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2425__26
timestamp 1688980957
transform 1 0 31464 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2426_
timestamp 1688980957
transform 1 0 33488 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2427__27
timestamp 1688980957
transform 1 0 32752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2428__28
timestamp 1688980957
transform 1 0 31556 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2429__29
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2430__30
timestamp 1688980957
transform 1 0 27600 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2431__31
timestamp 1688980957
transform 1 0 32200 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2432__32
timestamp 1688980957
transform 1 0 4784 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2433__33
timestamp 1688980957
transform 1 0 4692 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2434__34
timestamp 1688980957
transform 1 0 9936 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2435__35
timestamp 1688980957
transform 1 0 7728 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2436__36
timestamp 1688980957
transform 1 0 4232 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2437__37
timestamp 1688980957
transform 1 0 3956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2438__38
timestamp 1688980957
transform 1 0 12236 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2439__39
timestamp 1688980957
transform 1 0 20240 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2440__40
timestamp 1688980957
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2441__41
timestamp 1688980957
transform 1 0 30268 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2442__42
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2443__43
timestamp 1688980957
transform 1 0 34776 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2444__44
timestamp 1688980957
transform 1 0 34132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2445__45
timestamp 1688980957
transform 1 0 33764 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2446_
timestamp 1688980957
transform 1 0 29348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2447__46
timestamp 1688980957
transform 1 0 24748 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2448__47
timestamp 1688980957
transform 1 0 31832 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2449__48
timestamp 1688980957
transform 1 0 8004 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2450__49
timestamp 1688980957
transform 1 0 6992 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2451__50
timestamp 1688980957
transform 1 0 11592 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2452__51
timestamp 1688980957
transform 1 0 9476 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2453__52
timestamp 1688980957
transform 1 0 6808 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2454__53
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2455__54
timestamp 1688980957
transform 1 0 9844 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2456__55
timestamp 1688980957
transform 1 0 8464 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2457__56
timestamp 1688980957
transform 1 0 28152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2458__57
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2459__58
timestamp 1688980957
transform 1 0 27140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2460__59
timestamp 1688980957
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2461__60
timestamp 1688980957
transform 1 0 28704 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2462__61
timestamp 1688980957
transform 1 0 28244 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2463__62
timestamp 1688980957
transform 1 0 26680 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2464__63
timestamp 1688980957
transform 1 0 29164 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2465__64
timestamp 1688980957
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2466__1
timestamp 1688980957
transform 1 0 27048 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2467__2
timestamp 1688980957
transform 1 0 34776 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2468__3
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2469__4
timestamp 1688980957
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2470__5
timestamp 1688980957
transform 1 0 31648 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2471__6
timestamp 1688980957
transform 1 0 27048 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2472__7
timestamp 1688980957
transform 1 0 34960 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2473_
timestamp 1688980957
transform 1 0 17112 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2474_
timestamp 1688980957
transform 1 0 17664 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2475_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2476_
timestamp 1688980957
transform 1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2477_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2478_
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2479_
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2480_
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2481_
timestamp 1688980957
transform 1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2482_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2483_
timestamp 1688980957
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 1688980957
transform 1 0 10304 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2485_
timestamp 1688980957
transform 1 0 10212 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2486_
timestamp 1688980957
transform 1 0 11776 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2487_
timestamp 1688980957
transform 1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _2488_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2489_
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2490_
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _2491_
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2492_
timestamp 1688980957
transform 1 0 11592 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2493_
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2494_
timestamp 1688980957
transform 1 0 11224 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2495_
timestamp 1688980957
transform 1 0 9016 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2496_
timestamp 1688980957
transform 1 0 7636 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _2497_
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _2498_
timestamp 1688980957
transform 1 0 6624 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2499_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2500_
timestamp 1688980957
transform 1 0 17572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2501_
timestamp 1688980957
transform 1 0 17204 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2502_
timestamp 1688980957
transform 1 0 4416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2503_
timestamp 1688980957
transform 1 0 4876 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 1688980957
transform 1 0 3956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2505_
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 1688980957
transform 1 0 13800 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2507_
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2508_
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2509_
timestamp 1688980957
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 1688980957
transform 1 0 3956 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2511_
timestamp 1688980957
transform 1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2512_
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2513_
timestamp 1688980957
transform 1 0 13064 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2514_
timestamp 1688980957
transform 1 0 4232 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2515_
timestamp 1688980957
transform 1 0 4692 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2516_
timestamp 1688980957
transform 1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2518_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2519_
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2520_
timestamp 1688980957
transform 1 0 18216 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2521_
timestamp 1688980957
transform 1 0 3220 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2522_
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2524_
timestamp 1688980957
transform 1 0 1748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2525_
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2526_
timestamp 1688980957
transform 1 0 12420 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2527_
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2528_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2529_
timestamp 1688980957
transform 1 0 3864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2530_
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2531_
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2532_
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2533_
timestamp 1688980957
transform 1 0 12512 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2534_
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2535_
timestamp 1688980957
transform 1 0 4600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2536_
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2537_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 1688980957
transform 1 0 2576 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2539_
timestamp 1688980957
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2541_
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 1688980957
transform 1 0 5796 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2543_
timestamp 1688980957
transform 1 0 5336 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2544_
timestamp 1688980957
transform 1 0 5060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2545_
timestamp 1688980957
transform 1 0 4508 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2546_
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2547_
timestamp 1688980957
transform 1 0 3864 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _2548_
timestamp 1688980957
transform 1 0 9200 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2549_
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2550_
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2551_
timestamp 1688980957
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2552_
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2553_
timestamp 1688980957
transform 1 0 4232 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2554_
timestamp 1688980957
transform 1 0 4140 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2555_
timestamp 1688980957
transform 1 0 3404 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2556_
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2557_
timestamp 1688980957
transform 1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2558_
timestamp 1688980957
transform 1 0 3036 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2559_
timestamp 1688980957
transform 1 0 4048 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2560_
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2561_
timestamp 1688980957
transform 1 0 2392 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2562_
timestamp 1688980957
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2563_
timestamp 1688980957
transform 1 0 4508 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2564_
timestamp 1688980957
transform 1 0 4968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2565_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2566_
timestamp 1688980957
transform 1 0 3312 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 1688980957
transform 1 0 2300 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2568_
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2569_
timestamp 1688980957
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2570_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2571_
timestamp 1688980957
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2572_
timestamp 1688980957
transform 1 0 7176 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2573_
timestamp 1688980957
transform 1 0 6900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2574_
timestamp 1688980957
transform 1 0 6992 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2575_
timestamp 1688980957
transform 1 0 7452 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2576_
timestamp 1688980957
transform 1 0 7360 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2577_
timestamp 1688980957
transform 1 0 6624 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 1688980957
transform 1 0 6624 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2579_
timestamp 1688980957
transform 1 0 5336 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2580_
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2581_
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2582_
timestamp 1688980957
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2583_
timestamp 1688980957
transform 1 0 4416 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2584_
timestamp 1688980957
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2585_
timestamp 1688980957
transform 1 0 5428 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2586_
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2587_
timestamp 1688980957
transform 1 0 5428 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2588_
timestamp 1688980957
transform 1 0 4784 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2589_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2590_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2591_
timestamp 1688980957
transform 1 0 6440 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2592_
timestamp 1688980957
transform 1 0 6164 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2593_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4600 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2594_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2595_
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2596_
timestamp 1688980957
transform 1 0 6808 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2597_
timestamp 1688980957
transform 1 0 6900 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2598_
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2599_
timestamp 1688980957
transform 1 0 5704 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2600_
timestamp 1688980957
transform 1 0 6900 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2601_
timestamp 1688980957
transform 1 0 14720 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2602_
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2603_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2604_
timestamp 1688980957
transform 1 0 10212 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2605_
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2606_
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2607_
timestamp 1688980957
transform 1 0 12696 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2608_
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2609_
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2610_
timestamp 1688980957
transform 1 0 15272 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2611_
timestamp 1688980957
transform 1 0 14352 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2612_
timestamp 1688980957
transform 1 0 10304 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 1688980957
transform 1 0 7728 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2614_
timestamp 1688980957
transform 1 0 11500 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2616_
timestamp 1688980957
transform 1 0 11040 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2617_
timestamp 1688980957
transform 1 0 9844 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2618_
timestamp 1688980957
transform 1 0 9476 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2619_
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2620_
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2621_
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2622_
timestamp 1688980957
transform 1 0 5796 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2623_
timestamp 1688980957
transform 1 0 9476 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2624_
timestamp 1688980957
transform 1 0 7820 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2625_
timestamp 1688980957
transform 1 0 5244 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2626_
timestamp 1688980957
transform 1 0 4324 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2627_
timestamp 1688980957
transform 1 0 8096 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2628_
timestamp 1688980957
transform 1 0 10304 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2629_
timestamp 1688980957
transform 1 0 4140 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2630_
timestamp 1688980957
transform 1 0 4324 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2631_
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2632_
timestamp 1688980957
transform 1 0 10212 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2633_
timestamp 1688980957
transform 1 0 24288 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2634_
timestamp 1688980957
transform 1 0 31004 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2635_
timestamp 1688980957
transform 1 0 31372 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2636_
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2637_
timestamp 1688980957
transform 1 0 31464 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2638_
timestamp 1688980957
transform 1 0 32660 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2639_
timestamp 1688980957
transform 1 0 27508 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2640_
timestamp 1688980957
transform 1 0 32476 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2641_
timestamp 1688980957
transform 1 0 5060 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2642_
timestamp 1688980957
transform 1 0 4968 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 1688980957
transform 1 0 10212 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2644_
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2645_
timestamp 1688980957
transform 1 0 4140 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2646_
timestamp 1688980957
transform 1 0 3864 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2647_
timestamp 1688980957
transform 1 0 12052 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2648_
timestamp 1688980957
transform 1 0 20516 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2649_
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2650_
timestamp 1688980957
transform 1 0 30084 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2651_
timestamp 1688980957
transform 1 0 26772 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2652_
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2653_
timestamp 1688980957
transform 1 0 34040 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2654_
timestamp 1688980957
transform 1 0 32844 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2655_
timestamp 1688980957
transform 1 0 24656 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2656_
timestamp 1688980957
transform 1 0 29992 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2657_
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2658_
timestamp 1688980957
transform 1 0 6900 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2659_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 1688980957
transform 1 0 9384 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2661_
timestamp 1688980957
transform 1 0 6716 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2662_
timestamp 1688980957
transform 1 0 6992 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2663_
timestamp 1688980957
transform 1 0 10120 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2664_
timestamp 1688980957
transform 1 0 8372 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2665_
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2666_
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2667_
timestamp 1688980957
transform 1 0 27048 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2668_
timestamp 1688980957
transform 1 0 29072 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2669_
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2670_
timestamp 1688980957
transform 1 0 28152 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2671_
timestamp 1688980957
transform 1 0 26956 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2672_
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2673_
timestamp 1688980957
transform 1 0 29072 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2674_
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2675_
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2676_
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2677_
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2678_
timestamp 1688980957
transform 1 0 31188 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2679_
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2680_
timestamp 1688980957
transform 1 0 34592 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2681_
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2682_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 1688980957
transform 1 0 2760 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 1688980957
transform 1 0 5244 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2691_
timestamp 1688980957
transform 1 0 1656 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 1688980957
transform 1 0 6440 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 1688980957
transform 1 0 4784 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 1688980957
transform 1 0 3404 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 1688980957
transform 1 0 4232 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2697_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2698_
timestamp 1688980957
transform 1 0 11868 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2699_
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2700_
timestamp 1688980957
transform 1 0 9476 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0514_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0515_
timestamp 1688980957
transform 1 0 17940 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0516_
timestamp 1688980957
transform 1 0 19412 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0517_
timestamp 1688980957
transform 1 0 19412 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1688980957
transform 1 0 13892 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0514_
timestamp 1688980957
transform 1 0 28612 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0515_
timestamp 1688980957
transform 1 0 12972 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0516_
timestamp 1688980957
transform 1 0 12972 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0517_
timestamp 1688980957
transform 1 0 12972 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0514_
timestamp 1688980957
transform 1 0 31188 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0515_
timestamp 1688980957
transform 1 0 12972 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0516_
timestamp 1688980957
transform 1 0 23368 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0517_
timestamp 1688980957
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform 1 0 5244 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout55
timestamp 1688980957
transform 1 0 2024 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout57
timestamp 1688980957
transform 1 0 2576 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout58
timestamp 1688980957
transform 1 0 5612 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout59
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout60
timestamp 1688980957
transform 1 0 22356 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout61
timestamp 1688980957
transform 1 0 25852 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_217
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_287
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_117
timestamp 1688980957
transform 1 0 11868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_132
timestamp 1688980957
transform 1 0 13248 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_156
timestamp 1688980957
transform 1 0 15456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_180
timestamp 1688980957
transform 1 0 17664 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_192
timestamp 1688980957
transform 1 0 18768 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_204
timestamp 1688980957
transform 1 0 19872 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_216
timestamp 1688980957
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_256
timestamp 1688980957
transform 1 0 24656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_268
timestamp 1688980957
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_77
timestamp 1688980957
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_87
timestamp 1688980957
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_99
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_131
timestamp 1688980957
transform 1 0 13156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_143
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_155
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_247
timestamp 1688980957
transform 1 0 23828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_259
timestamp 1688980957
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_269
timestamp 1688980957
transform 1 0 25852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_275
timestamp 1688980957
transform 1 0 26404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_289
timestamp 1688980957
transform 1 0 27692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_294
timestamp 1688980957
transform 1 0 28152 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_300
timestamp 1688980957
transform 1 0 28704 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_312
timestamp 1688980957
transform 1 0 29808 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_324
timestamp 1688980957
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_57
timestamp 1688980957
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_78
timestamp 1688980957
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_90
timestamp 1688980957
transform 1 0 9384 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_112
timestamp 1688980957
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_116
timestamp 1688980957
transform 1 0 11776 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_169
timestamp 1688980957
transform 1 0 16652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1688980957
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_212
timestamp 1688980957
transform 1 0 20608 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_224
timestamp 1688980957
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_228
timestamp 1688980957
transform 1 0 22080 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_242
timestamp 1688980957
transform 1 0 23368 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_276
timestamp 1688980957
transform 1 0 26496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_284
timestamp 1688980957
transform 1 0 27232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_291
timestamp 1688980957
transform 1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_124
timestamp 1688980957
transform 1 0 12512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_142
timestamp 1688980957
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_216
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_233
timestamp 1688980957
transform 1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_254
timestamp 1688980957
transform 1 0 24472 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_266
timestamp 1688980957
transform 1 0 25576 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_323
timestamp 1688980957
transform 1 0 30820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_332
timestamp 1688980957
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_73
timestamp 1688980957
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_126
timestamp 1688980957
transform 1 0 12696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_157
timestamp 1688980957
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_167
timestamp 1688980957
transform 1 0 16468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_179
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_191
timestamp 1688980957
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_213
timestamp 1688980957
transform 1 0 20700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_225
timestamp 1688980957
transform 1 0 21804 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_244
timestamp 1688980957
transform 1 0 23552 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_264
timestamp 1688980957
transform 1 0 25392 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_276
timestamp 1688980957
transform 1 0 26496 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_288
timestamp 1688980957
transform 1 0 27600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_298
timestamp 1688980957
transform 1 0 28520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 1688980957
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_327
timestamp 1688980957
transform 1 0 31188 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_338
timestamp 1688980957
transform 1 0 32200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_350
timestamp 1688980957
transform 1 0 33304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_362
timestamp 1688980957
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_61
timestamp 1688980957
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_73
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_92
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_96
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_108
timestamp 1688980957
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_126
timestamp 1688980957
transform 1 0 12696 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_185
timestamp 1688980957
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_200
timestamp 1688980957
transform 1 0 19504 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_212
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_240
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_252
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_259
timestamp 1688980957
transform 1 0 24932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_271
timestamp 1688980957
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_289
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_296
timestamp 1688980957
transform 1 0 28336 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_308
timestamp 1688980957
transform 1 0 29440 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_319
timestamp 1688980957
transform 1 0 30452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_345
timestamp 1688980957
transform 1 0 32844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_357
timestamp 1688980957
transform 1 0 33948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_369
timestamp 1688980957
transform 1 0 35052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_381
timestamp 1688980957
transform 1 0 36156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_389
timestamp 1688980957
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_23
timestamp 1688980957
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_49
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_134
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_149
timestamp 1688980957
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_174
timestamp 1688980957
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1688980957
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_202
timestamp 1688980957
transform 1 0 19688 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_208
timestamp 1688980957
transform 1 0 20240 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_216
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_226
timestamp 1688980957
transform 1 0 21896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_246
timestamp 1688980957
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_270
timestamp 1688980957
transform 1 0 25944 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_282
timestamp 1688980957
transform 1 0 27048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_287
timestamp 1688980957
transform 1 0 27508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_304
timestamp 1688980957
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_315
timestamp 1688980957
transform 1 0 30084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_328
timestamp 1688980957
transform 1 0 31280 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_340
timestamp 1688980957
transform 1 0 32384 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_352
timestamp 1688980957
transform 1 0 33488 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_7
timestamp 1688980957
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_19
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_40
timestamp 1688980957
transform 1 0 4784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_50
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_60
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_72
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_84
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_91
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_182
timestamp 1688980957
transform 1 0 17848 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_194
timestamp 1688980957
transform 1 0 18952 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_219
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_238
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_246
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_271
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_289
timestamp 1688980957
transform 1 0 27692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_295
timestamp 1688980957
transform 1 0 28244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_321
timestamp 1688980957
transform 1 0 30636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_345
timestamp 1688980957
transform 1 0 32844 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_355
timestamp 1688980957
transform 1 0 33764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_367
timestamp 1688980957
transform 1 0 34868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_379
timestamp 1688980957
transform 1 0 35972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_35
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_43
timestamp 1688980957
transform 1 0 5060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_49
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_71
timestamp 1688980957
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_76
timestamp 1688980957
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_125
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_152
timestamp 1688980957
transform 1 0 15088 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_164
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_176
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_188
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1688980957
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_206
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_218
timestamp 1688980957
transform 1 0 21160 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_230
timestamp 1688980957
transform 1 0 22264 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_246
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_288
timestamp 1688980957
transform 1 0 27600 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_300
timestamp 1688980957
transform 1 0 28704 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_312
timestamp 1688980957
transform 1 0 29808 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_336
timestamp 1688980957
transform 1 0 32016 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_348
timestamp 1688980957
transform 1 0 33120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_360
timestamp 1688980957
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_11
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_14
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_24
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_32
timestamp 1688980957
transform 1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_40
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_80
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_97
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_127
timestamp 1688980957
transform 1 0 12788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_139
timestamp 1688980957
transform 1 0 13892 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_216
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_245
timestamp 1688980957
transform 1 0 23644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_266
timestamp 1688980957
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_286
timestamp 1688980957
transform 1 0 27416 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_294
timestamp 1688980957
transform 1 0 28152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_299
timestamp 1688980957
transform 1 0 28612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_304
timestamp 1688980957
transform 1 0 29072 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_312
timestamp 1688980957
transform 1 0 29808 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_318
timestamp 1688980957
transform 1 0 30360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_326
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_352
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_364
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_376
timestamp 1688980957
transform 1 0 35696 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_388
timestamp 1688980957
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_12
timestamp 1688980957
transform 1 0 2208 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_48
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_60
timestamp 1688980957
transform 1 0 6624 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_72
timestamp 1688980957
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1688980957
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_91
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_112
timestamp 1688980957
transform 1 0 11408 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_149
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_159
timestamp 1688980957
transform 1 0 15732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_171
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_175
timestamp 1688980957
transform 1 0 17204 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_186
timestamp 1688980957
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1688980957
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_243
timestamp 1688980957
transform 1 0 23460 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_248
timestamp 1688980957
transform 1 0 23920 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_261
timestamp 1688980957
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_278
timestamp 1688980957
transform 1 0 26680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_293
timestamp 1688980957
transform 1 0 28060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_302
timestamp 1688980957
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_314
timestamp 1688980957
transform 1 0 29992 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_326
timestamp 1688980957
transform 1 0 31096 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_340
timestamp 1688980957
transform 1 0 32384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_355
timestamp 1688980957
transform 1 0 33764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_31
timestamp 1688980957
transform 1 0 3956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_67
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_75
timestamp 1688980957
transform 1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_87
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_99
timestamp 1688980957
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_131
timestamp 1688980957
transform 1 0 13156 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_147
timestamp 1688980957
transform 1 0 14628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_159
timestamp 1688980957
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_190
timestamp 1688980957
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_198
timestamp 1688980957
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_211
timestamp 1688980957
transform 1 0 20516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_216
timestamp 1688980957
transform 1 0 20976 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_238
timestamp 1688980957
transform 1 0 23000 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_250
timestamp 1688980957
transform 1 0 24104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_265
timestamp 1688980957
transform 1 0 25484 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_276
timestamp 1688980957
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_289
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_301
timestamp 1688980957
transform 1 0 28796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_307
timestamp 1688980957
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_314
timestamp 1688980957
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_318
timestamp 1688980957
transform 1 0 30360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_348
timestamp 1688980957
transform 1 0 33120 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_360
timestamp 1688980957
transform 1 0 34224 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_372
timestamp 1688980957
transform 1 0 35328 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_384
timestamp 1688980957
transform 1 0 36432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_33
timestamp 1688980957
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_42
timestamp 1688980957
transform 1 0 4968 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_120
timestamp 1688980957
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_132
timestamp 1688980957
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_147
timestamp 1688980957
transform 1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_152
timestamp 1688980957
transform 1 0 15088 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_202
timestamp 1688980957
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_225
timestamp 1688980957
transform 1 0 21804 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_244
timestamp 1688980957
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_262
timestamp 1688980957
transform 1 0 25208 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_274
timestamp 1688980957
transform 1 0 26312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_286
timestamp 1688980957
transform 1 0 27416 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_306
timestamp 1688980957
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_313
timestamp 1688980957
transform 1 0 29900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_325
timestamp 1688980957
transform 1 0 31004 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_339
timestamp 1688980957
transform 1 0 32292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_351
timestamp 1688980957
transform 1 0 33396 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_372
timestamp 1688980957
transform 1 0 35328 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_384
timestamp 1688980957
transform 1 0 36432 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_396
timestamp 1688980957
transform 1 0 37536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_400
timestamp 1688980957
transform 1 0 37904 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_47
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_60
timestamp 1688980957
transform 1 0 6624 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_72
timestamp 1688980957
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_104
timestamp 1688980957
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_119
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_127
timestamp 1688980957
transform 1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_182
timestamp 1688980957
transform 1 0 17848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_199
timestamp 1688980957
transform 1 0 19412 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_211
timestamp 1688980957
transform 1 0 20516 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1688980957
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_238
timestamp 1688980957
transform 1 0 23000 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_247
timestamp 1688980957
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_259
timestamp 1688980957
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_271
timestamp 1688980957
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_290
timestamp 1688980957
transform 1 0 27784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_296
timestamp 1688980957
transform 1 0 28336 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_307
timestamp 1688980957
transform 1 0 29348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_319
timestamp 1688980957
transform 1 0 30452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_325
timestamp 1688980957
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_333
timestamp 1688980957
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_351
timestamp 1688980957
transform 1 0 33396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_359
timestamp 1688980957
transform 1 0 34132 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_368
timestamp 1688980957
transform 1 0 34960 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_380
timestamp 1688980957
transform 1 0 36064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_384
timestamp 1688980957
transform 1 0 36432 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1688980957
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_7
timestamp 1688980957
transform 1 0 1748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_18
timestamp 1688980957
transform 1 0 2760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_22
timestamp 1688980957
transform 1 0 3128 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1688980957
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_59
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_69
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_98
timestamp 1688980957
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_105
timestamp 1688980957
transform 1 0 10764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_144
timestamp 1688980957
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_158
timestamp 1688980957
transform 1 0 15640 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_170
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_212
timestamp 1688980957
transform 1 0 20608 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_224
timestamp 1688980957
transform 1 0 21712 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_236
timestamp 1688980957
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 1688980957
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_256
timestamp 1688980957
transform 1 0 24656 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_270
timestamp 1688980957
transform 1 0 25944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_297
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 1688980957
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_315
timestamp 1688980957
transform 1 0 30084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_327
timestamp 1688980957
transform 1 0 31188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_350
timestamp 1688980957
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_362
timestamp 1688980957
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_23
timestamp 1688980957
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_35
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_47
timestamp 1688980957
transform 1 0 5428 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_117
timestamp 1688980957
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_127
timestamp 1688980957
transform 1 0 12788 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_151
timestamp 1688980957
transform 1 0 14996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_155
timestamp 1688980957
transform 1 0 15364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_159
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_185
timestamp 1688980957
transform 1 0 18124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1688980957
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_233
timestamp 1688980957
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_239
timestamp 1688980957
transform 1 0 23092 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_247
timestamp 1688980957
transform 1 0 23828 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_256
timestamp 1688980957
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_269
timestamp 1688980957
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_277
timestamp 1688980957
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_286
timestamp 1688980957
transform 1 0 27416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_298
timestamp 1688980957
transform 1 0 28520 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_308
timestamp 1688980957
transform 1 0 29440 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_358
timestamp 1688980957
transform 1 0 34040 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_370
timestamp 1688980957
transform 1 0 35144 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_382
timestamp 1688980957
transform 1 0 36248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_390
timestamp 1688980957
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_10
timestamp 1688980957
transform 1 0 2024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_21
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_67
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_98
timestamp 1688980957
transform 1 0 10120 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_122
timestamp 1688980957
transform 1 0 12328 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_131
timestamp 1688980957
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_149
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_159
timestamp 1688980957
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1688980957
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_207
timestamp 1688980957
transform 1 0 20148 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_215
timestamp 1688980957
transform 1 0 20884 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_228
timestamp 1688980957
transform 1 0 22080 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_264
timestamp 1688980957
transform 1 0 25392 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_272
timestamp 1688980957
transform 1 0 26128 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_282
timestamp 1688980957
transform 1 0 27048 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_294
timestamp 1688980957
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_298
timestamp 1688980957
transform 1 0 28520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_317
timestamp 1688980957
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_323
timestamp 1688980957
transform 1 0 30820 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_335
timestamp 1688980957
transform 1 0 31924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_347
timestamp 1688980957
transform 1 0 33028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_359
timestamp 1688980957
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_22
timestamp 1688980957
transform 1 0 3128 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_47
timestamp 1688980957
transform 1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1688980957
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_66
timestamp 1688980957
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_78
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_92
timestamp 1688980957
transform 1 0 9568 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_136
timestamp 1688980957
transform 1 0 13616 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_148
timestamp 1688980957
transform 1 0 14720 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_160
timestamp 1688980957
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_203
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_207
timestamp 1688980957
transform 1 0 20148 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 1688980957
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_277
timestamp 1688980957
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_289
timestamp 1688980957
transform 1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_297
timestamp 1688980957
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_309
timestamp 1688980957
transform 1 0 29532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_327
timestamp 1688980957
transform 1 0 31188 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_342
timestamp 1688980957
transform 1 0 32568 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_358
timestamp 1688980957
transform 1 0 34040 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_370
timestamp 1688980957
transform 1 0 35144 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_382
timestamp 1688980957
transform 1 0 36248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_390
timestamp 1688980957
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_12
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 1688980957
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_33
timestamp 1688980957
transform 1 0 4140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_80
timestamp 1688980957
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_99
timestamp 1688980957
transform 1 0 10212 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_111
timestamp 1688980957
transform 1 0 11316 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_149
timestamp 1688980957
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_157
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_169
timestamp 1688980957
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_180
timestamp 1688980957
transform 1 0 17664 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_205
timestamp 1688980957
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_236
timestamp 1688980957
transform 1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_246
timestamp 1688980957
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_263
timestamp 1688980957
transform 1 0 25300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_269
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_287
timestamp 1688980957
transform 1 0 27508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_303
timestamp 1688980957
transform 1 0 28980 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_317
timestamp 1688980957
transform 1 0 30268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_328
timestamp 1688980957
transform 1 0 31280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_338
timestamp 1688980957
transform 1 0 32200 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_342
timestamp 1688980957
transform 1 0 32568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_361
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_23
timestamp 1688980957
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_41
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_48
timestamp 1688980957
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_66
timestamp 1688980957
transform 1 0 7176 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_92
timestamp 1688980957
transform 1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_100
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_126
timestamp 1688980957
transform 1 0 12696 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_146
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_153
timestamp 1688980957
transform 1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_158
timestamp 1688980957
transform 1 0 15640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_162
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1688980957
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_173
timestamp 1688980957
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_194
timestamp 1688980957
transform 1 0 18952 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_206
timestamp 1688980957
transform 1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_210
timestamp 1688980957
transform 1 0 20424 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_231
timestamp 1688980957
transform 1 0 22356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_270
timestamp 1688980957
transform 1 0 25944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_276
timestamp 1688980957
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_284
timestamp 1688980957
transform 1 0 27232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_296
timestamp 1688980957
transform 1 0 28336 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_300
timestamp 1688980957
transform 1 0 28704 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_312
timestamp 1688980957
transform 1 0 29808 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_320
timestamp 1688980957
transform 1 0 30544 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_328
timestamp 1688980957
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_345
timestamp 1688980957
transform 1 0 32844 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_355
timestamp 1688980957
transform 1 0 33764 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_367
timestamp 1688980957
transform 1 0 34868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_379
timestamp 1688980957
transform 1 0 35972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_33
timestamp 1688980957
transform 1 0 4140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_37
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_62
timestamp 1688980957
transform 1 0 6808 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_150
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_173
timestamp 1688980957
transform 1 0 17020 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_208
timestamp 1688980957
transform 1 0 20240 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_247
timestamp 1688980957
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_260
timestamp 1688980957
transform 1 0 25024 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_272
timestamp 1688980957
transform 1 0 26128 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_284
timestamp 1688980957
transform 1 0 27232 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_291
timestamp 1688980957
transform 1 0 27876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_300
timestamp 1688980957
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_317
timestamp 1688980957
transform 1 0 30268 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_336
timestamp 1688980957
transform 1 0 32016 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_353
timestamp 1688980957
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_361
timestamp 1688980957
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_12
timestamp 1688980957
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_25
timestamp 1688980957
transform 1 0 3404 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_33
timestamp 1688980957
transform 1 0 4140 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_40
timestamp 1688980957
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1688980957
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_78
timestamp 1688980957
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_90
timestamp 1688980957
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_100
timestamp 1688980957
transform 1 0 10304 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_122
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_128
timestamp 1688980957
transform 1 0 12880 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_157
timestamp 1688980957
transform 1 0 15548 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_165
timestamp 1688980957
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_184
timestamp 1688980957
transform 1 0 18032 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_204
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_209
timestamp 1688980957
transform 1 0 20332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_250
timestamp 1688980957
transform 1 0 24104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_254
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_260
timestamp 1688980957
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_264
timestamp 1688980957
transform 1 0 25392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_326
timestamp 1688980957
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_334
timestamp 1688980957
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_345
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_356
timestamp 1688980957
transform 1 0 33856 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_368
timestamp 1688980957
transform 1 0 34960 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_380
timestamp 1688980957
transform 1 0 36064 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_23
timestamp 1688980957
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_38
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_50
timestamp 1688980957
transform 1 0 5704 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_62
timestamp 1688980957
transform 1 0 6808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_74
timestamp 1688980957
transform 1 0 7912 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_80
timestamp 1688980957
transform 1 0 8464 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_128
timestamp 1688980957
transform 1 0 12880 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_173
timestamp 1688980957
transform 1 0 17020 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_179
timestamp 1688980957
transform 1 0 17572 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_191
timestamp 1688980957
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_219
timestamp 1688980957
transform 1 0 21252 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_244
timestamp 1688980957
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_275
timestamp 1688980957
transform 1 0 26404 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_283
timestamp 1688980957
transform 1 0 27140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_292
timestamp 1688980957
transform 1 0 27968 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_298
timestamp 1688980957
transform 1 0 28520 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_302
timestamp 1688980957
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_316
timestamp 1688980957
transform 1 0 30176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_325
timestamp 1688980957
transform 1 0 31004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_332
timestamp 1688980957
transform 1 0 31648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_342
timestamp 1688980957
transform 1 0 32568 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_352
timestamp 1688980957
transform 1 0 33488 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_21
timestamp 1688980957
transform 1 0 3036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_29
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_41
timestamp 1688980957
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_74
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_84
timestamp 1688980957
transform 1 0 8832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_94
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_106
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_134
timestamp 1688980957
transform 1 0 13432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_138
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_159
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_186
timestamp 1688980957
transform 1 0 18216 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_192
timestamp 1688980957
transform 1 0 18768 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_215
timestamp 1688980957
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_261
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_313
timestamp 1688980957
transform 1 0 29900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_324
timestamp 1688980957
transform 1 0 30912 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_362
timestamp 1688980957
transform 1 0 34408 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_374
timestamp 1688980957
transform 1 0 35512 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_386
timestamp 1688980957
transform 1 0 36616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_12
timestamp 1688980957
transform 1 0 2208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_24
timestamp 1688980957
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_44
timestamp 1688980957
transform 1 0 5152 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_50
timestamp 1688980957
transform 1 0 5704 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_60
timestamp 1688980957
transform 1 0 6624 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_92
timestamp 1688980957
transform 1 0 9568 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_104
timestamp 1688980957
transform 1 0 10672 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_116
timestamp 1688980957
transform 1 0 11776 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_150
timestamp 1688980957
transform 1 0 14904 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_162
timestamp 1688980957
transform 1 0 16008 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_174
timestamp 1688980957
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_178
timestamp 1688980957
transform 1 0 17480 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1688980957
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_219
timestamp 1688980957
transform 1 0 21252 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_229
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_240
timestamp 1688980957
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_331
timestamp 1688980957
transform 1 0 31556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_343
timestamp 1688980957
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_355
timestamp 1688980957
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_372
timestamp 1688980957
transform 1 0 35328 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_384
timestamp 1688980957
transform 1 0 36432 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_396
timestamp 1688980957
transform 1 0 37536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_400
timestamp 1688980957
transform 1 0 37904 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_23
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_29
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_42
timestamp 1688980957
transform 1 0 4968 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_87
timestamp 1688980957
transform 1 0 9108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_96
timestamp 1688980957
transform 1 0 9936 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_104
timestamp 1688980957
transform 1 0 10672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_122
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_135
timestamp 1688980957
transform 1 0 13524 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_147
timestamp 1688980957
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_154
timestamp 1688980957
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_185
timestamp 1688980957
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_194
timestamp 1688980957
transform 1 0 18952 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_200
timestamp 1688980957
transform 1 0 19504 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_252
timestamp 1688980957
transform 1 0 24288 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_264
timestamp 1688980957
transform 1 0 25392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_276
timestamp 1688980957
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_289
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_309
timestamp 1688980957
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_321
timestamp 1688980957
transform 1 0 30636 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_342
timestamp 1688980957
transform 1 0 32568 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_354
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_375
timestamp 1688980957
transform 1 0 35604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_387
timestamp 1688980957
transform 1 0 36708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_24
timestamp 1688980957
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_40
timestamp 1688980957
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_44
timestamp 1688980957
transform 1 0 5152 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_70
timestamp 1688980957
transform 1 0 7544 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_80
timestamp 1688980957
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_99
timestamp 1688980957
transform 1 0 10212 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_154
timestamp 1688980957
transform 1 0 15272 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_161
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_171
timestamp 1688980957
transform 1 0 16836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_183
timestamp 1688980957
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_188
timestamp 1688980957
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_203
timestamp 1688980957
transform 1 0 19780 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_217
timestamp 1688980957
transform 1 0 21068 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_229
timestamp 1688980957
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_242
timestamp 1688980957
transform 1 0 23368 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_260
timestamp 1688980957
transform 1 0 25024 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_283
timestamp 1688980957
transform 1 0 27140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_304
timestamp 1688980957
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_320
timestamp 1688980957
transform 1 0 30544 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_328
timestamp 1688980957
transform 1 0 31280 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_336
timestamp 1688980957
transform 1 0 32016 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_353
timestamp 1688980957
transform 1 0 33580 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_10
timestamp 1688980957
transform 1 0 2024 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_14
timestamp 1688980957
transform 1 0 2392 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_22
timestamp 1688980957
transform 1 0 3128 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_28
timestamp 1688980957
transform 1 0 3680 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_40
timestamp 1688980957
transform 1 0 4784 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 1688980957
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_71
timestamp 1688980957
transform 1 0 7636 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_103
timestamp 1688980957
transform 1 0 10580 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_123
timestamp 1688980957
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_135
timestamp 1688980957
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_147
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_155
timestamp 1688980957
transform 1 0 15364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_163
timestamp 1688980957
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_176
timestamp 1688980957
transform 1 0 17296 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_182
timestamp 1688980957
transform 1 0 17848 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_192
timestamp 1688980957
transform 1 0 18768 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_201
timestamp 1688980957
transform 1 0 19596 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_212
timestamp 1688980957
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_303
timestamp 1688980957
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_315
timestamp 1688980957
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_327
timestamp 1688980957
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_348
timestamp 1688980957
transform 1 0 33120 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_360
timestamp 1688980957
transform 1 0 34224 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_370
timestamp 1688980957
transform 1 0 35144 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_382
timestamp 1688980957
transform 1 0 36248 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_390
timestamp 1688980957
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_19
timestamp 1688980957
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_37
timestamp 1688980957
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_43
timestamp 1688980957
transform 1 0 5060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_56
timestamp 1688980957
transform 1 0 6256 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_62
timestamp 1688980957
transform 1 0 6808 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_182
timestamp 1688980957
transform 1 0 17848 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_207
timestamp 1688980957
transform 1 0 20148 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_213
timestamp 1688980957
transform 1 0 20700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_225
timestamp 1688980957
transform 1 0 21804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_261
timestamp 1688980957
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_279
timestamp 1688980957
transform 1 0 26772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_291
timestamp 1688980957
transform 1 0 27876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_302
timestamp 1688980957
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_338
timestamp 1688980957
transform 1 0 32200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_343
timestamp 1688980957
transform 1 0 32660 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_348
timestamp 1688980957
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_360
timestamp 1688980957
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_378
timestamp 1688980957
transform 1 0 35880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_390
timestamp 1688980957
transform 1 0 36984 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_398
timestamp 1688980957
transform 1 0 37720 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1688980957
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_64
timestamp 1688980957
transform 1 0 6992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_68
timestamp 1688980957
transform 1 0 7360 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_72
timestamp 1688980957
transform 1 0 7728 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_84
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_90
timestamp 1688980957
transform 1 0 9384 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_98
timestamp 1688980957
transform 1 0 10120 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_106
timestamp 1688980957
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_174
timestamp 1688980957
transform 1 0 17112 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_182
timestamp 1688980957
transform 1 0 17848 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_209
timestamp 1688980957
transform 1 0 20332 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_242
timestamp 1688980957
transform 1 0 23368 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_256
timestamp 1688980957
transform 1 0 24656 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_264
timestamp 1688980957
transform 1 0 25392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_270
timestamp 1688980957
transform 1 0 25944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 1688980957
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_288
timestamp 1688980957
transform 1 0 27600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_292
timestamp 1688980957
transform 1 0 27968 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_307
timestamp 1688980957
transform 1 0 29348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_334
timestamp 1688980957
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_347
timestamp 1688980957
transform 1 0 33028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_355
timestamp 1688980957
transform 1 0 33764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_359
timestamp 1688980957
transform 1 0 34132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_371
timestamp 1688980957
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_383
timestamp 1688980957
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1688980957
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_34
timestamp 1688980957
transform 1 0 4232 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_46
timestamp 1688980957
transform 1 0 5336 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_54
timestamp 1688980957
transform 1 0 6072 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_66
timestamp 1688980957
transform 1 0 7176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_71
timestamp 1688980957
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_128
timestamp 1688980957
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_146
timestamp 1688980957
transform 1 0 14536 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_166
timestamp 1688980957
transform 1 0 16376 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_174
timestamp 1688980957
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_184
timestamp 1688980957
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_205
timestamp 1688980957
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_215
timestamp 1688980957
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_223
timestamp 1688980957
transform 1 0 21620 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1688980957
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_260
timestamp 1688980957
transform 1 0 25024 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_264
timestamp 1688980957
transform 1 0 25392 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_272
timestamp 1688980957
transform 1 0 26128 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_276
timestamp 1688980957
transform 1 0 26496 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_285
timestamp 1688980957
transform 1 0 27324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_299
timestamp 1688980957
transform 1 0 28612 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_319
timestamp 1688980957
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_331
timestamp 1688980957
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_343
timestamp 1688980957
transform 1 0 32660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_347
timestamp 1688980957
transform 1 0 33028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_351
timestamp 1688980957
transform 1 0 33396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_373
timestamp 1688980957
transform 1 0 35420 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_385
timestamp 1688980957
transform 1 0 36524 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_397
timestamp 1688980957
transform 1 0 37628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_9
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_38
timestamp 1688980957
transform 1 0 4600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_50
timestamp 1688980957
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_61
timestamp 1688980957
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_83
timestamp 1688980957
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_131
timestamp 1688980957
transform 1 0 13156 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_156
timestamp 1688980957
transform 1 0 15456 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_174
timestamp 1688980957
transform 1 0 17112 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_186
timestamp 1688980957
transform 1 0 18216 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_198
timestamp 1688980957
transform 1 0 19320 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_210
timestamp 1688980957
transform 1 0 20424 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 1688980957
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_244
timestamp 1688980957
transform 1 0 23552 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_253
timestamp 1688980957
transform 1 0 24380 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_268
timestamp 1688980957
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_306
timestamp 1688980957
transform 1 0 29256 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_314
timestamp 1688980957
transform 1 0 29992 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_326
timestamp 1688980957
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1688980957
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_365
timestamp 1688980957
transform 1 0 34684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_383
timestamp 1688980957
transform 1 0 36340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_23
timestamp 1688980957
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_37
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_91
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_106
timestamp 1688980957
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_118
timestamp 1688980957
transform 1 0 11960 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_129
timestamp 1688980957
transform 1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1688980957
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_156
timestamp 1688980957
transform 1 0 15456 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_164
timestamp 1688980957
transform 1 0 16192 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_171
timestamp 1688980957
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_229
timestamp 1688980957
transform 1 0 22172 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_241
timestamp 1688980957
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_297
timestamp 1688980957
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 1688980957
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_317
timestamp 1688980957
transform 1 0 30268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_329
timestamp 1688980957
transform 1 0 31372 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_344
timestamp 1688980957
transform 1 0 32752 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_356
timestamp 1688980957
transform 1 0 33856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_372
timestamp 1688980957
transform 1 0 35328 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1688980957
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_389
timestamp 1688980957
transform 1 0 36892 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_11
timestamp 1688980957
transform 1 0 2116 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_24
timestamp 1688980957
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_36
timestamp 1688980957
transform 1 0 4416 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_52
timestamp 1688980957
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_85
timestamp 1688980957
transform 1 0 8924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_100
timestamp 1688980957
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_136
timestamp 1688980957
transform 1 0 13616 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_144
timestamp 1688980957
transform 1 0 14352 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_152
timestamp 1688980957
transform 1 0 15088 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_160
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_172
timestamp 1688980957
transform 1 0 16928 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_213
timestamp 1688980957
transform 1 0 20700 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_221
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_231
timestamp 1688980957
transform 1 0 22356 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_242
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_254
timestamp 1688980957
transform 1 0 24472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_263
timestamp 1688980957
transform 1 0 25300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_274
timestamp 1688980957
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_292
timestamp 1688980957
transform 1 0 27968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_300
timestamp 1688980957
transform 1 0 28704 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_306
timestamp 1688980957
transform 1 0 29256 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_318
timestamp 1688980957
transform 1 0 30360 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_326
timestamp 1688980957
transform 1 0 31096 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_347
timestamp 1688980957
transform 1 0 33028 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_355
timestamp 1688980957
transform 1 0 33764 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_364
timestamp 1688980957
transform 1 0 34592 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_368
timestamp 1688980957
transform 1 0 34960 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_380
timestamp 1688980957
transform 1 0 36064 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_36
timestamp 1688980957
transform 1 0 4416 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_43
timestamp 1688980957
transform 1 0 5060 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_58
timestamp 1688980957
transform 1 0 6440 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_90
timestamp 1688980957
transform 1 0 9384 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_102
timestamp 1688980957
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_115
timestamp 1688980957
transform 1 0 11684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_129
timestamp 1688980957
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1688980957
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_183
timestamp 1688980957
transform 1 0 17940 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_226
timestamp 1688980957
transform 1 0 21896 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_235
timestamp 1688980957
transform 1 0 22724 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_247
timestamp 1688980957
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_268
timestamp 1688980957
transform 1 0 25760 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_285
timestamp 1688980957
transform 1 0 27324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_313
timestamp 1688980957
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_323
timestamp 1688980957
transform 1 0 30820 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_380
timestamp 1688980957
transform 1 0 36064 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_392
timestamp 1688980957
transform 1 0 37168 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_400
timestamp 1688980957
transform 1 0 37904 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_19
timestamp 1688980957
transform 1 0 2852 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_45
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_49
timestamp 1688980957
transform 1 0 5612 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_74
timestamp 1688980957
transform 1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_80
timestamp 1688980957
transform 1 0 8464 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_92
timestamp 1688980957
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_96
timestamp 1688980957
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_106
timestamp 1688980957
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_122
timestamp 1688980957
transform 1 0 12328 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_134
timestamp 1688980957
transform 1 0 13432 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_146
timestamp 1688980957
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_155
timestamp 1688980957
transform 1 0 15364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_183
timestamp 1688980957
transform 1 0 17940 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_199
timestamp 1688980957
transform 1 0 19412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_234
timestamp 1688980957
transform 1 0 22632 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_246
timestamp 1688980957
transform 1 0 23736 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_258
timestamp 1688980957
transform 1 0 24840 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_270
timestamp 1688980957
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_278
timestamp 1688980957
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_288
timestamp 1688980957
transform 1 0 27600 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_309
timestamp 1688980957
transform 1 0 29532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_321
timestamp 1688980957
transform 1 0 30636 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_344
timestamp 1688980957
transform 1 0 32752 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_356
timestamp 1688980957
transform 1 0 33856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_366
timestamp 1688980957
transform 1 0 34776 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_380
timestamp 1688980957
transform 1 0 36064 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_10
timestamp 1688980957
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_22
timestamp 1688980957
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_37
timestamp 1688980957
transform 1 0 4508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_69
timestamp 1688980957
transform 1 0 7452 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_90
timestamp 1688980957
transform 1 0 9384 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_118
timestamp 1688980957
transform 1 0 11960 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_130
timestamp 1688980957
transform 1 0 13064 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_156
timestamp 1688980957
transform 1 0 15456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_206
timestamp 1688980957
transform 1 0 20056 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_218
timestamp 1688980957
transform 1 0 21160 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1688980957
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_259
timestamp 1688980957
transform 1 0 24932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_270
timestamp 1688980957
transform 1 0 25944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_278
timestamp 1688980957
transform 1 0 26680 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_287
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_299
timestamp 1688980957
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_336
timestamp 1688980957
transform 1 0 32016 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_348
timestamp 1688980957
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_360
timestamp 1688980957
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_385
timestamp 1688980957
transform 1 0 36524 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_393
timestamp 1688980957
transform 1 0 37260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_397
timestamp 1688980957
transform 1 0 37628 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_23
timestamp 1688980957
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_35
timestamp 1688980957
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_47
timestamp 1688980957
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_75
timestamp 1688980957
transform 1 0 8004 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_87
timestamp 1688980957
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_99
timestamp 1688980957
transform 1 0 10212 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_103
timestamp 1688980957
transform 1 0 10580 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_107
timestamp 1688980957
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_133
timestamp 1688980957
transform 1 0 13340 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_143
timestamp 1688980957
transform 1 0 14260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_155
timestamp 1688980957
transform 1 0 15364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_159
timestamp 1688980957
transform 1 0 15732 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_201
timestamp 1688980957
transform 1 0 19596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_213
timestamp 1688980957
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_229
timestamp 1688980957
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_272
timestamp 1688980957
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_288
timestamp 1688980957
transform 1 0 27600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_292
timestamp 1688980957
transform 1 0 27968 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_314
timestamp 1688980957
transform 1 0 29992 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_326
timestamp 1688980957
transform 1 0 31096 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_342
timestamp 1688980957
transform 1 0 32568 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_354
timestamp 1688980957
transform 1 0 33672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_362
timestamp 1688980957
transform 1 0 34408 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 1688980957
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 1688980957
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_34
timestamp 1688980957
transform 1 0 4232 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_45
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_57
timestamp 1688980957
transform 1 0 6348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_78
timestamp 1688980957
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_119
timestamp 1688980957
transform 1 0 12052 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_123
timestamp 1688980957
transform 1 0 12420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_157
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_176
timestamp 1688980957
transform 1 0 17296 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_193
timestamp 1688980957
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_223
timestamp 1688980957
transform 1 0 21620 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_244
timestamp 1688980957
transform 1 0 23552 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_248
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_263
timestamp 1688980957
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_267
timestamp 1688980957
transform 1 0 25668 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_276
timestamp 1688980957
transform 1 0 26496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_285
timestamp 1688980957
transform 1 0 27324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_304
timestamp 1688980957
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_313
timestamp 1688980957
transform 1 0 29900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_351
timestamp 1688980957
transform 1 0 33396 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_378
timestamp 1688980957
transform 1 0 35880 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_390
timestamp 1688980957
transform 1 0 36984 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_398
timestamp 1688980957
transform 1 0 37720 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_9
timestamp 1688980957
transform 1 0 1932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_23
timestamp 1688980957
transform 1 0 3220 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_45
timestamp 1688980957
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_103
timestamp 1688980957
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_153
timestamp 1688980957
transform 1 0 15180 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_187
timestamp 1688980957
transform 1 0 18308 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_202
timestamp 1688980957
transform 1 0 19688 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_208
timestamp 1688980957
transform 1 0 20240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_236
timestamp 1688980957
transform 1 0 22816 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_248
timestamp 1688980957
transform 1 0 23920 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_260
timestamp 1688980957
transform 1 0 25024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_264
timestamp 1688980957
transform 1 0 25392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_272
timestamp 1688980957
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_300
timestamp 1688980957
transform 1 0 28704 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_304
timestamp 1688980957
transform 1 0 29072 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_311
timestamp 1688980957
transform 1 0 29716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_323
timestamp 1688980957
transform 1 0 30820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_346
timestamp 1688980957
transform 1 0 32936 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_358
timestamp 1688980957
transform 1 0 34040 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_369
timestamp 1688980957
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_381
timestamp 1688980957
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_389
timestamp 1688980957
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_78
timestamp 1688980957
transform 1 0 8280 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_82
timestamp 1688980957
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_89
timestamp 1688980957
transform 1 0 9292 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_123
timestamp 1688980957
transform 1 0 12420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_157
timestamp 1688980957
transform 1 0 15548 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_183
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1688980957
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_223
timestamp 1688980957
transform 1 0 21620 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_231
timestamp 1688980957
transform 1 0 22356 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_239
timestamp 1688980957
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_262
timestamp 1688980957
transform 1 0 25208 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_278
timestamp 1688980957
transform 1 0 26680 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_290
timestamp 1688980957
transform 1 0 27784 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_305
timestamp 1688980957
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_361
timestamp 1688980957
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_54
timestamp 1688980957
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_67
timestamp 1688980957
transform 1 0 7268 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_79
timestamp 1688980957
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_91
timestamp 1688980957
transform 1 0 9476 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_102
timestamp 1688980957
transform 1 0 10488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_110
timestamp 1688980957
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_120
timestamp 1688980957
transform 1 0 12144 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_128
timestamp 1688980957
transform 1 0 12880 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_160
timestamp 1688980957
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_185
timestamp 1688980957
transform 1 0 18124 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_191
timestamp 1688980957
transform 1 0 18676 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_203
timestamp 1688980957
transform 1 0 19780 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_209
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_216
timestamp 1688980957
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_257
timestamp 1688980957
transform 1 0 24748 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_265
timestamp 1688980957
transform 1 0 25484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_275
timestamp 1688980957
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_286
timestamp 1688980957
transform 1 0 27416 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_296
timestamp 1688980957
transform 1 0 28336 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_300
timestamp 1688980957
transform 1 0 28704 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_327
timestamp 1688980957
transform 1 0 31188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_346
timestamp 1688980957
transform 1 0 32936 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_384
timestamp 1688980957
transform 1 0 36432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_37
timestamp 1688980957
transform 1 0 4508 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_66
timestamp 1688980957
transform 1 0 7176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_78
timestamp 1688980957
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_88
timestamp 1688980957
transform 1 0 9200 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_119
timestamp 1688980957
transform 1 0 12052 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_131
timestamp 1688980957
transform 1 0 13156 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_154
timestamp 1688980957
transform 1 0 15272 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_162
timestamp 1688980957
transform 1 0 16008 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_171
timestamp 1688980957
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_186
timestamp 1688980957
transform 1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1688980957
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_213
timestamp 1688980957
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_226
timestamp 1688980957
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_238
timestamp 1688980957
transform 1 0 23000 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_246
timestamp 1688980957
transform 1 0 23736 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_303
timestamp 1688980957
transform 1 0 28980 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_319
timestamp 1688980957
transform 1 0 30452 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_328
timestamp 1688980957
transform 1 0 31280 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_359
timestamp 1688980957
transform 1 0 34132 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_388
timestamp 1688980957
transform 1 0 36800 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_400
timestamp 1688980957
transform 1 0 37904 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_47
timestamp 1688980957
transform 1 0 5428 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_53
timestamp 1688980957
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_75
timestamp 1688980957
transform 1 0 8004 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_108
timestamp 1688980957
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_122
timestamp 1688980957
transform 1 0 12328 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_136
timestamp 1688980957
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_162
timestamp 1688980957
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_180
timestamp 1688980957
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_184
timestamp 1688980957
transform 1 0 18032 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_199
timestamp 1688980957
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_211
timestamp 1688980957
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_265
timestamp 1688980957
transform 1 0 25484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_276
timestamp 1688980957
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_285
timestamp 1688980957
transform 1 0 27324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_289
timestamp 1688980957
transform 1 0 27692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_297
timestamp 1688980957
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_307
timestamp 1688980957
transform 1 0 29348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_319
timestamp 1688980957
transform 1 0 30452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_331
timestamp 1688980957
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_357
timestamp 1688980957
transform 1 0 33948 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_362
timestamp 1688980957
transform 1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_369
timestamp 1688980957
transform 1 0 35052 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_381
timestamp 1688980957
transform 1 0 36156 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_389
timestamp 1688980957
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_42
timestamp 1688980957
transform 1 0 4968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_46
timestamp 1688980957
transform 1 0 5336 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_56
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_69
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_113
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_123
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_129
timestamp 1688980957
transform 1 0 12972 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_145
timestamp 1688980957
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_166
timestamp 1688980957
transform 1 0 16376 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_206
timestamp 1688980957
transform 1 0 20056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_210
timestamp 1688980957
transform 1 0 20424 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_218
timestamp 1688980957
transform 1 0 21160 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_234
timestamp 1688980957
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_246
timestamp 1688980957
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_292
timestamp 1688980957
transform 1 0 27968 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_304
timestamp 1688980957
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_317
timestamp 1688980957
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_330
timestamp 1688980957
transform 1 0 31464 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_342
timestamp 1688980957
transform 1 0 32568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_350
timestamp 1688980957
transform 1 0 33304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_355
timestamp 1688980957
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_54
timestamp 1688980957
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_82
timestamp 1688980957
transform 1 0 8648 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_94
timestamp 1688980957
transform 1 0 9752 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_106
timestamp 1688980957
transform 1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_133
timestamp 1688980957
transform 1 0 13340 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_141
timestamp 1688980957
transform 1 0 14076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_158
timestamp 1688980957
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_166
timestamp 1688980957
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_173
timestamp 1688980957
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_232
timestamp 1688980957
transform 1 0 22448 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_250
timestamp 1688980957
transform 1 0 24104 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_262
timestamp 1688980957
transform 1 0 25208 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_276
timestamp 1688980957
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_285
timestamp 1688980957
transform 1 0 27324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_297
timestamp 1688980957
transform 1 0 28428 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_309
timestamp 1688980957
transform 1 0 29532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_324
timestamp 1688980957
transform 1 0 30912 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_332
timestamp 1688980957
transform 1 0 31648 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_346
timestamp 1688980957
transform 1 0 32936 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_379
timestamp 1688980957
transform 1 0 35972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_10
timestamp 1688980957
transform 1 0 2024 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_22
timestamp 1688980957
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_33
timestamp 1688980957
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_37
timestamp 1688980957
transform 1 0 4508 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_45
timestamp 1688980957
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_57
timestamp 1688980957
transform 1 0 6348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_61
timestamp 1688980957
transform 1 0 6716 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_94
timestamp 1688980957
transform 1 0 9752 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_111
timestamp 1688980957
transform 1 0 11316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_117
timestamp 1688980957
transform 1 0 11868 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_125
timestamp 1688980957
transform 1 0 12604 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_171
timestamp 1688980957
transform 1 0 16836 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_188
timestamp 1688980957
transform 1 0 18400 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_205
timestamp 1688980957
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_213
timestamp 1688980957
transform 1 0 20700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_225
timestamp 1688980957
transform 1 0 21804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_243
timestamp 1688980957
transform 1 0 23460 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_261
timestamp 1688980957
transform 1 0 25116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_278
timestamp 1688980957
transform 1 0 26680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_306
timestamp 1688980957
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_351
timestamp 1688980957
transform 1 0 33396 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_362
timestamp 1688980957
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_368
timestamp 1688980957
transform 1 0 34960 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_380
timestamp 1688980957
transform 1 0 36064 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_392
timestamp 1688980957
transform 1 0 37168 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_400
timestamp 1688980957
transform 1 0 37904 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_66
timestamp 1688980957
transform 1 0 7176 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_90
timestamp 1688980957
transform 1 0 9384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_126
timestamp 1688980957
transform 1 0 12696 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_134
timestamp 1688980957
transform 1 0 13432 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_146
timestamp 1688980957
transform 1 0 14536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_158
timestamp 1688980957
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1688980957
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_197
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_209
timestamp 1688980957
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1688980957
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_246
timestamp 1688980957
transform 1 0 23736 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_258
timestamp 1688980957
transform 1 0 24840 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_268
timestamp 1688980957
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_284
timestamp 1688980957
transform 1 0 27232 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_296
timestamp 1688980957
transform 1 0 28336 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_319
timestamp 1688980957
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_334
timestamp 1688980957
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_346
timestamp 1688980957
transform 1 0 32936 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_358
timestamp 1688980957
transform 1 0 34040 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_384
timestamp 1688980957
transform 1 0 36432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_35
timestamp 1688980957
transform 1 0 4324 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_39
timestamp 1688980957
transform 1 0 4692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_47
timestamp 1688980957
transform 1 0 5428 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_58
timestamp 1688980957
transform 1 0 6440 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_73
timestamp 1688980957
transform 1 0 7820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1688980957
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_91
timestamp 1688980957
transform 1 0 9476 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_95
timestamp 1688980957
transform 1 0 9844 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_107
timestamp 1688980957
transform 1 0 10948 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_119
timestamp 1688980957
transform 1 0 12052 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_125
timestamp 1688980957
transform 1 0 12604 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_155
timestamp 1688980957
transform 1 0 15364 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_172
timestamp 1688980957
transform 1 0 16928 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_180
timestamp 1688980957
transform 1 0 17664 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_191
timestamp 1688980957
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_203
timestamp 1688980957
transform 1 0 19780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_216
timestamp 1688980957
transform 1 0 20976 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_228
timestamp 1688980957
transform 1 0 22080 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_237
timestamp 1688980957
transform 1 0 22908 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_261
timestamp 1688980957
transform 1 0 25116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_270
timestamp 1688980957
transform 1 0 25944 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_274
timestamp 1688980957
transform 1 0 26312 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_278
timestamp 1688980957
transform 1 0 26680 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_290
timestamp 1688980957
transform 1 0 27784 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_305
timestamp 1688980957
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_347
timestamp 1688980957
transform 1 0 33028 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_371
timestamp 1688980957
transform 1 0 35236 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_383
timestamp 1688980957
transform 1 0 36340 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_395
timestamp 1688980957
transform 1 0 37444 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_85
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_100
timestamp 1688980957
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_156
timestamp 1688980957
transform 1 0 15456 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_180
timestamp 1688980957
transform 1 0 17664 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_209
timestamp 1688980957
transform 1 0 20332 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_216
timestamp 1688980957
transform 1 0 20976 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_241
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_262
timestamp 1688980957
transform 1 0 25208 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_270
timestamp 1688980957
transform 1 0 25944 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_331
timestamp 1688980957
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_367
timestamp 1688980957
transform 1 0 34868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_379
timestamp 1688980957
transform 1 0 35972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_57
timestamp 1688980957
transform 1 0 6348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_61
timestamp 1688980957
transform 1 0 6716 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_94
timestamp 1688980957
transform 1 0 9752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_100
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_112
timestamp 1688980957
transform 1 0 11408 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_120
timestamp 1688980957
transform 1 0 12144 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_145
timestamp 1688980957
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_155
timestamp 1688980957
transform 1 0 15364 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_193
timestamp 1688980957
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_202
timestamp 1688980957
transform 1 0 19688 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_210
timestamp 1688980957
transform 1 0 20424 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_225
timestamp 1688980957
transform 1 0 21804 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_243
timestamp 1688980957
transform 1 0 23460 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_270
timestamp 1688980957
transform 1 0 25944 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_285
timestamp 1688980957
transform 1 0 27324 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_297
timestamp 1688980957
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_302
timestamp 1688980957
transform 1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_347
timestamp 1688980957
transform 1 0 33028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_362
timestamp 1688980957
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_388
timestamp 1688980957
transform 1 0 36800 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_400
timestamp 1688980957
transform 1 0 37904 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_34
timestamp 1688980957
transform 1 0 4232 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_40
timestamp 1688980957
transform 1 0 4784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_44
timestamp 1688980957
transform 1 0 5152 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_66
timestamp 1688980957
transform 1 0 7176 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_110
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_122
timestamp 1688980957
transform 1 0 12328 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_128
timestamp 1688980957
transform 1 0 12880 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_189
timestamp 1688980957
transform 1 0 18492 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_219
timestamp 1688980957
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_241
timestamp 1688980957
transform 1 0 23276 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_267
timestamp 1688980957
transform 1 0 25668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_287
timestamp 1688980957
transform 1 0 27508 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_296
timestamp 1688980957
transform 1 0 28336 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_310
timestamp 1688980957
transform 1 0 29624 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_318
timestamp 1688980957
transform 1 0 30360 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_322
timestamp 1688980957
transform 1 0 30728 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_340
timestamp 1688980957
transform 1 0 32384 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_352
timestamp 1688980957
transform 1 0 33488 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_364
timestamp 1688980957
transform 1 0 34592 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_369
timestamp 1688980957
transform 1 0 35052 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_381
timestamp 1688980957
transform 1 0 36156 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_389
timestamp 1688980957
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_94
timestamp 1688980957
transform 1 0 9752 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_129
timestamp 1688980957
transform 1 0 12972 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_136
timestamp 1688980957
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_151
timestamp 1688980957
transform 1 0 14996 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_163
timestamp 1688980957
transform 1 0 16100 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_175
timestamp 1688980957
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_187
timestamp 1688980957
transform 1 0 18308 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_194
timestamp 1688980957
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_228
timestamp 1688980957
transform 1 0 22080 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_234
timestamp 1688980957
transform 1 0 22632 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_242
timestamp 1688980957
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_250
timestamp 1688980957
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_261
timestamp 1688980957
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_271
timestamp 1688980957
transform 1 0 26036 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_283
timestamp 1688980957
transform 1 0 27140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_295
timestamp 1688980957
transform 1 0 28244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_350
timestamp 1688980957
transform 1 0 33304 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1688980957
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_75
timestamp 1688980957
transform 1 0 8004 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_87
timestamp 1688980957
transform 1 0 9108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_99
timestamp 1688980957
transform 1 0 10212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_103
timestamp 1688980957
transform 1 0 10580 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_107
timestamp 1688980957
transform 1 0 10948 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_219
timestamp 1688980957
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_233
timestamp 1688980957
transform 1 0 22540 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_252
timestamp 1688980957
transform 1 0 24288 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_260
timestamp 1688980957
transform 1 0 25024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_304
timestamp 1688980957
transform 1 0 29072 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_324
timestamp 1688980957
transform 1 0 30912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_340
timestamp 1688980957
transform 1 0 32384 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_387
timestamp 1688980957
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1688980957
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_47
timestamp 1688980957
transform 1 0 5428 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_59
timestamp 1688980957
transform 1 0 6532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_67
timestamp 1688980957
transform 1 0 7268 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_82
timestamp 1688980957
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_93
timestamp 1688980957
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_104
timestamp 1688980957
transform 1 0 10672 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_116
timestamp 1688980957
transform 1 0 11776 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_129
timestamp 1688980957
transform 1 0 12972 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_137
timestamp 1688980957
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_169
timestamp 1688980957
transform 1 0 16652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_176
timestamp 1688980957
transform 1 0 17296 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_190
timestamp 1688980957
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_226
timestamp 1688980957
transform 1 0 21896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_273
timestamp 1688980957
transform 1 0 26220 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_278
timestamp 1688980957
transform 1 0 26680 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_285
timestamp 1688980957
transform 1 0 27324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_303
timestamp 1688980957
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_318
timestamp 1688980957
transform 1 0 30360 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_330
timestamp 1688980957
transform 1 0 31464 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_342
timestamp 1688980957
transform 1 0 32568 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_371
timestamp 1688980957
transform 1 0 35236 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_383
timestamp 1688980957
transform 1 0 36340 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_395
timestamp 1688980957
transform 1 0 37444 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_63
timestamp 1688980957
transform 1 0 6900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_85
timestamp 1688980957
transform 1 0 8924 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_121
timestamp 1688980957
transform 1 0 12236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_133
timestamp 1688980957
transform 1 0 13340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_141
timestamp 1688980957
transform 1 0 14076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_182
timestamp 1688980957
transform 1 0 17848 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_206
timestamp 1688980957
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_218
timestamp 1688980957
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_232
timestamp 1688980957
transform 1 0 22448 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_244
timestamp 1688980957
transform 1 0 23552 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_250
timestamp 1688980957
transform 1 0 24104 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_256
timestamp 1688980957
transform 1 0 24656 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_268
timestamp 1688980957
transform 1 0 25760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_315
timestamp 1688980957
transform 1 0 30084 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_327
timestamp 1688980957
transform 1 0 31188 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_366
timestamp 1688980957
transform 1 0 34776 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_378
timestamp 1688980957
transform 1 0 35880 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_390
timestamp 1688980957
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_397
timestamp 1688980957
transform 1 0 37628 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_35
timestamp 1688980957
transform 1 0 4324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_39
timestamp 1688980957
transform 1 0 4692 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_45
timestamp 1688980957
transform 1 0 5244 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_49
timestamp 1688980957
transform 1 0 5612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_61
timestamp 1688980957
transform 1 0 6716 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_68
timestamp 1688980957
transform 1 0 7360 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_76
timestamp 1688980957
transform 1 0 8096 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_82
timestamp 1688980957
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_101
timestamp 1688980957
transform 1 0 10396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_113
timestamp 1688980957
transform 1 0 11500 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_126
timestamp 1688980957
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_138
timestamp 1688980957
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_154
timestamp 1688980957
transform 1 0 15272 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_162
timestamp 1688980957
transform 1 0 16008 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_178
timestamp 1688980957
transform 1 0 17480 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_187
timestamp 1688980957
transform 1 0 18308 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_193
timestamp 1688980957
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_216
timestamp 1688980957
transform 1 0 20976 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_228
timestamp 1688980957
transform 1 0 22080 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_240
timestamp 1688980957
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_269
timestamp 1688980957
transform 1 0 25852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_290
timestamp 1688980957
transform 1 0 27784 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_294
timestamp 1688980957
transform 1 0 28152 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_298
timestamp 1688980957
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 1688980957
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_318
timestamp 1688980957
transform 1 0 30360 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_361
timestamp 1688980957
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_66
timestamp 1688980957
transform 1 0 7176 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_72
timestamp 1688980957
transform 1 0 7728 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_94
timestamp 1688980957
transform 1 0 9752 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_106
timestamp 1688980957
transform 1 0 10856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_119
timestamp 1688980957
transform 1 0 12052 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_128
timestamp 1688980957
transform 1 0 12880 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_140
timestamp 1688980957
transform 1 0 13984 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_152
timestamp 1688980957
transform 1 0 15088 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_164
timestamp 1688980957
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_184
timestamp 1688980957
transform 1 0 18032 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_196
timestamp 1688980957
transform 1 0 19136 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_215
timestamp 1688980957
transform 1 0 20884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_232
timestamp 1688980957
transform 1 0 22448 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_250
timestamp 1688980957
transform 1 0 24104 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_258
timestamp 1688980957
transform 1 0 24840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_268
timestamp 1688980957
transform 1 0 25760 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_277
timestamp 1688980957
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_302
timestamp 1688980957
transform 1 0 28888 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_312
timestamp 1688980957
transform 1 0 29808 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_320
timestamp 1688980957
transform 1 0 30544 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_333
timestamp 1688980957
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1688980957
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1688980957
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_35
timestamp 1688980957
transform 1 0 4324 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_39
timestamp 1688980957
transform 1 0 4692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_51
timestamp 1688980957
transform 1 0 5796 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_62
timestamp 1688980957
transform 1 0 6808 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_93
timestamp 1688980957
transform 1 0 9660 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_120
timestamp 1688980957
transform 1 0 12144 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_132
timestamp 1688980957
transform 1 0 13248 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_148
timestamp 1688980957
transform 1 0 14720 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_160
timestamp 1688980957
transform 1 0 15824 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_172
timestamp 1688980957
transform 1 0 16928 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_184
timestamp 1688980957
transform 1 0 18032 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_205
timestamp 1688980957
transform 1 0 19964 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_213
timestamp 1688980957
transform 1 0 20700 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_224
timestamp 1688980957
transform 1 0 21712 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_228
timestamp 1688980957
transform 1 0 22080 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_237
timestamp 1688980957
transform 1 0 22908 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_247
timestamp 1688980957
transform 1 0 23828 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_272
timestamp 1688980957
transform 1 0 26128 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_280
timestamp 1688980957
transform 1 0 26864 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_292
timestamp 1688980957
transform 1 0 27968 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_304
timestamp 1688980957
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_330
timestamp 1688980957
transform 1 0 31464 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_342
timestamp 1688980957
transform 1 0 32568 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_354
timestamp 1688980957
transform 1 0 33672 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_362
timestamp 1688980957
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_47
timestamp 1688980957
transform 1 0 5428 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_68
timestamp 1688980957
transform 1 0 7360 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_72
timestamp 1688980957
transform 1 0 7728 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_82
timestamp 1688980957
transform 1 0 8648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_92
timestamp 1688980957
transform 1 0 9568 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_106
timestamp 1688980957
transform 1 0 10856 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_122
timestamp 1688980957
transform 1 0 12328 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_136
timestamp 1688980957
transform 1 0 13616 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_151
timestamp 1688980957
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_163
timestamp 1688980957
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_243
timestamp 1688980957
transform 1 0 23460 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_255
timestamp 1688980957
transform 1 0 24564 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_269
timestamp 1688980957
transform 1 0 25852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_277
timestamp 1688980957
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_312
timestamp 1688980957
transform 1 0 29808 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_343
timestamp 1688980957
transform 1 0 32660 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_353
timestamp 1688980957
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_365
timestamp 1688980957
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_377
timestamp 1688980957
transform 1 0 35788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_389
timestamp 1688980957
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_37
timestamp 1688980957
transform 1 0 4508 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_106
timestamp 1688980957
transform 1 0 10856 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_118
timestamp 1688980957
transform 1 0 11960 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_137
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_149
timestamp 1688980957
transform 1 0 14812 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_158
timestamp 1688980957
transform 1 0 15640 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_170
timestamp 1688980957
transform 1 0 16744 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_176
timestamp 1688980957
transform 1 0 17296 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_187
timestamp 1688980957
transform 1 0 18308 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_201
timestamp 1688980957
transform 1 0 19596 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_216
timestamp 1688980957
transform 1 0 20976 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_228
timestamp 1688980957
transform 1 0 22080 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_236
timestamp 1688980957
transform 1 0 22816 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_244
timestamp 1688980957
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_273
timestamp 1688980957
transform 1 0 26220 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_282
timestamp 1688980957
transform 1 0 27048 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_320
timestamp 1688980957
transform 1 0 30544 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_325
timestamp 1688980957
transform 1 0 31004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_337
timestamp 1688980957
transform 1 0 32108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_362
timestamp 1688980957
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_63
timestamp 1688980957
transform 1 0 6900 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_67
timestamp 1688980957
transform 1 0 7268 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_79
timestamp 1688980957
transform 1 0 8372 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_91
timestamp 1688980957
transform 1 0 9476 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_103
timestamp 1688980957
transform 1 0 10580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_233
timestamp 1688980957
transform 1 0 22540 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_240
timestamp 1688980957
transform 1 0 23184 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_252
timestamp 1688980957
transform 1 0 24288 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_260
timestamp 1688980957
transform 1 0 25024 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_269
timestamp 1688980957
transform 1 0 25852 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_277
timestamp 1688980957
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_287
timestamp 1688980957
transform 1 0 27508 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_291
timestamp 1688980957
transform 1 0 27876 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_303
timestamp 1688980957
transform 1 0 28980 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_315
timestamp 1688980957
transform 1 0 30084 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_327
timestamp 1688980957
transform 1 0 31188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_343
timestamp 1688980957
transform 1 0 32660 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_347
timestamp 1688980957
transform 1 0 33028 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_359
timestamp 1688980957
transform 1 0 34132 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_371
timestamp 1688980957
transform 1 0 35236 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_383
timestamp 1688980957
transform 1 0 36340 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_9
timestamp 1688980957
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_21
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_88
timestamp 1688980957
transform 1 0 9200 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_100
timestamp 1688980957
transform 1 0 10304 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_112
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_124
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_136
timestamp 1688980957
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_154
timestamp 1688980957
transform 1 0 15272 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_166
timestamp 1688980957
transform 1 0 16376 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_178
timestamp 1688980957
transform 1 0 17480 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_190
timestamp 1688980957
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_205
timestamp 1688980957
transform 1 0 19964 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_217
timestamp 1688980957
transform 1 0 21068 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_225
timestamp 1688980957
transform 1 0 21804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_241
timestamp 1688980957
transform 1 0 23276 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_250
timestamp 1688980957
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_262
timestamp 1688980957
transform 1 0 25208 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_274
timestamp 1688980957
transform 1 0 26312 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_280
timestamp 1688980957
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_286
timestamp 1688980957
transform 1 0 27416 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_298
timestamp 1688980957
transform 1 0 28520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_306
timestamp 1688980957
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_331
timestamp 1688980957
transform 1 0 31556 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_343
timestamp 1688980957
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_355
timestamp 1688980957
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_395
timestamp 1688980957
transform 1 0 37444 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_77
timestamp 1688980957
transform 1 0 8188 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_116
timestamp 1688980957
transform 1 0 11776 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_120
timestamp 1688980957
transform 1 0 12144 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_130
timestamp 1688980957
transform 1 0 13064 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_138
timestamp 1688980957
transform 1 0 13800 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_151
timestamp 1688980957
transform 1 0 14996 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_164
timestamp 1688980957
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_175
timestamp 1688980957
transform 1 0 17204 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_183
timestamp 1688980957
transform 1 0 17940 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_191
timestamp 1688980957
transform 1 0 18676 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_204
timestamp 1688980957
transform 1 0 19872 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_232
timestamp 1688980957
transform 1 0 22448 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_240
timestamp 1688980957
transform 1 0 23184 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_252
timestamp 1688980957
transform 1 0 24288 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_296
timestamp 1688980957
transform 1 0 28336 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_300
timestamp 1688980957
transform 1 0 28704 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_313
timestamp 1688980957
transform 1 0 29900 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 1688980957
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_340
timestamp 1688980957
transform 1 0 32384 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_352
timestamp 1688980957
transform 1 0 33488 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_364
timestamp 1688980957
transform 1 0 34592 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_376
timestamp 1688980957
transform 1 0 35696 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_388
timestamp 1688980957
transform 1 0 36800 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_45
timestamp 1688980957
transform 1 0 5244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_57
timestamp 1688980957
transform 1 0 6348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_69
timestamp 1688980957
transform 1 0 7452 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_92
timestamp 1688980957
transform 1 0 9568 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_243
timestamp 1688980957
transform 1 0 23460 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_277
timestamp 1688980957
transform 1 0 26588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_302
timestamp 1688980957
transform 1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_330
timestamp 1688980957
transform 1 0 31464 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_340
timestamp 1688980957
transform 1 0 32384 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_352
timestamp 1688980957
transform 1 0 33488 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_368
timestamp 1688980957
transform 1 0 34960 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_380
timestamp 1688980957
transform 1 0 36064 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_392
timestamp 1688980957
transform 1 0 37168 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_9
timestamp 1688980957
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_21
timestamp 1688980957
transform 1 0 3036 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_29
timestamp 1688980957
transform 1 0 3772 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_37
timestamp 1688980957
transform 1 0 4508 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_44
timestamp 1688980957
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_85
timestamp 1688980957
transform 1 0 8924 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_119
timestamp 1688980957
transform 1 0 12052 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_127
timestamp 1688980957
transform 1 0 12788 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_133
timestamp 1688980957
transform 1 0 13340 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_139
timestamp 1688980957
transform 1 0 13892 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_141
timestamp 1688980957
transform 1 0 14076 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_153
timestamp 1688980957
transform 1 0 15180 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_177
timestamp 1688980957
transform 1 0 17388 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_184
timestamp 1688980957
transform 1 0 18032 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_197
timestamp 1688980957
transform 1 0 19228 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_216
timestamp 1688980957
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_233
timestamp 1688980957
transform 1 0 22540 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_245
timestamp 1688980957
transform 1 0 23644 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_251
timestamp 1688980957
transform 1 0 24196 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_253
timestamp 1688980957
transform 1 0 24380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_260
timestamp 1688980957
transform 1 0 25024 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_268
timestamp 1688980957
transform 1 0 25760 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_275
timestamp 1688980957
transform 1 0 26404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_287
timestamp 1688980957
transform 1 0 27508 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_299
timestamp 1688980957
transform 1 0 28612 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_307
timestamp 1688980957
transform 1 0 29348 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_309
timestamp 1688980957
transform 1 0 29532 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_321
timestamp 1688980957
transform 1 0 30636 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_345
timestamp 1688980957
transform 1 0 32844 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_352
timestamp 1688980957
transform 1 0 33488 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_365
timestamp 1688980957
transform 1 0 34684 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_380
timestamp 1688980957
transform 1 0 36064 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_399
timestamp 1688980957
transform 1 0 37812 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 8096 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 9016 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 8004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1688980957
transform 1 0 37444 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1688980957
transform 1 0 31004 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform 1 0 15548 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 37444 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1688980957
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap47
timestamp 1688980957
transform 1 0 7084 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  max_cap48
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  max_cap49
timestamp 1688980957
transform 1 0 22264 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap51
timestamp 1688980957
transform 1 0 19136 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap52
timestamp 1688980957
transform 1 0 18584 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap53
timestamp 1688980957
transform 1 0 17020 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  max_cap54
timestamp 1688980957
transform 1 0 21528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1688980957
transform 1 0 17664 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1688980957
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 21988 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 37444 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1688980957
transform 1 0 12972 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform 1 0 3956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1688980957
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 37444 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1688980957
transform 1 0 9292 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 6532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1688980957
transform 1 0 37628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 19412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 35512 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform 1 0 32936 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1688980957
transform 1 0 4784 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 1688980957
transform 1 0 37444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 38272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 38272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 38272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 38272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 38272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 38272 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 38272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 38272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 38272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 38272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 38272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 38272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 38272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 38272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 38272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 38272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 38272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 38272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 38272 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 38272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 38272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 38272 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 38272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 38272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 38272 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 38272 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 38272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 38272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 38272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 38272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 38272 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 38272 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 38272 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 38272 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 38272 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 38272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 38272 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 38272 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 38272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 38272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 38272 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 38272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 38272 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 38272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 38272 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 38272 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 38272 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 38272 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 3680 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 8832 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 13984 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 19136 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 24288 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 29440 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 34592 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire50
timestamp 1688980957
transform 1 0 23184 0 1 23936
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 38618 8848 39418 8968 0 FreeSans 480 0 0 0 cs
port 1 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 gpi[0]
port 2 nsew signal input
flabel metal3 s 38618 29248 39418 29368 0 FreeSans 480 0 0 0 gpi[10]
port 3 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 gpi[11]
port 4 nsew signal input
flabel metal3 s 38618 13608 39418 13728 0 FreeSans 480 0 0 0 gpi[12]
port 5 nsew signal input
flabel metal2 s 1950 40762 2006 41562 0 FreeSans 224 90 0 0 gpi[13]
port 6 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 gpi[14]
port 7 nsew signal input
flabel metal3 s 38618 25168 39418 25288 0 FreeSans 480 0 0 0 gpi[15]
port 8 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 gpi[16]
port 9 nsew signal input
flabel metal3 s 38618 4088 39418 4208 0 FreeSans 480 0 0 0 gpi[17]
port 10 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 gpi[18]
port 11 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 gpi[19]
port 12 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 gpi[1]
port 13 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 gpi[20]
port 14 nsew signal input
flabel metal3 s 38618 6128 39418 6248 0 FreeSans 480 0 0 0 gpi[21]
port 15 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 gpi[22]
port 16 nsew signal input
flabel metal2 s 30930 40762 30986 41562 0 FreeSans 224 90 0 0 gpi[23]
port 17 nsew signal input
flabel metal2 s 28354 40762 28410 41562 0 FreeSans 224 90 0 0 gpi[24]
port 18 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 gpi[25]
port 19 nsew signal input
flabel metal3 s 38618 27208 39418 27328 0 FreeSans 480 0 0 0 gpi[26]
port 20 nsew signal input
flabel metal3 s 38618 31968 39418 32088 0 FreeSans 480 0 0 0 gpi[27]
port 21 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpi[28]
port 22 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpi[29]
port 23 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpi[2]
port 24 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 gpi[30]
port 25 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 gpi[31]
port 26 nsew signal input
flabel metal2 s 24490 40762 24546 41562 0 FreeSans 224 90 0 0 gpi[32]
port 27 nsew signal input
flabel metal2 s 6458 40762 6514 41562 0 FreeSans 224 90 0 0 gpi[33]
port 28 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpi[3]
port 29 nsew signal input
flabel metal2 s 15474 40762 15530 41562 0 FreeSans 224 90 0 0 gpi[4]
port 30 nsew signal input
flabel metal2 s 37370 40762 37426 41562 0 FreeSans 224 90 0 0 gpi[5]
port 31 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 gpi[6]
port 32 nsew signal input
flabel metal2 s 19982 40762 20038 41562 0 FreeSans 224 90 0 0 gpi[7]
port 33 nsew signal input
flabel metal2 s 39302 40762 39358 41562 0 FreeSans 224 90 0 0 gpi[8]
port 34 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gpi[9]
port 35 nsew signal input
flabel metal2 s 17406 40762 17462 41562 0 FreeSans 224 90 0 0 gpo[0]
port 36 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 gpo[10]
port 37 nsew signal tristate
flabel metal3 s 38618 10888 39418 11008 0 FreeSans 480 0 0 0 gpo[11]
port 38 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gpo[12]
port 39 nsew signal tristate
flabel metal3 s 38618 15648 39418 15768 0 FreeSans 480 0 0 0 gpo[13]
port 40 nsew signal tristate
flabel metal2 s 18 40762 74 41562 0 FreeSans 224 90 0 0 gpo[14]
port 41 nsew signal tristate
flabel metal2 s 26422 40762 26478 41562 0 FreeSans 224 90 0 0 gpo[15]
port 42 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpo[16]
port 43 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpo[17]
port 44 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 gpo[18]
port 45 nsew signal tristate
flabel metal2 s 21914 40762 21970 41562 0 FreeSans 224 90 0 0 gpo[19]
port 46 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gpo[1]
port 47 nsew signal tristate
flabel metal3 s 38618 38768 39418 38888 0 FreeSans 480 0 0 0 gpo[20]
port 48 nsew signal tristate
flabel metal2 s 12898 40762 12954 41562 0 FreeSans 224 90 0 0 gpo[21]
port 49 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpo[22]
port 50 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpo[23]
port 51 nsew signal tristate
flabel metal3 s 38618 36728 39418 36848 0 FreeSans 480 0 0 0 gpo[24]
port 52 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 gpo[25]
port 53 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpo[26]
port 54 nsew signal tristate
flabel metal3 s 38618 34008 39418 34128 0 FreeSans 480 0 0 0 gpo[27]
port 55 nsew signal tristate
flabel metal3 s 38618 1368 39418 1488 0 FreeSans 480 0 0 0 gpo[28]
port 56 nsew signal tristate
flabel metal2 s 9034 40762 9090 41562 0 FreeSans 224 90 0 0 gpo[29]
port 57 nsew signal tristate
flabel metal3 s 38618 20408 39418 20528 0 FreeSans 480 0 0 0 gpo[2]
port 58 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpo[30]
port 59 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpo[31]
port 60 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 gpo[32]
port 61 nsew signal tristate
flabel metal3 s 38618 22448 39418 22568 0 FreeSans 480 0 0 0 gpo[33]
port 62 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpo[3]
port 63 nsew signal tristate
flabel metal2 s 35438 40762 35494 41562 0 FreeSans 224 90 0 0 gpo[4]
port 64 nsew signal tristate
flabel metal2 s 32862 40762 32918 41562 0 FreeSans 224 90 0 0 gpo[5]
port 65 nsew signal tristate
flabel metal2 s 4526 40762 4582 41562 0 FreeSans 224 90 0 0 gpo[6]
port 66 nsew signal tristate
flabel metal2 s 10966 40762 11022 41562 0 FreeSans 224 90 0 0 gpo[7]
port 67 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 gpo[8]
port 68 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 gpo[9]
port 69 nsew signal tristate
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 nrst
port 70 nsew signal input
flabel metal3 s 38618 17688 39418 17808 0 FreeSans 480 0 0 0 store_en
port 71 nsew signal tristate
flabel metal4 s 4208 2128 4528 39216 0 FreeSans 1920 90 0 0 vccd1
port 72 nsew power bidirectional
flabel metal4 s 34928 2128 35248 39216 0 FreeSans 1920 90 0 0 vccd1
port 72 nsew power bidirectional
flabel metal4 s 19568 2128 19888 39216 0 FreeSans 1920 90 0 0 vssd1
port 73 nsew ground bidirectional
rlabel metal1 19688 38624 19688 38624 0 vccd1
rlabel via1 19688 39168 19688 39168 0 vssd1
rlabel metal1 15548 23698 15548 23698 0 ALU.flags_to_alu\[0\]
rlabel metal2 17986 33626 17986 33626 0 ALU.flags_to_alu\[1\]
rlabel metal1 17710 26282 17710 26282 0 ALU.flags_to_alu\[2\]
rlabel metal1 8832 30022 8832 30022 0 ALU.flags_to_alu\[3\]
rlabel metal1 18584 28118 18584 28118 0 ALU.flags_to_alu\[4\]
rlabel metal1 8786 31790 8786 31790 0 ALU.flags_to_alu\[5\]
rlabel metal1 19458 37910 19458 37910 0 ALU.flags_to_alu\[6\]
rlabel metal1 21390 35156 21390 35156 0 ALU.flags_to_alu\[7\]
rlabel metal1 17158 10234 17158 10234 0 ALU.immediate\[0\]
rlabel metal1 7774 11662 7774 11662 0 ALU.immediate\[10\]
rlabel metal1 18814 22168 18814 22168 0 ALU.immediate\[11\]
rlabel metal1 14214 22474 14214 22474 0 ALU.immediate\[12\]
rlabel metal1 7774 15130 7774 15130 0 ALU.immediate\[13\]
rlabel metal2 5934 21862 5934 21862 0 ALU.immediate\[14\]
rlabel via1 8694 19363 8694 19363 0 ALU.immediate\[15\]
rlabel metal2 17066 7140 17066 7140 0 ALU.immediate\[1\]
rlabel metal2 14766 8092 14766 8092 0 ALU.immediate\[2\]
rlabel metal1 14030 10642 14030 10642 0 ALU.immediate\[3\]
rlabel metal2 9522 13464 9522 13464 0 ALU.immediate\[4\]
rlabel metal1 12650 13158 12650 13158 0 ALU.immediate\[5\]
rlabel via2 12926 16405 12926 16405 0 ALU.immediate\[6\]
rlabel metal1 22080 15640 22080 15640 0 ALU.immediate\[7\]
rlabel metal2 26450 17935 26450 17935 0 ALU.immediate\[8\]
rlabel via2 4094 20451 4094 20451 0 ALU.immediate\[9\]
rlabel metal2 11638 7616 11638 7616 0 ByteBuffer.counter\[0\]
rlabel metal1 11362 7888 11362 7888 0 ByteBuffer.counter\[1\]
rlabel metal1 16698 10642 16698 10642 0 ByteBuffer.instr\[16\]
rlabel metal2 18078 18292 18078 18292 0 ByteBuffer.instr\[17\]
rlabel metal1 18492 8466 18492 8466 0 ByteBuffer.instr\[18\]
rlabel viali 19734 17170 19734 17170 0 ByteBuffer.instr\[19\]
rlabel metal1 14214 20400 14214 20400 0 ByteBuffer.instr\[20\]
rlabel metal1 16192 19346 16192 19346 0 ByteBuffer.instr\[21\]
rlabel metal1 13110 7922 13110 7922 0 ByteBuffer.instr\[22\]
rlabel metal1 14122 14994 14122 14994 0 ByteBuffer.instr\[23\]
rlabel metal1 11040 7854 11040 7854 0 ByteBuffer.next_counter\[0\]
rlabel metal1 9292 7514 9292 7514 0 ByteBuffer.next_counter\[1\]
rlabel metal1 8464 6290 8464 6290 0 ByteDecoder.num_bytes\[1\]
rlabel metal1 8280 4454 8280 4454 0 ByteDecoder.num_bytes\[2\]
rlabel metal1 8188 5678 8188 5678 0 ByteDecoder.num_bytes\[3\]
rlabel metal2 9338 5440 9338 5440 0 ByteDecoder.state\[0\]
rlabel metal1 12466 5168 12466 5168 0 ByteDecoder.state\[1\]
rlabel metal1 9660 5746 9660 5746 0 FSM.next_state\[0\]
rlabel metal1 9522 4760 9522 4760 0 FSM.next_state\[1\]
rlabel metal1 14950 5576 14950 5576 0 MemControl.state\[0\]
rlabel metal1 13800 5202 13800 5202 0 MemControl.state\[1\]
rlabel metal1 13708 5338 13708 5338 0 MemControl.state\[2\]
rlabel metal1 4784 8262 4784 8262 0 PC.i_mem_addr\[0\]
rlabel metal1 2438 22678 2438 22678 0 PC.i_mem_addr\[10\]
rlabel metal1 4554 21998 4554 21998 0 PC.i_mem_addr\[11\]
rlabel metal1 7728 22610 7728 22610 0 PC.i_mem_addr\[12\]
rlabel metal1 6808 23018 6808 23018 0 PC.i_mem_addr\[13\]
rlabel metal2 4830 24378 4830 24378 0 PC.i_mem_addr\[14\]
rlabel metal1 5750 19822 5750 19822 0 PC.i_mem_addr\[15\]
rlabel metal1 4554 7378 4554 7378 0 PC.i_mem_addr\[1\]
rlabel metal1 4140 9554 4140 9554 0 PC.i_mem_addr\[2\]
rlabel metal1 5244 10506 5244 10506 0 PC.i_mem_addr\[3\]
rlabel metal1 2530 11152 2530 11152 0 PC.i_mem_addr\[4\]
rlabel metal1 4692 13702 4692 13702 0 PC.i_mem_addr\[5\]
rlabel metal1 4278 17068 4278 17068 0 PC.i_mem_addr\[6\]
rlabel metal1 7176 17510 7176 17510 0 PC.i_mem_addr\[7\]
rlabel via2 17986 16507 17986 16507 0 PC.i_mem_addr\[8\]
rlabel metal1 3864 20978 3864 20978 0 PC.i_mem_addr\[9\]
rlabel metal3 20401 17340 20401 17340 0 RegFile.A\[0\]
rlabel metal1 24610 33456 24610 33456 0 RegFile.A\[1\]
rlabel metal1 16146 25908 16146 25908 0 RegFile.A\[2\]
rlabel metal2 28934 29274 28934 29274 0 RegFile.A\[3\]
rlabel metal1 17250 25772 17250 25772 0 RegFile.A\[4\]
rlabel metal1 32890 31858 32890 31858 0 RegFile.A\[5\]
rlabel metal1 14490 35666 14490 35666 0 RegFile.A\[6\]
rlabel metal1 35236 31654 35236 31654 0 RegFile.A\[7\]
rlabel metal1 29578 24752 29578 24752 0 RegFile.B\[0\]
rlabel viali 29210 34578 29210 34578 0 RegFile.B\[1\]
rlabel metal1 16422 26282 16422 26282 0 RegFile.B\[2\]
rlabel metal1 16422 29614 16422 29614 0 RegFile.B\[3\]
rlabel metal2 26358 28220 26358 28220 0 RegFile.B\[4\]
rlabel via1 29762 32402 29762 32402 0 RegFile.B\[5\]
rlabel metal1 25254 36176 25254 36176 0 RegFile.B\[6\]
rlabel metal1 25530 35598 25530 35598 0 RegFile.B\[7\]
rlabel metal1 19642 24344 19642 24344 0 RegFile.C\[0\]
rlabel metal1 8464 35802 8464 35802 0 RegFile.C\[1\]
rlabel metal1 17250 27370 17250 27370 0 RegFile.C\[2\]
rlabel metal1 17020 30702 17020 30702 0 RegFile.C\[3\]
rlabel metal1 10028 27846 10028 27846 0 RegFile.C\[4\]
rlabel metal1 8510 32878 8510 32878 0 RegFile.C\[5\]
rlabel metal1 17618 37944 17618 37944 0 RegFile.C\[6\]
rlabel metal1 19274 37264 19274 37264 0 RegFile.C\[7\]
rlabel metal2 23138 25602 23138 25602 0 RegFile.D\[0\]
rlabel metal1 25162 34544 25162 34544 0 RegFile.D\[1\]
rlabel metal1 26588 27302 26588 27302 0 RegFile.D\[2\]
rlabel metal1 19366 30192 19366 30192 0 RegFile.D\[3\]
rlabel viali 25438 28523 25438 28523 0 RegFile.D\[4\]
rlabel metal1 25300 31790 25300 31790 0 RegFile.D\[5\]
rlabel metal1 25346 37910 25346 37910 0 RegFile.D\[6\]
rlabel metal2 31786 37264 31786 37264 0 RegFile.D\[7\]
rlabel metal1 7176 26282 7176 26282 0 RegFile.E\[0\]
rlabel metal1 7912 34986 7912 34986 0 RegFile.E\[1\]
rlabel metal1 11960 27030 11960 27030 0 RegFile.E\[2\]
rlabel metal1 15088 30566 15088 30566 0 RegFile.E\[3\]
rlabel metal1 6992 27846 6992 27846 0 RegFile.E\[4\]
rlabel metal1 6210 31654 6210 31654 0 RegFile.E\[5\]
rlabel metal1 18492 37842 18492 37842 0 RegFile.E\[6\]
rlabel metal1 21160 37910 21160 37910 0 RegFile.E\[7\]
rlabel metal2 22494 23698 22494 23698 0 RegFile.H\[0\]
rlabel via1 31418 34170 31418 34170 0 RegFile.H\[1\]
rlabel metal2 32614 26384 32614 26384 0 RegFile.H\[2\]
rlabel metal1 21482 30668 21482 30668 0 RegFile.H\[3\]
rlabel metal2 25714 28152 25714 28152 0 RegFile.H\[4\]
rlabel metal1 34224 32266 34224 32266 0 RegFile.H\[5\]
rlabel metal1 29141 36278 29141 36278 0 RegFile.H\[6\]
rlabel metal1 25852 36822 25852 36822 0 RegFile.H\[7\]
rlabel metal1 16146 23732 16146 23732 0 RegFile.L\[0\]
rlabel metal1 7314 34578 7314 34578 0 RegFile.L\[1\]
rlabel metal1 16846 27370 16846 27370 0 RegFile.L\[2\]
rlabel metal1 16791 30634 16791 30634 0 RegFile.L\[3\]
rlabel metal2 16330 28594 16330 28594 0 RegFile.L\[4\]
rlabel metal2 6210 32606 6210 32606 0 RegFile.L\[5\]
rlabel metal1 20010 36142 20010 36142 0 RegFile.L\[6\]
rlabel metal2 12006 35496 12006 35496 0 RegFile.L\[7\]
rlabel metal1 15778 5780 15778 5780 0 _0000_
rlabel metal1 12558 4250 12558 4250 0 _0001_
rlabel metal1 14306 4658 14306 4658 0 _0066_
rlabel metal1 6670 5304 6670 5304 0 _0067_
rlabel metal1 7491 4794 7491 4794 0 _0068_
rlabel metal1 6670 6426 6670 6426 0 _0069_
rlabel metal1 5106 14042 5106 14042 0 _0070_
rlabel metal1 5612 12138 5612 12138 0 _0071_
rlabel metal1 6670 11832 6670 11832 0 _0072_
rlabel metal1 7268 20026 7268 20026 0 _0073_
rlabel metal1 7452 16218 7452 16218 0 _0074_
rlabel metal1 6624 14586 6624 14586 0 _0075_
rlabel metal1 6203 10234 6203 10234 0 _0076_
rlabel metal1 7360 18666 7360 18666 0 _0077_
rlabel metal1 15180 10710 15180 10710 0 _0078_
rlabel metal1 15870 11866 15870 11866 0 _0079_
rlabel metal1 16606 8398 16606 8398 0 _0080_
rlabel metal1 10396 12614 10396 12614 0 _0081_
rlabel metal1 9246 15368 9246 15368 0 _0082_
rlabel metal1 13202 11832 13202 11832 0 _0083_
rlabel metal1 13156 7446 13156 7446 0 _0084_
rlabel metal2 11822 14178 11822 14178 0 _0085_
rlabel metal1 15502 9928 15502 9928 0 _0086_
rlabel metal1 15318 6698 15318 6698 0 _0087_
rlabel metal1 14582 8398 14582 8398 0 _0088_
rlabel metal1 10350 9962 10350 9962 0 _0089_
rlabel metal2 8234 13600 8234 13600 0 _0090_
rlabel metal2 11822 10914 11822 10914 0 _0091_
rlabel metal1 12180 9146 12180 9146 0 _0092_
rlabel metal1 11132 15130 11132 15130 0 _0093_
rlabel metal1 10212 23154 10212 23154 0 _0094_
rlabel metal2 9798 33252 9798 33252 0 _0095_
rlabel metal1 10028 25330 10028 25330 0 _0096_
rlabel metal1 7176 30158 7176 30158 0 _0097_
rlabel metal1 8280 28730 8280 28730 0 _0098_
rlabel metal1 7774 31926 7774 31926 0 _0099_
rlabel metal1 10488 28730 10488 28730 0 _0100_
rlabel metal1 8280 34170 8280 34170 0 _0101_
rlabel metal1 5605 25466 5605 25466 0 _0102_
rlabel metal1 5014 34170 5014 34170 0 _0103_
rlabel metal1 8694 26486 8694 26486 0 _0104_
rlabel metal2 10718 31969 10718 31969 0 _0105_
rlabel metal2 5014 28832 5014 28832 0 _0106_
rlabel metal1 4922 33082 4922 33082 0 _0107_
rlabel metal1 9292 35802 9292 35802 0 _0108_
rlabel metal1 10580 35122 10580 35122 0 _0109_
rlabel metal1 24656 23290 24656 23290 0 _0110_
rlabel metal1 31188 34034 31188 34034 0 _0111_
rlabel metal2 31786 26146 31786 26146 0 _0112_
rlabel metal2 32430 30634 32430 30634 0 _0113_
rlabel metal2 31786 28322 31786 28322 0 _0114_
rlabel metal1 33350 32334 33350 32334 0 _0115_
rlabel metal1 27554 36074 27554 36074 0 _0116_
rlabel metal2 32798 36380 32798 36380 0 _0117_
rlabel metal1 5428 26282 5428 26282 0 _0118_
rlabel metal2 5566 35938 5566 35938 0 _0119_
rlabel metal1 10573 26554 10573 26554 0 _0120_
rlabel metal2 7774 31518 7774 31518 0 _0121_
rlabel metal2 4738 27880 4738 27880 0 _0122_
rlabel metal1 4554 31450 4554 31450 0 _0123_
rlabel metal1 12512 38726 12512 38726 0 _0124_
rlabel metal1 20838 38216 20838 38216 0 _0125_
rlabel metal1 24610 26010 24610 26010 0 _0126_
rlabel metal1 30590 35598 30590 35598 0 _0127_
rlabel metal2 27094 28322 27094 28322 0 _0128_
rlabel metal1 34592 30634 34592 30634 0 _0129_
rlabel metal1 34362 28152 34362 28152 0 _0130_
rlabel metal1 33672 33422 33672 33422 0 _0131_
rlabel metal1 25254 37978 25254 37978 0 _0132_
rlabel metal1 32154 37740 32154 37740 0 _0133_
rlabel metal1 8280 24854 8280 24854 0 _0134_
rlabel metal1 7360 35802 7360 35802 0 _0135_
rlabel metal1 11730 27982 11730 27982 0 _0136_
rlabel metal1 9890 30906 9890 30906 0 _0137_
rlabel metal1 7130 27642 7130 27642 0 _0138_
rlabel metal1 7452 33082 7452 33082 0 _0139_
rlabel metal1 10396 37978 10396 37978 0 _0140_
rlabel metal1 8832 37434 8832 37434 0 _0141_
rlabel metal1 28336 23766 28336 23766 0 _0142_
rlabel metal1 26818 34510 26818 34510 0 _0143_
rlabel metal1 27416 26418 27416 26418 0 _0144_
rlabel metal1 29348 30294 29348 30294 0 _0145_
rlabel metal1 29670 28458 29670 28458 0 _0146_
rlabel metal1 28198 33082 28198 33082 0 _0147_
rlabel metal1 26956 37978 26956 37978 0 _0148_
rlabel metal1 29762 37978 29762 37978 0 _0149_
rlabel metal1 29394 25976 29394 25976 0 _0150_
rlabel metal1 27094 32334 27094 32334 0 _0151_
rlabel metal1 34822 26282 34822 26282 0 _0152_
rlabel metal1 34822 29070 34822 29070 0 _0153_
rlabel metal1 34362 25466 34362 25466 0 _0154_
rlabel metal2 32154 32096 32154 32096 0 _0155_
rlabel metal1 26864 29818 26864 29818 0 _0156_
rlabel metal2 34270 32164 34270 32164 0 _0157_
rlabel metal1 6210 7514 6210 7514 0 _0158_
rlabel metal1 3772 6698 3772 6698 0 _0159_
rlabel metal1 1840 9146 1840 9146 0 _0160_
rlabel metal1 3174 10710 3174 10710 0 _0161_
rlabel metal1 1748 11798 1748 11798 0 _0162_
rlabel metal1 1840 13498 1840 13498 0 _0163_
rlabel metal1 1840 15130 1840 15130 0 _0164_
rlabel metal2 5106 17272 5106 17272 0 _0165_
rlabel metal1 1840 16762 1840 16762 0 _0166_
rlabel metal1 2024 20570 2024 20570 0 _0167_
rlabel metal1 2070 24922 2070 24922 0 _0168_
rlabel metal2 1794 23460 1794 23460 0 _0169_
rlabel metal1 6854 23834 6854 23834 0 _0170_
rlabel metal1 5244 22746 5244 22746 0 _0171_
rlabel metal1 3864 24378 3864 24378 0 _0172_
rlabel metal1 4738 18938 4738 18938 0 _0173_
rlabel metal2 28566 4454 28566 4454 0 _0174_
rlabel metal2 29302 6018 29302 6018 0 _0175_
rlabel metal1 26450 8908 26450 8908 0 _0176_
rlabel metal1 26404 7854 26404 7854 0 _0177_
rlabel metal1 27508 6834 27508 6834 0 _0178_
rlabel metal1 27738 6732 27738 6732 0 _0179_
rlabel metal1 28934 6732 28934 6732 0 _0180_
rlabel metal1 28106 6256 28106 6256 0 _0181_
rlabel metal1 28612 6766 28612 6766 0 _0182_
rlabel metal2 15134 19380 15134 19380 0 _0183_
rlabel metal1 35512 21862 35512 21862 0 _0184_
rlabel metal1 34178 21590 34178 21590 0 _0185_
rlabel metal2 34178 21522 34178 21522 0 _0186_
rlabel metal1 33166 21352 33166 21352 0 _0187_
rlabel metal1 28382 29478 28382 29478 0 _0188_
rlabel metal1 35190 29682 35190 29682 0 _0189_
rlabel metal1 22770 5236 22770 5236 0 _0190_
rlabel metal1 22954 5134 22954 5134 0 _0191_
rlabel metal1 24426 4624 24426 4624 0 _0192_
rlabel metal1 24794 4624 24794 4624 0 _0193_
rlabel metal1 20930 4794 20930 4794 0 _0194_
rlabel metal1 21873 4998 21873 4998 0 _0195_
rlabel metal1 25530 7412 25530 7412 0 _0196_
rlabel metal1 22402 8500 22402 8500 0 _0197_
rlabel metal1 25116 8806 25116 8806 0 _0198_
rlabel metal1 25530 7310 25530 7310 0 _0199_
rlabel metal1 25024 7446 25024 7446 0 _0200_
rlabel metal1 24886 5644 24886 5644 0 _0201_
rlabel metal1 24702 4726 24702 4726 0 _0202_
rlabel metal1 23920 4794 23920 4794 0 _0203_
rlabel via2 21942 18955 21942 18955 0 _0204_
rlabel metal1 34914 19958 34914 19958 0 _0205_
rlabel via1 35374 20298 35374 20298 0 _0206_
rlabel metal1 35696 20026 35696 20026 0 _0207_
rlabel via2 2438 21539 2438 21539 0 _0208_
rlabel metal1 24196 20842 24196 20842 0 _0209_
rlabel metal1 26128 20774 26128 20774 0 _0210_
rlabel metal1 33856 26554 33856 26554 0 _0211_
rlabel metal1 21206 6732 21206 6732 0 _0212_
rlabel metal1 22448 6766 22448 6766 0 _0213_
rlabel metal1 20056 5746 20056 5746 0 _0214_
rlabel metal2 22770 6086 22770 6086 0 _0215_
rlabel metal1 22310 7310 22310 7310 0 _0216_
rlabel metal1 20378 7412 20378 7412 0 _0217_
rlabel metal2 20562 7650 20562 7650 0 _0218_
rlabel metal1 22954 8398 22954 8398 0 _0219_
rlabel metal1 23230 7820 23230 7820 0 _0220_
rlabel metal1 22954 7378 22954 7378 0 _0221_
rlabel metal1 22494 6358 22494 6358 0 _0222_
rlabel metal1 23184 6426 23184 6426 0 _0223_
rlabel metal2 14030 19567 14030 19567 0 _0224_
rlabel metal1 34408 18666 34408 18666 0 _0225_
rlabel metal1 34914 18870 34914 18870 0 _0226_
rlabel metal1 35328 18326 35328 18326 0 _0227_
rlabel viali 33389 17612 33389 17612 0 _0228_
rlabel metal2 3174 19261 3174 19261 0 _0229_
rlabel metal1 26542 19482 26542 19482 0 _0230_
rlabel metal1 26220 32538 26220 32538 0 _0231_
rlabel metal1 22402 10064 22402 10064 0 _0232_
rlabel metal1 20930 9350 20930 9350 0 _0233_
rlabel metal1 21482 10132 21482 10132 0 _0234_
rlabel metal1 21620 10098 21620 10098 0 _0235_
rlabel metal1 22678 9996 22678 9996 0 _0236_
rlabel metal1 22816 9554 22816 9554 0 _0237_
rlabel metal2 22770 9248 22770 9248 0 _0238_
rlabel metal1 22356 10642 22356 10642 0 _0239_
rlabel metal1 23736 11730 23736 11730 0 _0240_
rlabel metal1 22494 9554 22494 9554 0 _0241_
rlabel metal1 22862 9690 22862 9690 0 _0242_
rlabel metal2 10304 12580 10304 12580 0 _0243_
rlabel metal2 28750 17340 28750 17340 0 _0244_
rlabel metal1 31970 17136 31970 17136 0 _0245_
rlabel metal1 32154 17102 32154 17102 0 _0246_
rlabel metal1 32338 17204 32338 17204 0 _0247_
rlabel metal1 18078 16660 18078 16660 0 _0248_
rlabel metal1 24564 19482 24564 19482 0 _0249_
rlabel metal1 28704 25466 28704 25466 0 _0250_
rlabel metal1 18262 22542 18262 22542 0 _0251_
rlabel metal1 27646 37740 27646 37740 0 _0252_
rlabel metal1 29854 37876 29854 37876 0 _0253_
rlabel metal1 26956 37842 26956 37842 0 _0254_
rlabel metal1 27968 32878 27968 32878 0 _0255_
rlabel metal1 28980 28186 28980 28186 0 _0256_
rlabel metal1 28612 29818 28612 29818 0 _0257_
rlabel metal1 27600 26010 27600 26010 0 _0258_
rlabel metal1 26772 34170 26772 34170 0 _0259_
rlabel metal1 28474 24378 28474 24378 0 _0260_
rlabel metal1 14490 17510 14490 17510 0 _0261_
rlabel metal1 9430 20400 9430 20400 0 _0262_
rlabel metal1 9246 20366 9246 20366 0 _0263_
rlabel metal1 12650 21114 12650 21114 0 _0264_
rlabel metal1 13662 24786 13662 24786 0 _0265_
rlabel metal1 13156 23630 13156 23630 0 _0266_
rlabel metal2 13386 24021 13386 24021 0 _0267_
rlabel metal1 13294 24650 13294 24650 0 _0268_
rlabel viali 13662 24169 13662 24169 0 _0269_
rlabel metal1 8418 35564 8418 35564 0 _0270_
rlabel metal1 9338 37230 9338 37230 0 _0271_
rlabel metal1 10166 35598 10166 35598 0 _0272_
rlabel metal1 10580 37842 10580 37842 0 _0273_
rlabel metal1 8924 21658 8924 21658 0 _0274_
rlabel metal1 7820 32878 7820 32878 0 _0275_
rlabel metal1 8142 27540 8142 27540 0 _0276_
rlabel metal1 7544 27438 7544 27438 0 _0277_
rlabel metal1 9706 21114 9706 21114 0 _0278_
rlabel metal1 10442 30702 10442 30702 0 _0279_
rlabel metal1 11454 24038 11454 24038 0 _0280_
rlabel metal1 11500 27642 11500 27642 0 _0281_
rlabel metal1 9568 20570 9568 20570 0 _0282_
rlabel metal1 7774 35666 7774 35666 0 _0283_
rlabel metal1 10810 21930 10810 21930 0 _0284_
rlabel metal1 9752 24922 9752 24922 0 _0285_
rlabel metal1 12696 24310 12696 24310 0 _0286_
rlabel metal1 13478 25228 13478 25228 0 _0287_
rlabel metal1 13892 25262 13892 25262 0 _0288_
rlabel metal1 33672 34034 33672 34034 0 _0289_
rlabel metal2 32338 37502 32338 37502 0 _0290_
rlabel metal1 25760 37842 25760 37842 0 _0291_
rlabel metal1 34270 34034 34270 34034 0 _0292_
rlabel metal1 33396 27914 33396 27914 0 _0293_
rlabel metal1 34224 30362 34224 30362 0 _0294_
rlabel metal1 27232 27642 27232 27642 0 _0295_
rlabel metal1 30820 35258 30820 35258 0 _0296_
rlabel metal1 24564 25466 24564 25466 0 _0297_
rlabel metal1 13386 37774 13386 37774 0 _0298_
rlabel metal1 20332 37978 20332 37978 0 _0299_
rlabel metal2 12742 38454 12742 38454 0 _0300_
rlabel metal1 5106 31280 5106 31280 0 _0301_
rlabel metal1 5198 27438 5198 27438 0 _0302_
rlabel metal1 8464 31858 8464 31858 0 _0303_
rlabel metal2 10994 27132 10994 27132 0 _0304_
rlabel metal1 5888 35258 5888 35258 0 _0305_
rlabel metal1 6210 26010 6210 26010 0 _0306_
rlabel metal1 14582 24344 14582 24344 0 _0307_
rlabel metal2 17158 24565 17158 24565 0 _0308_
rlabel metal1 32890 35802 32890 35802 0 _0309_
rlabel metal1 27370 35802 27370 35802 0 _0310_
rlabel metal1 33902 32946 33902 32946 0 _0311_
rlabel metal1 32062 28050 32062 28050 0 _0312_
rlabel metal1 32246 29002 32246 29002 0 _0313_
rlabel metal1 32062 25874 32062 25874 0 _0314_
rlabel metal1 30912 34578 30912 34578 0 _0315_
rlabel metal2 24886 23698 24886 23698 0 _0316_
rlabel metal1 6532 32946 6532 32946 0 _0317_
rlabel metal1 11178 35666 11178 35666 0 _0318_
rlabel metal1 9660 35666 9660 35666 0 _0319_
rlabel metal1 5566 32878 5566 32878 0 _0320_
rlabel metal1 5198 28560 5198 28560 0 _0321_
rlabel metal1 11224 32402 11224 32402 0 _0322_
rlabel metal1 9338 26350 9338 26350 0 _0323_
rlabel metal1 5980 33966 5980 33966 0 _0324_
rlabel metal1 6624 25466 6624 25466 0 _0325_
rlabel metal3 12420 19312 12420 19312 0 _0326_
rlabel metal1 15042 19380 15042 19380 0 _0327_
rlabel metal2 9844 33524 9844 33524 0 _0328_
rlabel metal1 15594 17034 15594 17034 0 _0329_
rlabel metal2 15778 17850 15778 17850 0 _0330_
rlabel metal1 15180 17170 15180 17170 0 _0331_
rlabel metal2 14398 16796 14398 16796 0 _0332_
rlabel metal1 13662 16422 13662 16422 0 _0333_
rlabel metal2 13386 19652 13386 19652 0 _0334_
rlabel metal1 12650 17238 12650 17238 0 _0335_
rlabel metal1 8970 33966 8970 33966 0 _0336_
rlabel metal1 10350 30022 10350 30022 0 _0337_
rlabel metal1 24518 19958 24518 19958 0 _0338_
rlabel metal1 23828 20026 23828 20026 0 _0339_
rlabel metal2 23782 19652 23782 19652 0 _0340_
rlabel metal1 22816 18666 22816 18666 0 _0341_
rlabel metal2 23690 19720 23690 19720 0 _0342_
rlabel metal2 12190 19635 12190 19635 0 _0343_
rlabel metal1 10580 23834 10580 23834 0 _0344_
rlabel metal1 10166 28458 10166 28458 0 _0345_
rlabel metal2 33350 17850 33350 17850 0 _0346_
rlabel metal1 29026 14960 29026 14960 0 _0347_
rlabel metal1 30222 7820 30222 7820 0 _0348_
rlabel metal1 33350 7446 33350 7446 0 _0349_
rlabel metal1 24426 5882 24426 5882 0 _0350_
rlabel metal1 24935 6426 24935 6426 0 _0351_
rlabel metal1 24242 7412 24242 7412 0 _0352_
rlabel metal1 25024 6834 25024 6834 0 _0353_
rlabel metal2 33350 6664 33350 6664 0 _0354_
rlabel metal2 33718 9078 33718 9078 0 _0355_
rlabel metal1 33902 9962 33902 9962 0 _0356_
rlabel metal1 34592 10166 34592 10166 0 _0357_
rlabel metal1 24610 10200 24610 10200 0 _0358_
rlabel metal1 34914 10234 34914 10234 0 _0359_
rlabel metal2 34868 11220 34868 11220 0 _0360_
rlabel metal1 34960 16762 34960 16762 0 _0361_
rlabel metal1 32890 20774 32890 20774 0 _0362_
rlabel metal1 33718 17816 33718 17816 0 _0363_
rlabel metal1 33902 17646 33902 17646 0 _0364_
rlabel metal1 34132 17306 34132 17306 0 _0365_
rlabel metal1 34362 17170 34362 17170 0 _0366_
rlabel metal1 29854 15062 29854 15062 0 _0367_
rlabel metal1 31234 14416 31234 14416 0 _0368_
rlabel metal1 32016 14586 32016 14586 0 _0369_
rlabel metal1 32752 15538 32752 15538 0 _0370_
rlabel metal1 33626 15674 33626 15674 0 _0371_
rlabel metal1 33994 17136 33994 17136 0 _0372_
rlabel metal1 34730 16966 34730 16966 0 _0373_
rlabel metal1 34822 17204 34822 17204 0 _0374_
rlabel metal1 30912 16966 30912 16966 0 _0375_
rlabel metal1 29264 17238 29264 17238 0 _0376_
rlabel metal2 29164 8908 29164 8908 0 _0377_
rlabel metal2 28014 17340 28014 17340 0 _0378_
rlabel metal2 29486 17510 29486 17510 0 _0379_
rlabel metal1 23690 17102 23690 17102 0 _0380_
rlabel metal1 24426 17306 24426 17306 0 _0381_
rlabel metal1 24334 17714 24334 17714 0 _0382_
rlabel metal1 26082 17612 26082 17612 0 _0383_
rlabel metal1 25898 17714 25898 17714 0 _0384_
rlabel metal1 26634 17748 26634 17748 0 _0385_
rlabel metal1 27186 17646 27186 17646 0 _0386_
rlabel metal1 28842 17612 28842 17612 0 _0387_
rlabel metal1 12144 18190 12144 18190 0 _0388_
rlabel metal1 11684 24378 11684 24378 0 _0389_
rlabel metal1 11040 25466 11040 25466 0 _0390_
rlabel metal1 10396 32946 10396 32946 0 _0391_
rlabel metal1 30038 16116 30038 16116 0 _0392_
rlabel metal2 30130 17204 30130 17204 0 _0393_
rlabel metal1 29348 11866 29348 11866 0 _0394_
rlabel metal1 23322 12274 23322 12274 0 _0395_
rlabel metal2 25990 12087 25990 12087 0 _0396_
rlabel metal1 25254 11526 25254 11526 0 _0397_
rlabel metal1 28750 12410 28750 12410 0 _0398_
rlabel metal2 28382 17748 28382 17748 0 _0399_
rlabel metal1 28244 19346 28244 19346 0 _0400_
rlabel metal1 28474 19278 28474 19278 0 _0401_
rlabel metal1 28749 19346 28749 19346 0 _0402_
rlabel metal1 28934 18292 28934 18292 0 _0403_
rlabel metal2 11362 20591 11362 20591 0 _0404_
rlabel metal1 11454 22202 11454 22202 0 _0405_
rlabel metal2 11546 23188 11546 23188 0 _0406_
rlabel metal1 8188 19890 8188 19890 0 _0407_
rlabel metal1 12236 6358 12236 6358 0 _0408_
rlabel metal2 12834 7684 12834 7684 0 _0409_
rlabel metal1 13202 5610 13202 5610 0 _0410_
rlabel metal1 16100 12682 16100 12682 0 _0411_
rlabel metal2 13202 6596 13202 6596 0 _0412_
rlabel metal2 12834 16932 12834 16932 0 _0413_
rlabel metal1 8832 5610 8832 5610 0 _0414_
rlabel metal2 9430 5984 9430 5984 0 _0415_
rlabel metal2 8694 4998 8694 4998 0 _0416_
rlabel metal1 12489 19822 12489 19822 0 _0417_
rlabel metal1 12696 19686 12696 19686 0 _0418_
rlabel metal1 8142 10030 8142 10030 0 _0419_
rlabel metal1 8970 12206 8970 12206 0 _0420_
rlabel metal2 9246 12002 9246 12002 0 _0421_
rlabel metal2 9384 13158 9384 13158 0 _0422_
rlabel metal1 10074 12172 10074 12172 0 _0423_
rlabel metal1 9522 12206 9522 12206 0 _0424_
rlabel metal2 8050 10744 8050 10744 0 _0425_
rlabel metal1 14214 10778 14214 10778 0 _0426_
rlabel metal1 9108 9894 9108 9894 0 _0427_
rlabel metal1 9016 11526 9016 11526 0 _0428_
rlabel metal1 12926 9554 12926 9554 0 _0429_
rlabel metal2 8234 9180 8234 9180 0 _0430_
rlabel metal2 8602 7888 8602 7888 0 _0431_
rlabel metal1 8142 6324 8142 6324 0 _0432_
rlabel metal1 8970 12614 8970 12614 0 _0433_
rlabel metal1 8372 10234 8372 10234 0 _0434_
rlabel metal1 14812 8942 14812 8942 0 _0435_
rlabel metal2 15318 9792 15318 9792 0 _0436_
rlabel metal1 8878 10098 8878 10098 0 _0437_
rlabel metal1 8326 6834 8326 6834 0 _0438_
rlabel metal1 8464 5202 8464 5202 0 _0439_
rlabel metal1 6670 18122 6670 18122 0 _0440_
rlabel metal1 13984 18734 13984 18734 0 _0441_
rlabel metal2 12650 20893 12650 20893 0 _0442_
rlabel metal1 15042 5644 15042 5644 0 _0443_
rlabel metal2 14490 5474 14490 5474 0 _0444_
rlabel metal1 2530 18700 2530 18700 0 _0445_
rlabel metal1 16468 3026 16468 3026 0 _0446_
rlabel metal2 37582 33286 37582 33286 0 _0447_
rlabel metal1 37030 3026 37030 3026 0 _0448_
rlabel metal2 12558 31586 12558 31586 0 _0449_
rlabel via3 11845 4012 11845 4012 0 _0450_
rlabel metal3 13271 4012 13271 4012 0 _0451_
rlabel metal1 1978 28594 1978 28594 0 _0452_
rlabel metal1 37444 23086 37444 23086 0 _0453_
rlabel metal1 2162 18938 2162 18938 0 _0454_
rlabel metal1 8050 8398 8050 8398 0 _0455_
rlabel metal1 9476 8602 9476 8602 0 _0456_
rlabel metal1 5106 9146 5106 9146 0 _0457_
rlabel metal1 3082 8500 3082 8500 0 _0458_
rlabel metal1 13478 10540 13478 10540 0 _0459_
rlabel metal2 2990 10540 2990 10540 0 _0460_
rlabel metal1 5796 15130 5796 15130 0 _0461_
rlabel metal1 3956 18394 3956 18394 0 _0462_
rlabel via2 7498 17731 7498 17731 0 _0463_
rlabel metal2 17618 14421 17618 14421 0 _0464_
rlabel metal1 17664 3026 17664 3026 0 _0465_
rlabel metal1 2484 19346 2484 19346 0 _0466_
rlabel metal1 1794 18292 1794 18292 0 _0467_
rlabel metal1 2530 21658 2530 21658 0 _0468_
rlabel metal3 17204 21896 17204 21896 0 _0469_
rlabel via2 9338 22083 9338 22083 0 _0470_
rlabel metal1 12742 22032 12742 22032 0 _0471_
rlabel metal1 5750 20944 5750 20944 0 _0472_
rlabel metal1 5474 18394 5474 18394 0 _0473_
rlabel metal1 2461 18258 2461 18258 0 _0474_
rlabel metal1 26082 21488 26082 21488 0 _0475_
rlabel metal1 26542 21998 26542 21998 0 _0476_
rlabel metal1 25024 37434 25024 37434 0 _0477_
rlabel metal2 2254 20519 2254 20519 0 _0478_
rlabel metal1 37398 20978 37398 20978 0 _0479_
rlabel metal2 25346 16932 25346 16932 0 _0480_
rlabel metal2 34546 37774 34546 37774 0 _0481_
rlabel metal2 32062 38012 32062 38012 0 _0482_
rlabel metal2 5198 38369 5198 38369 0 _0483_
rlabel via2 11730 37859 11730 37859 0 _0484_
rlabel metal1 13800 4590 13800 4590 0 _0485_
rlabel metal1 7038 6324 7038 6324 0 _0486_
rlabel metal1 5474 13974 5474 13974 0 _0487_
rlabel metal1 6164 12818 6164 12818 0 _0488_
rlabel metal1 6440 11322 6440 11322 0 _0489_
rlabel metal2 9338 19584 9338 19584 0 _0490_
rlabel metal1 7682 19822 7682 19822 0 _0491_
rlabel metal1 7682 16082 7682 16082 0 _0492_
rlabel metal1 6854 14382 6854 14382 0 _0493_
rlabel metal1 6532 9690 6532 9690 0 _0494_
rlabel metal1 7636 17850 7636 17850 0 _0495_
rlabel metal2 11914 7548 11914 7548 0 _0496_
rlabel metal2 13294 8092 13294 8092 0 _0497_
rlabel metal1 15594 11186 15594 11186 0 _0498_
rlabel metal1 15456 11730 15456 11730 0 _0499_
rlabel metal1 16146 8466 16146 8466 0 _0500_
rlabel metal1 10580 12818 10580 12818 0 _0501_
rlabel metal1 9154 15130 9154 15130 0 _0502_
rlabel metal1 12972 12206 12972 12206 0 _0503_
rlabel metal1 13754 7922 13754 7922 0 _0504_
rlabel metal1 12558 13906 12558 13906 0 _0505_
rlabel metal1 14858 10030 14858 10030 0 _0506_
rlabel metal2 15226 6970 15226 6970 0 _0507_
rlabel metal2 14306 8262 14306 8262 0 _0508_
rlabel metal1 10442 9690 10442 9690 0 _0509_
rlabel metal1 8694 13294 8694 13294 0 _0510_
rlabel metal1 12006 10710 12006 10710 0 _0511_
rlabel metal1 12328 9554 12328 9554 0 _0512_
rlabel metal1 11316 14994 11316 14994 0 _0513_
rlabel metal1 29992 30634 29992 30634 0 _0514_
rlabel metal2 17986 30736 17986 30736 0 _0515_
rlabel metal2 19458 30736 19458 30736 0 _0516_
rlabel metal1 29578 31416 29578 31416 0 _0517_
rlabel metal1 17664 15674 17664 15674 0 _0518_
rlabel metal1 14766 9486 14766 9486 0 _0519_
rlabel metal1 14536 10030 14536 10030 0 _0520_
rlabel metal1 14306 9962 14306 9962 0 _0521_
rlabel metal1 13271 10166 13271 10166 0 _0522_
rlabel metal1 10488 18190 10488 18190 0 _0523_
rlabel metal1 11822 17544 11822 17544 0 _0524_
rlabel via1 11546 19278 11546 19278 0 _0525_
rlabel metal1 11086 18224 11086 18224 0 _0526_
rlabel metal1 11546 17306 11546 17306 0 _0527_
rlabel metal1 11224 17306 11224 17306 0 _0528_
rlabel metal1 10258 17850 10258 17850 0 _0529_
rlabel metal1 11040 19414 11040 19414 0 _0530_
rlabel metal2 11822 18292 11822 18292 0 _0531_
rlabel viali 10902 18735 10902 18735 0 _0532_
rlabel metal1 10534 18360 10534 18360 0 _0533_
rlabel metal1 9936 18122 9936 18122 0 _0534_
rlabel metal1 10718 18360 10718 18360 0 _0535_
rlabel metal2 12742 18496 12742 18496 0 _0536_
rlabel metal1 11362 18122 11362 18122 0 _0537_
rlabel metal1 11316 17646 11316 17646 0 _0538_
rlabel metal1 9982 17714 9982 17714 0 _0539_
rlabel metal1 7130 22678 7130 22678 0 _0540_
rlabel metal1 7406 8602 7406 8602 0 _0541_
rlabel metal2 3082 19584 3082 19584 0 _0542_
rlabel metal1 6624 7378 6624 7378 0 _0543_
rlabel metal1 17250 7480 17250 7480 0 _0544_
rlabel metal2 17250 7072 17250 7072 0 _0545_
rlabel metal1 5198 7514 5198 7514 0 _0546_
rlabel metal1 4692 7514 4692 7514 0 _0547_
rlabel metal1 3680 6766 3680 6766 0 _0548_
rlabel metal2 13846 8976 13846 8976 0 _0549_
rlabel metal1 5428 8942 5428 8942 0 _0550_
rlabel metal1 5014 8942 5014 8942 0 _0551_
rlabel metal1 4462 9044 4462 9044 0 _0552_
rlabel metal1 2806 9044 2806 9044 0 _0553_
rlabel metal1 2254 8942 2254 8942 0 _0554_
rlabel metal1 9246 10540 9246 10540 0 _0555_
rlabel metal1 4370 13294 4370 13294 0 _0556_
rlabel metal1 4784 10234 4784 10234 0 _0557_
rlabel metal1 4922 10778 4922 10778 0 _0558_
rlabel metal2 4646 10880 4646 10880 0 _0559_
rlabel metal1 3634 11118 3634 11118 0 _0560_
rlabel metal1 5060 12954 5060 12954 0 _0561_
rlabel metal1 4094 12750 4094 12750 0 _0562_
rlabel metal1 3312 12206 3312 12206 0 _0563_
rlabel metal1 2116 12206 2116 12206 0 _0564_
rlabel metal1 12972 13362 12972 13362 0 _0565_
rlabel metal2 11178 13770 11178 13770 0 _0566_
rlabel metal1 4094 14348 4094 14348 0 _0567_
rlabel metal1 3864 14382 3864 14382 0 _0568_
rlabel metal1 4048 14042 4048 14042 0 _0569_
rlabel metal2 2990 13566 2990 13566 0 _0570_
rlabel metal1 2346 13294 2346 13294 0 _0571_
rlabel metal1 5520 15470 5520 15470 0 _0572_
rlabel metal1 4646 16660 4646 16660 0 _0573_
rlabel metal1 4370 16116 4370 16116 0 _0574_
rlabel metal1 4278 15572 4278 15572 0 _0575_
rlabel metal1 3450 15130 3450 15130 0 _0576_
rlabel metal1 2392 14994 2392 14994 0 _0577_
rlabel metal1 12535 15946 12535 15946 0 _0578_
rlabel metal1 5704 16626 5704 16626 0 _0579_
rlabel metal2 5842 16898 5842 16898 0 _0580_
rlabel metal1 5336 17170 5336 17170 0 _0581_
rlabel viali 4554 17651 4554 17651 0 _0582_
rlabel metal1 4094 17544 4094 17544 0 _0583_
rlabel metal1 3956 17102 3956 17102 0 _0584_
rlabel metal1 5776 22066 5776 22066 0 _0585_
rlabel metal1 3404 17510 3404 17510 0 _0586_
rlabel metal2 2530 17136 2530 17136 0 _0587_
rlabel via2 4094 22627 4094 22627 0 _0588_
rlabel metal2 3726 20604 3726 20604 0 _0589_
rlabel metal1 3634 20366 3634 20366 0 _0590_
rlabel metal1 3220 20570 3220 20570 0 _0591_
rlabel metal1 2530 20502 2530 20502 0 _0592_
rlabel metal1 3404 22678 3404 22678 0 _0593_
rlabel metal1 4232 22746 4232 22746 0 _0594_
rlabel metal1 3358 23290 3358 23290 0 _0595_
rlabel metal1 2392 24786 2392 24786 0 _0596_
rlabel viali 8237 22610 8237 22610 0 _0597_
rlabel metal1 3634 22542 3634 22542 0 _0598_
rlabel metal1 3680 22202 3680 22202 0 _0599_
rlabel metal1 3082 22746 3082 22746 0 _0600_
rlabel metal1 2162 23086 2162 23086 0 _0601_
rlabel metal2 8326 22882 8326 22882 0 _0602_
rlabel viali 8237 23086 8237 23086 0 _0603_
rlabel metal1 7866 23290 7866 23290 0 _0604_
rlabel metal1 7176 23698 7176 23698 0 _0605_
rlabel metal2 6026 21760 6026 21760 0 _0606_
rlabel metal1 7268 22134 7268 22134 0 _0607_
rlabel metal1 6854 22576 6854 22576 0 _0608_
rlabel metal1 6716 22610 6716 22610 0 _0609_
rlabel metal1 5566 22678 5566 22678 0 _0610_
rlabel metal2 5750 20604 5750 20604 0 _0611_
rlabel metal1 5474 21930 5474 21930 0 _0612_
rlabel metal1 5106 22066 5106 22066 0 _0613_
rlabel metal1 4324 24174 4324 24174 0 _0614_
rlabel metal1 6302 19414 6302 19414 0 _0615_
rlabel metal1 5934 18836 5934 18836 0 _0616_
rlabel metal1 5244 18734 5244 18734 0 _0617_
rlabel metal1 15594 17578 15594 17578 0 _0618_
rlabel metal1 20102 20842 20102 20842 0 _0619_
rlabel via1 20104 17170 20104 17170 0 _0620_
rlabel metal1 20746 18326 20746 18326 0 _0621_
rlabel metal1 20608 19822 20608 19822 0 _0622_
rlabel metal1 15180 21998 15180 21998 0 _0623_
rlabel metal1 18906 19822 18906 19822 0 _0624_
rlabel metal1 14766 15130 14766 15130 0 _0625_
rlabel metal2 17158 22039 17158 22039 0 _0626_
rlabel metal1 14168 14586 14168 14586 0 _0627_
rlabel metal2 15042 16592 15042 16592 0 _0628_
rlabel metal1 15134 26996 15134 26996 0 _0629_
rlabel via2 16606 19499 16606 19499 0 _0630_
rlabel metal1 24288 20910 24288 20910 0 _0631_
rlabel metal1 15502 14348 15502 14348 0 _0632_
rlabel metal1 16744 20502 16744 20502 0 _0633_
rlabel metal2 17342 21284 17342 21284 0 _0634_
rlabel metal1 18262 13872 18262 13872 0 _0635_
rlabel metal1 14168 18938 14168 18938 0 _0636_
rlabel via1 17801 20910 17801 20910 0 _0637_
rlabel metal1 18722 21590 18722 21590 0 _0638_
rlabel metal1 14996 16082 14996 16082 0 _0639_
rlabel metal2 18906 19346 18906 19346 0 _0640_
rlabel metal1 19596 19346 19596 19346 0 _0641_
rlabel metal1 16422 19822 16422 19822 0 _0642_
rlabel metal2 18722 18870 18722 18870 0 _0643_
rlabel metal1 19550 20911 19550 20911 0 _0644_
rlabel metal1 20424 16082 20424 16082 0 _0645_
rlabel metal1 21528 21998 21528 21998 0 _0646_
rlabel metal2 19918 17119 19918 17119 0 _0647_
rlabel metal1 14582 17714 14582 17714 0 _0648_
rlabel metal2 20654 19312 20654 19312 0 _0649_
rlabel metal1 21620 20910 21620 20910 0 _0650_
rlabel metal1 23782 23732 23782 23732 0 _0651_
rlabel metal2 28750 24106 28750 24106 0 _0652_
rlabel metal1 15272 21658 15272 21658 0 _0653_
rlabel metal2 15778 23426 15778 23426 0 _0654_
rlabel metal1 13156 19754 13156 19754 0 _0655_
rlabel metal1 17112 13294 17112 13294 0 _0656_
rlabel metal1 17894 13498 17894 13498 0 _0657_
rlabel metal2 11638 6086 11638 6086 0 _0658_
rlabel metal1 14582 12614 14582 12614 0 _0659_
rlabel metal1 16514 14382 16514 14382 0 _0660_
rlabel metal2 16238 15504 16238 15504 0 _0661_
rlabel metal2 16146 14076 16146 14076 0 _0662_
rlabel metal1 16928 14042 16928 14042 0 _0663_
rlabel metal1 18814 14382 18814 14382 0 _0664_
rlabel metal1 15548 20910 15548 20910 0 _0665_
rlabel metal1 17986 15028 17986 15028 0 _0666_
rlabel metal1 17066 17306 17066 17306 0 _0667_
rlabel metal1 16330 17204 16330 17204 0 _0668_
rlabel metal1 17250 16116 17250 16116 0 _0669_
rlabel metal1 16146 16014 16146 16014 0 _0670_
rlabel metal1 17342 16048 17342 16048 0 _0671_
rlabel metal1 17434 16014 17434 16014 0 _0672_
rlabel metal1 17342 14994 17342 14994 0 _0673_
rlabel metal1 18630 10642 18630 10642 0 _0674_
rlabel metal1 19734 8432 19734 8432 0 _0675_
rlabel metal2 30728 29614 30728 29614 0 _0676_
rlabel metal2 18998 21692 18998 21692 0 _0677_
rlabel metal2 20930 15572 20930 15572 0 _0678_
rlabel metal1 18952 22066 18952 22066 0 _0679_
rlabel metal1 13570 27438 13570 27438 0 _0680_
rlabel metal1 19504 21658 19504 21658 0 _0681_
rlabel metal2 14306 37536 14306 37536 0 _0682_
rlabel metal1 22494 35122 22494 35122 0 _0683_
rlabel metal1 21850 21998 21850 21998 0 _0684_
rlabel metal1 12972 27370 12972 27370 0 _0685_
rlabel metal1 18262 23290 18262 23290 0 _0686_
rlabel metal1 13018 32810 13018 32810 0 _0687_
rlabel metal1 27186 35054 27186 35054 0 _0688_
rlabel metal2 28290 33218 28290 33218 0 _0689_
rlabel metal1 28934 22576 28934 22576 0 _0690_
rlabel metal2 29210 21801 29210 21801 0 _0691_
rlabel metal1 18630 14280 18630 14280 0 _0692_
rlabel metal1 20056 16558 20056 16558 0 _0693_
rlabel metal1 16606 23086 16606 23086 0 _0694_
rlabel metal2 17526 18938 17526 18938 0 _0695_
rlabel metal1 17020 18394 17020 18394 0 _0696_
rlabel metal1 15088 18598 15088 18598 0 _0697_
rlabel metal1 16928 18802 16928 18802 0 _0698_
rlabel metal1 19826 32402 19826 32402 0 _0699_
rlabel metal2 19642 14688 19642 14688 0 _0700_
rlabel metal1 17296 21658 17296 21658 0 _0701_
rlabel metal1 16606 17850 16606 17850 0 _0702_
rlabel metal1 17296 24038 17296 24038 0 _0703_
rlabel metal1 18124 25874 18124 25874 0 _0704_
rlabel metal2 17894 27948 17894 27948 0 _0705_
rlabel metal1 16974 25262 16974 25262 0 _0706_
rlabel metal2 17434 34782 17434 34782 0 _0707_
rlabel metal2 20378 33184 20378 33184 0 _0708_
rlabel metal1 25162 24854 25162 24854 0 _0709_
rlabel viali 25430 36142 25430 36142 0 _0710_
rlabel metal1 19826 26350 19826 26350 0 _0711_
rlabel metal2 25162 35530 25162 35530 0 _0712_
rlabel metal1 24748 34918 24748 34918 0 _0713_
rlabel metal1 28750 22644 28750 22644 0 _0714_
rlabel metal1 29716 20366 29716 20366 0 _0715_
rlabel metal1 29532 21998 29532 21998 0 _0716_
rlabel metal1 29302 22644 29302 22644 0 _0717_
rlabel metal2 29762 22202 29762 22202 0 _0718_
rlabel metal1 30590 29818 30590 29818 0 _0719_
rlabel metal1 30498 29648 30498 29648 0 _0720_
rlabel metal1 33902 24786 33902 24786 0 _0721_
rlabel metal1 25806 29648 25806 29648 0 _0722_
rlabel metal2 25530 29308 25530 29308 0 _0723_
rlabel metal1 25070 21454 25070 21454 0 _0724_
rlabel metal1 34638 23630 34638 23630 0 _0725_
rlabel metal1 34684 22746 34684 22746 0 _0726_
rlabel metal1 29716 26350 29716 26350 0 _0727_
rlabel metal1 31188 26350 31188 26350 0 _0728_
rlabel metal1 34040 24106 34040 24106 0 _0729_
rlabel metal1 26220 25874 26220 25874 0 _0730_
rlabel metal1 25852 26010 25852 26010 0 _0731_
rlabel metal1 26956 22066 26956 22066 0 _0732_
rlabel metal1 27554 22440 27554 22440 0 _0733_
rlabel metal1 35696 22066 35696 22066 0 _0734_
rlabel metal1 35834 22610 35834 22610 0 _0735_
rlabel metal1 35098 21930 35098 21930 0 _0736_
rlabel metal1 35374 20978 35374 20978 0 _0737_
rlabel metal1 29900 33966 29900 33966 0 _0738_
rlabel metal1 30636 31790 30636 31790 0 _0739_
rlabel metal1 33304 19822 33304 19822 0 _0740_
rlabel metal1 24426 33626 24426 33626 0 _0741_
rlabel metal2 25714 34170 25714 34170 0 _0742_
rlabel metal1 25116 34170 25116 34170 0 _0743_
rlabel metal2 25070 23579 25070 23579 0 _0744_
rlabel metal1 33626 19958 33626 19958 0 _0745_
rlabel metal1 35098 19856 35098 19856 0 _0746_
rlabel metal1 26588 24378 26588 24378 0 _0747_
rlabel metal2 30682 24378 30682 24378 0 _0748_
rlabel metal1 31602 19380 31602 19380 0 _0749_
rlabel metal1 26082 24684 26082 24684 0 _0750_
rlabel metal1 25806 25228 25806 25228 0 _0751_
rlabel metal3 25093 34476 25093 34476 0 _0752_
rlabel metal2 31970 19006 31970 19006 0 _0753_
rlabel metal1 32062 18666 32062 18666 0 _0754_
rlabel metal1 31740 18734 31740 18734 0 _0755_
rlabel metal1 32706 19380 32706 19380 0 _0756_
rlabel metal2 20746 19414 20746 19414 0 _0757_
rlabel metal1 20608 20026 20608 20026 0 _0758_
rlabel metal1 20838 20400 20838 20400 0 _0759_
rlabel metal1 14950 35054 14950 35054 0 _0760_
rlabel metal1 20838 22066 20838 22066 0 _0761_
rlabel metal2 14582 28169 14582 28169 0 _0762_
rlabel metal1 23322 27302 23322 27302 0 _0763_
rlabel metal1 23552 31994 23552 31994 0 _0764_
rlabel metal2 18078 35632 18078 35632 0 _0765_
rlabel metal1 22172 21998 22172 21998 0 _0766_
rlabel metal1 15502 33966 15502 33966 0 _0767_
rlabel metal1 22908 32878 22908 32878 0 _0768_
rlabel viali 23230 32403 23230 32403 0 _0769_
rlabel metal2 21666 25976 21666 25976 0 _0770_
rlabel metal2 15962 27115 15962 27115 0 _0771_
rlabel metal1 21988 21386 21988 21386 0 _0772_
rlabel metal1 23322 32300 23322 32300 0 _0773_
rlabel metal1 15916 26962 15916 26962 0 _0774_
rlabel metal2 13846 19635 13846 19635 0 _0775_
rlabel metal1 13156 31790 13156 31790 0 _0776_
rlabel metal2 12834 32266 12834 32266 0 _0777_
rlabel metal1 13432 19346 13432 19346 0 _0778_
rlabel metal1 19090 11050 19090 11050 0 _0779_
rlabel metal1 23276 19346 23276 19346 0 _0780_
rlabel metal1 33212 11662 33212 11662 0 _0781_
rlabel metal2 27186 11424 27186 11424 0 _0782_
rlabel metal1 18170 24106 18170 24106 0 _0783_
rlabel metal1 18078 30702 18078 30702 0 _0784_
rlabel metal1 17664 20026 17664 20026 0 _0785_
rlabel metal2 17526 38216 17526 38216 0 _0786_
rlabel metal1 24058 32198 24058 32198 0 _0787_
rlabel metal1 20148 34646 20148 34646 0 _0788_
rlabel metal2 16560 33966 16560 33966 0 _0789_
rlabel metal1 22862 31382 22862 31382 0 _0790_
rlabel metal1 23552 30838 23552 30838 0 _0791_
rlabel metal1 18492 25670 18492 25670 0 _0792_
rlabel metal1 18124 36142 18124 36142 0 _0793_
rlabel metal1 22908 25942 22908 25942 0 _0794_
rlabel metal1 21850 32470 21850 32470 0 _0795_
rlabel metal2 23966 30804 23966 30804 0 _0796_
rlabel metal1 24058 30736 24058 30736 0 _0797_
rlabel metal1 24794 30668 24794 30668 0 _0798_
rlabel metal1 21482 32198 21482 32198 0 _0799_
rlabel metal1 21390 31654 21390 31654 0 _0800_
rlabel metal1 25254 30804 25254 30804 0 _0801_
rlabel metal1 27554 11152 27554 11152 0 _0802_
rlabel metal1 33350 11764 33350 11764 0 _0803_
rlabel metal1 33304 11866 33304 11866 0 _0804_
rlabel metal1 34086 13328 34086 13328 0 _0805_
rlabel metal1 33212 10642 33212 10642 0 _0806_
rlabel metal1 14904 27574 14904 27574 0 _0807_
rlabel metal1 14996 27914 14996 27914 0 _0808_
rlabel metal1 15364 26962 15364 26962 0 _0809_
rlabel metal1 15594 26792 15594 26792 0 _0810_
rlabel metal2 15686 27132 15686 27132 0 _0811_
rlabel metal1 15042 26928 15042 26928 0 _0812_
rlabel metal1 14030 26826 14030 26826 0 _0813_
rlabel metal1 14168 26962 14168 26962 0 _0814_
rlabel metal1 14306 9452 14306 9452 0 _0815_
rlabel metal2 22494 7650 22494 7650 0 _0816_
rlabel metal1 21758 29478 21758 29478 0 _0817_
rlabel metal1 16928 26350 16928 26350 0 _0818_
rlabel metal1 17894 26452 17894 26452 0 _0819_
rlabel viali 18998 26961 18998 26961 0 _0820_
rlabel metal1 18630 26554 18630 26554 0 _0821_
rlabel metal2 17802 27234 17802 27234 0 _0822_
rlabel metal1 18354 25194 18354 25194 0 _0823_
rlabel metal1 18538 25262 18538 25262 0 _0824_
rlabel metal2 16698 27268 16698 27268 0 _0825_
rlabel metal2 18078 26044 18078 26044 0 _0826_
rlabel metal1 18170 24718 18170 24718 0 _0827_
rlabel metal1 19044 14586 19044 14586 0 _0828_
rlabel metal2 17894 10268 17894 10268 0 _0829_
rlabel metal1 17894 10030 17894 10030 0 _0830_
rlabel metal2 20332 9996 20332 9996 0 _0831_
rlabel metal2 25622 4692 25622 4692 0 _0832_
rlabel metal1 16928 29818 16928 29818 0 _0833_
rlabel metal1 18400 30090 18400 30090 0 _0834_
rlabel metal1 17802 30702 17802 30702 0 _0835_
rlabel metal1 18722 30906 18722 30906 0 _0836_
rlabel metal1 19136 30702 19136 30702 0 _0837_
rlabel viali 18356 29137 18356 29137 0 _0838_
rlabel viali 18262 29138 18262 29138 0 _0839_
rlabel metal1 16698 30668 16698 30668 0 _0840_
rlabel metal1 18492 29614 18492 29614 0 _0841_
rlabel metal1 18630 29206 18630 29206 0 _0842_
rlabel metal3 18561 10948 18561 10948 0 _0843_
rlabel metal1 19090 10200 19090 10200 0 _0844_
rlabel metal1 15226 30294 15226 30294 0 _0845_
rlabel metal2 14950 31212 14950 31212 0 _0846_
rlabel metal1 14720 29614 14720 29614 0 _0847_
rlabel metal1 15594 29750 15594 29750 0 _0848_
rlabel metal1 15318 29682 15318 29682 0 _0849_
rlabel metal1 14260 29682 14260 29682 0 _0850_
rlabel metal1 13248 29614 13248 29614 0 _0851_
rlabel metal2 13662 30090 13662 30090 0 _0852_
rlabel metal1 14260 10710 14260 10710 0 _0853_
rlabel metal1 19504 9622 19504 9622 0 _0854_
rlabel metal1 29486 7378 29486 7378 0 _0855_
rlabel metal1 30222 5542 30222 5542 0 _0856_
rlabel metal1 14858 33626 14858 33626 0 _0857_
rlabel metal1 14766 34170 14766 34170 0 _0858_
rlabel metal1 16652 34034 16652 34034 0 _0859_
rlabel metal1 18630 33898 18630 33898 0 _0860_
rlabel metal1 18400 33966 18400 33966 0 _0861_
rlabel metal1 18354 33524 18354 33524 0 _0862_
rlabel metal1 18630 33490 18630 33490 0 _0863_
rlabel metal2 12558 34170 12558 34170 0 _0864_
rlabel metal2 18814 33643 18814 33643 0 _0865_
rlabel metal1 19262 33490 19262 33490 0 _0866_
rlabel metal3 20171 33252 20171 33252 0 _0867_
rlabel metal1 19412 4590 19412 4590 0 _0868_
rlabel metal1 17756 6834 17756 6834 0 _0869_
rlabel metal1 19642 35088 19642 35088 0 _0870_
rlabel metal1 19550 34952 19550 34952 0 _0871_
rlabel metal1 17066 34476 17066 34476 0 _0872_
rlabel metal1 17204 34170 17204 34170 0 _0873_
rlabel metal1 16514 34170 16514 34170 0 _0874_
rlabel via2 19458 34731 19458 34731 0 _0875_
rlabel metal1 18400 32402 18400 32402 0 _0876_
rlabel metal1 17112 33490 17112 33490 0 _0877_
rlabel metal2 18354 33184 18354 33184 0 _0878_
rlabel metal2 18722 32606 18722 32606 0 _0879_
rlabel metal3 18469 32028 18469 32028 0 _0880_
rlabel metal1 19458 5236 19458 5236 0 _0881_
rlabel metal1 20424 5202 20424 5202 0 _0882_
rlabel metal1 21620 6766 21620 6766 0 _0883_
rlabel metal1 19458 6834 19458 6834 0 _0884_
rlabel metal1 20286 10608 20286 10608 0 _0885_
rlabel viali 22402 25873 22402 25873 0 _0886_
rlabel metal1 21850 24378 21850 24378 0 _0887_
rlabel metal1 22632 24922 22632 24922 0 _0888_
rlabel metal1 21068 26350 21068 26350 0 _0889_
rlabel metal2 22586 26044 22586 26044 0 _0890_
rlabel metal1 22908 25466 22908 25466 0 _0891_
rlabel metal1 21022 25296 21022 25296 0 _0892_
rlabel metal2 20378 25704 20378 25704 0 _0893_
rlabel metal1 20930 24922 20930 24922 0 _0894_
rlabel metal1 21298 25228 21298 25228 0 _0895_
rlabel metal1 21068 9010 21068 9010 0 _0896_
rlabel metal1 20240 24174 20240 24174 0 _0897_
rlabel metal2 20470 22899 20470 22899 0 _0898_
rlabel metal1 21482 22202 21482 22202 0 _0899_
rlabel metal2 21022 22576 21022 22576 0 _0900_
rlabel metal1 20884 22202 20884 22202 0 _0901_
rlabel metal1 20516 22202 20516 22202 0 _0902_
rlabel metal2 19320 17510 19320 17510 0 _0903_
rlabel metal1 16376 24378 16376 24378 0 _0904_
rlabel metal1 16284 23494 16284 23494 0 _0905_
rlabel metal1 18676 13770 18676 13770 0 _0906_
rlabel metal1 20240 11118 20240 11118 0 _0907_
rlabel metal1 20102 10710 20102 10710 0 _0908_
rlabel metal1 19504 7378 19504 7378 0 _0909_
rlabel metal1 20562 7310 20562 7310 0 _0910_
rlabel metal1 20056 4794 20056 4794 0 _0911_
rlabel metal1 21160 5270 21160 5270 0 _0912_
rlabel metal1 30590 5168 30590 5168 0 _0913_
rlabel metal2 23230 27914 23230 27914 0 _0914_
rlabel metal1 22540 28050 22540 28050 0 _0915_
rlabel metal2 23322 27676 23322 27676 0 _0916_
rlabel metal1 23598 27506 23598 27506 0 _0917_
rlabel metal2 21482 27676 21482 27676 0 _0918_
rlabel metal1 21022 28050 21022 28050 0 _0919_
rlabel metal1 21206 27642 21206 27642 0 _0920_
rlabel metal2 20378 14331 20378 14331 0 _0921_
rlabel metal2 29026 9775 29026 9775 0 _0922_
rlabel metal1 24150 26010 24150 26010 0 _0923_
rlabel metal2 24242 28832 24242 28832 0 _0924_
rlabel metal1 23092 29002 23092 29002 0 _0925_
rlabel metal1 22356 29274 22356 29274 0 _0926_
rlabel metal1 23046 29138 23046 29138 0 _0927_
rlabel metal1 23966 25908 23966 25908 0 _0928_
rlabel metal1 22954 15504 22954 15504 0 _0929_
rlabel metal1 19596 28050 19596 28050 0 _0930_
rlabel metal1 19918 27642 19918 27642 0 _0931_
rlabel metal1 19964 27914 19964 27914 0 _0932_
rlabel metal2 21942 16031 21942 16031 0 _0933_
rlabel metal1 23276 15334 23276 15334 0 _0934_
rlabel metal2 32338 10880 32338 10880 0 _0935_
rlabel metal1 32154 8976 32154 8976 0 _0936_
rlabel metal2 28566 8636 28566 8636 0 _0937_
rlabel metal1 30636 10642 30636 10642 0 _0938_
rlabel metal1 23322 35088 23322 35088 0 _0939_
rlabel metal1 22494 37230 22494 37230 0 _0940_
rlabel metal2 23414 34986 23414 34986 0 _0941_
rlabel metal1 23506 35156 23506 35156 0 _0942_
rlabel metal1 23276 34510 23276 34510 0 _0943_
rlabel metal1 22954 34578 22954 34578 0 _0944_
rlabel metal1 23138 34612 23138 34612 0 _0945_
rlabel metal2 13110 15861 13110 15861 0 _0946_
rlabel metal1 24794 15470 24794 15470 0 _0947_
rlabel metal1 23736 29750 23736 29750 0 _0948_
rlabel metal1 23506 36890 23506 36890 0 _0949_
rlabel metal1 23368 37434 23368 37434 0 _0950_
rlabel metal2 22126 37434 22126 37434 0 _0951_
rlabel metal1 23506 37230 23506 37230 0 _0952_
rlabel metal1 23552 36346 23552 36346 0 _0953_
rlabel metal1 23874 37094 23874 37094 0 _0954_
rlabel metal3 23299 16524 23299 16524 0 _0955_
rlabel metal1 20930 34714 20930 34714 0 _0956_
rlabel metal2 22310 34748 22310 34748 0 _0957_
rlabel metal3 21919 33252 21919 33252 0 _0958_
rlabel metal1 25254 15470 25254 15470 0 _0959_
rlabel metal1 28888 12818 28888 12818 0 _0960_
rlabel metal2 15318 36346 15318 36346 0 _0961_
rlabel metal1 15272 37842 15272 37842 0 _0962_
rlabel metal2 15226 36890 15226 36890 0 _0963_
rlabel metal1 19458 36108 19458 36108 0 _0964_
rlabel metal1 15226 35802 15226 35802 0 _0965_
rlabel metal1 14076 36006 14076 36006 0 _0966_
rlabel metal1 13616 35802 13616 35802 0 _0967_
rlabel metal1 13202 36278 13202 36278 0 _0968_
rlabel metal1 13110 16558 13110 16558 0 _0969_
rlabel metal1 29854 16116 29854 16116 0 _0970_
rlabel metal1 20240 29818 20240 29818 0 _0971_
rlabel metal1 19780 37230 19780 37230 0 _0972_
rlabel metal1 18676 37434 18676 37434 0 _0973_
rlabel metal1 18814 37910 18814 37910 0 _0974_
rlabel metal1 19458 37298 19458 37298 0 _0975_
rlabel metal1 20194 36346 20194 36346 0 _0976_
rlabel metal2 20286 30668 20286 30668 0 _0977_
rlabel metal1 19872 16558 19872 16558 0 _0978_
rlabel metal1 18446 36108 18446 36108 0 _0979_
rlabel metal2 19366 17765 19366 17765 0 _0980_
rlabel metal1 19596 16558 19596 16558 0 _0981_
rlabel metal1 29164 14994 29164 14994 0 _0982_
rlabel metal1 30682 12818 30682 12818 0 _0983_
rlabel metal1 30866 11662 30866 11662 0 _0984_
rlabel metal2 31142 11492 31142 11492 0 _0985_
rlabel metal1 30590 16048 30590 16048 0 _0986_
rlabel metal1 26726 15130 26726 15130 0 _0987_
rlabel metal1 27186 15334 27186 15334 0 _0988_
rlabel metal1 30912 11730 30912 11730 0 _0989_
rlabel metal1 32614 18700 32614 18700 0 _0990_
rlabel metal1 32890 19380 32890 19380 0 _0991_
rlabel metal1 32338 19380 32338 19380 0 _0992_
rlabel metal1 32614 19278 32614 19278 0 _0993_
rlabel metal1 34914 19754 34914 19754 0 _0994_
rlabel metal1 35466 23120 35466 23120 0 _0995_
rlabel metal2 35282 20910 35282 20910 0 _0996_
rlabel metal1 34776 21114 34776 21114 0 _0997_
rlabel metal1 35374 23766 35374 23766 0 _0998_
rlabel metal1 34638 22678 34638 22678 0 _0999_
rlabel metal1 33534 21998 33534 21998 0 _1000_
rlabel metal1 30452 32402 30452 32402 0 _1001_
rlabel metal1 30958 32198 30958 32198 0 _1002_
rlabel metal1 31510 31110 31510 31110 0 _1003_
rlabel metal1 26036 31994 26036 31994 0 _1004_
rlabel metal1 25806 32436 25806 32436 0 _1005_
rlabel metal1 25806 32198 25806 32198 0 _1006_
rlabel metal1 27554 23596 27554 23596 0 _1007_
rlabel metal1 32476 24038 32476 24038 0 _1008_
rlabel metal1 33074 24378 33074 24378 0 _1009_
rlabel metal1 32568 24650 32568 24650 0 _1010_
rlabel metal2 32062 24412 32062 24412 0 _1011_
rlabel metal1 30452 28050 30452 28050 0 _1012_
rlabel metal1 30498 27574 30498 27574 0 _1013_
rlabel metal1 30912 24174 30912 24174 0 _1014_
rlabel metal1 26542 28492 26542 28492 0 _1015_
rlabel metal1 26266 28118 26266 28118 0 _1016_
rlabel metal2 26910 36108 26910 36108 0 _1017_
rlabel metal1 30774 24140 30774 24140 0 _1018_
rlabel metal1 31280 23698 31280 23698 0 _1019_
rlabel metal1 31970 23834 31970 23834 0 _1020_
rlabel metal1 31234 22678 31234 22678 0 _1021_
rlabel metal1 32430 22644 32430 22644 0 _1022_
rlabel metal2 32430 24004 32430 24004 0 _1023_
rlabel metal2 31878 23018 31878 23018 0 _1024_
rlabel metal2 30406 22100 30406 22100 0 _1025_
rlabel metal1 29992 20434 29992 20434 0 _1026_
rlabel metal2 29486 35972 29486 35972 0 _1027_
rlabel metal2 29302 33601 29302 33601 0 _1028_
rlabel metal1 28060 19822 28060 19822 0 _1029_
rlabel metal1 25714 35700 25714 35700 0 _1030_
rlabel metal1 25898 35088 25898 35088 0 _1031_
rlabel metal1 25576 19822 25576 19822 0 _1032_
rlabel metal1 26082 19720 26082 19720 0 _1033_
rlabel metal1 28704 20026 28704 20026 0 _1034_
rlabel metal1 29210 19346 29210 19346 0 _1035_
rlabel metal1 28658 18700 28658 18700 0 _1036_
rlabel metal1 28842 19822 28842 19822 0 _1037_
rlabel metal2 29486 19788 29486 19788 0 _1038_
rlabel metal1 20884 16966 20884 16966 0 _1039_
rlabel metal2 20286 17442 20286 17442 0 _1040_
rlabel metal1 20544 17170 20544 17170 0 _1041_
rlabel metal1 21298 17204 21298 17204 0 _1042_
rlabel metal1 28842 10642 28842 10642 0 _1043_
rlabel metal1 20746 14416 20746 14416 0 _1044_
rlabel metal1 21022 15028 21022 15028 0 _1045_
rlabel metal1 20562 13974 20562 13974 0 _1046_
rlabel metal1 22034 14348 22034 14348 0 _1047_
rlabel metal1 22586 12818 22586 12818 0 _1048_
rlabel metal2 33212 8942 33212 8942 0 _1049_
rlabel metal1 30774 14382 30774 14382 0 _1050_
rlabel metal1 30176 19346 30176 19346 0 _1051_
rlabel metal1 34592 21658 34592 21658 0 _1052_
rlabel metal1 35006 19380 35006 19380 0 _1053_
rlabel metal1 34960 19142 34960 19142 0 _1054_
rlabel metal1 32752 18190 32752 18190 0 _1055_
rlabel metal2 28382 8092 28382 8092 0 _1056_
rlabel metal1 25622 6800 25622 6800 0 _1057_
rlabel metal1 21850 6800 21850 6800 0 _1058_
rlabel metal1 21344 7310 21344 7310 0 _1059_
rlabel metal1 26772 3910 26772 3910 0 _1060_
rlabel metal1 27462 7446 27462 7446 0 _1061_
rlabel metal1 25990 7310 25990 7310 0 _1062_
rlabel metal1 28520 7854 28520 7854 0 _1063_
rlabel metal1 29854 8942 29854 8942 0 _1064_
rlabel metal1 29900 9690 29900 9690 0 _1065_
rlabel metal1 25990 14960 25990 14960 0 _1066_
rlabel metal1 26542 12886 26542 12886 0 _1067_
rlabel metal1 26588 15062 26588 15062 0 _1068_
rlabel metal1 31786 14484 31786 14484 0 _1069_
rlabel metal1 27232 13294 27232 13294 0 _1070_
rlabel metal1 27554 11050 27554 11050 0 _1071_
rlabel metal1 27094 15402 27094 15402 0 _1072_
rlabel metal1 27186 11594 27186 11594 0 _1073_
rlabel metal1 27324 13158 27324 13158 0 _1074_
rlabel metal2 25806 14042 25806 14042 0 _1075_
rlabel metal1 26220 13294 26220 13294 0 _1076_
rlabel metal2 26358 12988 26358 12988 0 _1077_
rlabel metal1 28106 12240 28106 12240 0 _1078_
rlabel metal1 30268 17646 30268 17646 0 _1079_
rlabel metal2 35190 18598 35190 18598 0 _1080_
rlabel metal1 34454 19346 34454 19346 0 _1081_
rlabel metal1 34868 20366 34868 20366 0 _1082_
rlabel metal1 34684 23698 34684 23698 0 _1083_
rlabel metal1 34546 22066 34546 22066 0 _1084_
rlabel metal2 32338 22066 32338 22066 0 _1085_
rlabel metal1 32798 24140 32798 24140 0 _1086_
rlabel metal2 32614 21801 32614 21801 0 _1087_
rlabel metal2 30498 21624 30498 21624 0 _1088_
rlabel metal1 28842 20468 28842 20468 0 _1089_
rlabel metal1 30406 19380 30406 19380 0 _1090_
rlabel metal1 22862 14586 22862 14586 0 _1091_
rlabel metal1 33626 21522 33626 21522 0 _1092_
rlabel metal1 31372 14382 31372 14382 0 _1093_
rlabel metal1 30866 19278 30866 19278 0 _1094_
rlabel metal1 29900 15470 29900 15470 0 _1095_
rlabel metal1 30774 16014 30774 16014 0 _1096_
rlabel metal1 31418 15504 31418 15504 0 _1097_
rlabel metal1 33120 14450 33120 14450 0 _1098_
rlabel metal1 29670 15538 29670 15538 0 _1099_
rlabel metal1 31050 13328 31050 13328 0 _1100_
rlabel metal1 33810 14042 33810 14042 0 _1101_
rlabel metal1 33810 12852 33810 12852 0 _1102_
rlabel metal2 33534 13124 33534 13124 0 _1103_
rlabel metal1 30130 6324 30130 6324 0 _1104_
rlabel metal1 32706 6834 32706 6834 0 _1105_
rlabel metal1 26818 4046 26818 4046 0 _1106_
rlabel metal1 20102 4556 20102 4556 0 _1107_
rlabel metal1 20010 5644 20010 5644 0 _1108_
rlabel metal1 20240 9894 20240 9894 0 _1109_
rlabel metal1 19826 5746 19826 5746 0 _1110_
rlabel metal1 19182 4760 19182 4760 0 _1111_
rlabel metal1 26634 4148 26634 4148 0 _1112_
rlabel metal1 28704 4590 28704 4590 0 _1113_
rlabel metal1 32338 5678 32338 5678 0 _1114_
rlabel metal2 31970 5508 31970 5508 0 _1115_
rlabel metal1 32614 6256 32614 6256 0 _1116_
rlabel metal1 33212 6766 33212 6766 0 _1117_
rlabel metal1 33258 8908 33258 8908 0 _1118_
rlabel metal1 33626 13226 33626 13226 0 _1119_
rlabel metal1 33396 14382 33396 14382 0 _1120_
rlabel metal1 33304 14518 33304 14518 0 _1121_
rlabel metal1 21390 13294 21390 13294 0 _1122_
rlabel metal1 29118 10676 29118 10676 0 _1123_
rlabel metal1 33350 13838 33350 13838 0 _1124_
rlabel metal1 33220 15062 33220 15062 0 _1125_
rlabel metal1 27830 15062 27830 15062 0 _1126_
rlabel metal1 29670 10103 29670 10103 0 _1127_
rlabel metal1 30544 12750 30544 12750 0 _1128_
rlabel metal2 29026 12869 29026 12869 0 _1129_
rlabel metal1 28750 13328 28750 13328 0 _1130_
rlabel metal2 31510 13600 31510 13600 0 _1131_
rlabel metal1 32614 10642 32614 10642 0 _1132_
rlabel metal1 30084 9894 30084 9894 0 _1133_
rlabel metal1 32200 9894 32200 9894 0 _1134_
rlabel metal1 29946 8534 29946 8534 0 _1135_
rlabel metal2 30590 8126 30590 8126 0 _1136_
rlabel metal1 23000 5678 23000 5678 0 _1137_
rlabel metal1 19826 6698 19826 6698 0 _1138_
rlabel metal1 20838 7446 20838 7446 0 _1139_
rlabel metal1 21260 9622 21260 9622 0 _1140_
rlabel metal1 21528 9350 21528 9350 0 _1141_
rlabel metal1 22586 5644 22586 5644 0 _1142_
rlabel metal2 22954 5474 22954 5474 0 _1143_
rlabel metal1 26588 4250 26588 4250 0 _1144_
rlabel metal2 28106 5202 28106 5202 0 _1145_
rlabel metal2 31786 8160 31786 8160 0 _1146_
rlabel metal1 31050 8602 31050 8602 0 _1147_
rlabel metal2 29302 12971 29302 12971 0 _1148_
rlabel metal1 28658 13260 28658 13260 0 _1149_
rlabel metal1 21344 16558 21344 16558 0 _1150_
rlabel metal2 32936 12818 32936 12818 0 _1151_
rlabel metal1 28106 13498 28106 13498 0 _1152_
rlabel metal1 28704 14382 28704 14382 0 _1153_
rlabel metal1 33074 11084 33074 11084 0 _1154_
rlabel metal2 31786 14416 31786 14416 0 _1155_
rlabel metal1 30958 14280 30958 14280 0 _1156_
rlabel metal2 28198 15062 28198 15062 0 _1157_
rlabel metal1 28474 15029 28474 15029 0 _1158_
rlabel via1 21858 12070 21858 12070 0 _1159_
rlabel metal1 22632 13906 22632 13906 0 _1160_
rlabel via1 27904 6766 27904 6766 0 _1161_
rlabel metal1 22770 8466 22770 8466 0 _1162_
rlabel metal1 21275 12954 21275 12954 0 _1163_
rlabel metal2 23414 13056 23414 13056 0 _1164_
rlabel metal1 25162 12886 25162 12886 0 _1165_
rlabel metal1 33028 13226 33028 13226 0 _1166_
rlabel metal1 25162 13328 25162 13328 0 _1167_
rlabel metal2 22034 7446 22034 7446 0 _1168_
rlabel metal1 25254 13328 25254 13328 0 _1169_
rlabel metal1 25116 13498 25116 13498 0 _1170_
rlabel metal1 21344 11730 21344 11730 0 _1171_
rlabel metal2 20746 8364 20746 8364 0 _1172_
rlabel metal1 21988 12614 21988 12614 0 _1173_
rlabel metal1 25392 11730 25392 11730 0 _1174_
rlabel metal1 22954 8942 22954 8942 0 _1175_
rlabel metal1 25208 11866 25208 11866 0 _1176_
rlabel metal1 24886 12308 24886 12308 0 _1177_
rlabel metal2 24426 12614 24426 12614 0 _1178_
rlabel metal2 25070 14212 25070 14212 0 _1179_
rlabel metal1 27692 14586 27692 14586 0 _1180_
rlabel metal2 28290 14518 28290 14518 0 _1181_
rlabel metal2 17894 21182 17894 21182 0 _1182_
rlabel metal1 25944 19482 25944 19482 0 _1183_
rlabel metal2 33166 36448 33166 36448 0 _1184_
rlabel via1 15136 20434 15136 20434 0 _1185_
rlabel metal1 14789 20910 14789 20910 0 _1186_
rlabel metal1 14398 20842 14398 20842 0 _1187_
rlabel metal1 14536 22610 14536 22610 0 _1188_
rlabel metal1 15640 18394 15640 18394 0 _1189_
rlabel metal1 14398 20026 14398 20026 0 _1190_
rlabel metal2 14306 21488 14306 21488 0 _1191_
rlabel metal2 14674 24820 14674 24820 0 _1192_
rlabel metal1 15226 20570 15226 20570 0 _1193_
rlabel metal1 14996 13498 14996 13498 0 _1194_
rlabel metal1 15134 13940 15134 13940 0 _1195_
rlabel via1 14953 14042 14953 14042 0 _1196_
rlabel metal2 15502 16082 15502 16082 0 _1197_
rlabel metal1 15410 14042 15410 14042 0 _1198_
rlabel metal1 14306 14416 14306 14416 0 _1199_
rlabel metal1 14490 13974 14490 13974 0 _1200_
rlabel metal1 13294 17306 13294 17306 0 _1201_
rlabel metal1 15134 25371 15134 25371 0 _1202_
rlabel metal1 33120 32198 33120 32198 0 _1203_
rlabel metal1 34454 31858 34454 31858 0 _1204_
rlabel metal2 32982 13498 32982 13498 0 _1205_
rlabel metal1 31878 13396 31878 13396 0 _1206_
rlabel metal1 30820 12682 30820 12682 0 _1207_
rlabel metal1 32170 12954 32170 12954 0 _1208_
rlabel metal2 31970 13090 31970 13090 0 _1209_
rlabel metal1 30866 13226 30866 13226 0 _1210_
rlabel metal1 31004 14042 31004 14042 0 _1211_
rlabel metal1 30498 14450 30498 14450 0 _1212_
rlabel metal1 30590 13226 30590 13226 0 _1213_
rlabel metal1 25944 9078 25944 9078 0 _1214_
rlabel metal1 26036 13294 26036 13294 0 _1215_
rlabel metal1 27462 12852 27462 12852 0 _1216_
rlabel metal1 26956 12410 26956 12410 0 _1217_
rlabel metal1 28198 12614 28198 12614 0 _1218_
rlabel metal1 31418 13294 31418 13294 0 _1219_
rlabel metal2 32154 15028 32154 15028 0 _1220_
rlabel metal1 7130 18632 7130 18632 0 _1221_
rlabel metal1 29992 21862 29992 21862 0 _1222_
rlabel metal1 30038 20842 30038 20842 0 _1223_
rlabel metal2 17618 21148 17618 21148 0 _1224_
rlabel metal1 27232 21114 27232 21114 0 _1225_
rlabel metal1 26358 29614 26358 29614 0 _1226_
rlabel metal1 31924 8058 31924 8058 0 _1227_
rlabel metal2 30866 9350 30866 9350 0 _1228_
rlabel metal1 31786 10506 31786 10506 0 _1229_
rlabel metal1 26450 10642 26450 10642 0 _1230_
rlabel metal1 27186 10064 27186 10064 0 _1231_
rlabel metal1 27370 9996 27370 9996 0 _1232_
rlabel metal1 30222 9996 30222 9996 0 _1233_
rlabel metal1 31096 9554 31096 9554 0 _1234_
rlabel metal1 33534 9622 33534 9622 0 _1235_
rlabel metal1 33074 6695 33074 6695 0 _1236_
rlabel metal2 32522 7888 32522 7888 0 _1237_
rlabel metal2 32614 9350 32614 9350 0 _1238_
rlabel metal2 13110 19006 13110 19006 0 _1239_
rlabel metal1 32614 22644 32614 22644 0 _1240_
rlabel metal1 31694 21556 31694 21556 0 _1241_
rlabel metal1 31694 22542 31694 22542 0 _1242_
rlabel metal1 31556 21522 31556 21522 0 _1243_
rlabel metal1 32062 22100 32062 22100 0 _1244_
rlabel metal1 31326 21658 31326 21658 0 _1245_
rlabel metal1 15778 21998 15778 21998 0 _1246_
rlabel metal1 28474 32878 28474 32878 0 _1247_
rlabel metal1 31786 32334 31786 32334 0 _1248_
rlabel metal1 31970 7412 31970 7412 0 _1249_
rlabel metal1 30406 4624 30406 4624 0 _1250_
rlabel metal1 30590 4794 30590 4794 0 _1251_
rlabel metal1 30682 6732 30682 6732 0 _1252_
rlabel metal1 23736 9146 23736 9146 0 _1253_
rlabel metal1 23575 9962 23575 9962 0 _1254_
rlabel metal1 22632 10642 22632 10642 0 _1255_
rlabel metal1 24656 8602 24656 8602 0 _1256_
rlabel metal1 27692 8534 27692 8534 0 _1257_
rlabel metal1 27140 8602 27140 8602 0 _1258_
rlabel metal1 28658 8908 28658 8908 0 _1259_
rlabel metal1 27186 9588 27186 9588 0 _1260_
rlabel metal2 28842 9146 28842 9146 0 _1261_
rlabel metal1 29716 6766 29716 6766 0 _1262_
rlabel metal1 31142 6902 31142 6902 0 _1263_
rlabel metal2 32154 6868 32154 6868 0 _1264_
rlabel metal2 9890 16575 9890 16575 0 _1265_
rlabel metal1 32798 21930 32798 21930 0 _1266_
rlabel metal2 32890 21828 32890 21828 0 _1267_
rlabel metal1 32476 20978 32476 20978 0 _1268_
rlabel metal2 29118 25364 29118 25364 0 _1269_
rlabel metal1 33902 25262 33902 25262 0 _1270_
rlabel metal1 27094 4182 27094 4182 0 _1271_
rlabel metal1 28106 4148 28106 4148 0 _1272_
rlabel metal1 28244 3910 28244 3910 0 _1273_
rlabel metal1 27968 5882 27968 5882 0 _1274_
rlabel metal2 13938 19856 13938 19856 0 clk
rlabel metal2 32246 30090 32246 30090 0 clknet_0__0514_
rlabel metal1 13386 25942 13386 25942 0 clknet_0__0515_
rlabel metal1 20332 31926 20332 31926 0 clknet_0__0516_
rlabel metal1 14122 32402 14122 32402 0 clknet_0__0517_
rlabel metal2 9798 8160 9798 8160 0 clknet_0_clk
rlabel metal1 29394 31280 29394 31280 0 clknet_1_0__leaf__0514_
rlabel metal1 14306 31790 14306 31790 0 clknet_1_0__leaf__0515_
rlabel metal1 20286 38284 20286 38284 0 clknet_1_0__leaf__0516_
rlabel metal1 9522 31892 9522 31892 0 clknet_1_0__leaf__0517_
rlabel metal1 34132 27438 34132 27438 0 clknet_1_1__leaf__0514_
rlabel metal1 15548 25670 15548 25670 0 clknet_1_1__leaf__0515_
rlabel metal1 33626 28526 33626 28526 0 clknet_1_1__leaf__0516_
rlabel metal1 31878 38352 31878 38352 0 clknet_1_1__leaf__0517_
rlabel metal1 1426 17238 1426 17238 0 clknet_2_0__leaf_clk
rlabel metal1 1426 23732 1426 23732 0 clknet_2_1__leaf_clk
rlabel metal2 1426 12784 1426 12784 0 clknet_2_2__leaf_clk
rlabel metal1 14720 10642 14720 10642 0 clknet_2_3__leaf_clk
rlabel metal1 37812 8942 37812 8942 0 cs
rlabel metal3 820 11628 820 11628 0 gpi[0]
rlabel metal3 1096 6868 1096 6868 0 gpi[1]
rlabel metal1 31050 38998 31050 38998 0 gpi[23]
rlabel metal2 10994 1095 10994 1095 0 gpi[2]
rlabel metal2 8418 1027 8418 1027 0 gpi[3]
rlabel metal1 15594 38998 15594 38998 0 gpi[4]
rlabel metal1 37444 38930 37444 38930 0 gpi[5]
rlabel metal2 37398 1027 37398 1027 0 gpi[6]
rlabel metal1 20056 38930 20056 38930 0 gpi[7]
rlabel metal1 17664 39066 17664 39066 0 gpo[0]
rlabel metal3 820 4148 820 4148 0 gpo[10]
rlabel metal2 37950 10999 37950 10999 0 gpo[11]
rlabel metal3 820 8908 820 8908 0 gpo[12]
rlabel metal2 37858 15793 37858 15793 0 gpo[13]
rlabel metal1 828 39066 828 39066 0 gpo[14]
rlabel metal1 26818 39066 26818 39066 0 gpo[15]
rlabel metal2 17434 1520 17434 1520 0 gpo[16]
rlabel metal2 46 1520 46 1520 0 gpo[17]
rlabel metal3 751 25228 751 25228 0 gpo[18]
rlabel metal2 21942 39960 21942 39960 0 gpo[19]
rlabel metal3 820 15708 820 15708 0 gpo[1]
rlabel metal1 37904 38522 37904 38522 0 gpo[20]
rlabel metal1 13064 39066 13064 39066 0 gpo[21]
rlabel metal2 3910 1571 3910 1571 0 gpo[22]
rlabel metal2 1978 1520 1978 1520 0 gpo[23]
rlabel metal2 37858 36941 37858 36941 0 gpo[24]
rlabel metal3 820 18428 820 18428 0 gpo[25]
rlabel metal2 14858 1520 14858 1520 0 gpo[26]
rlabel metal1 37904 34510 37904 34510 0 gpo[27]
rlabel metal3 37958 1428 37958 1428 0 gpo[28]
rlabel metal1 9292 39066 9292 39066 0 gpo[29]
rlabel metal1 38134 20774 38134 20774 0 gpo[2]
rlabel metal2 6486 823 6486 823 0 gpo[30]
rlabel metal2 12926 1520 12926 1520 0 gpo[31]
rlabel metal3 820 20468 820 20468 0 gpo[32]
rlabel via2 37858 22491 37858 22491 0 gpo[33]
rlabel metal2 19366 1520 19366 1520 0 gpo[3]
rlabel metal1 35972 38998 35972 38998 0 gpo[4]
rlabel metal1 33028 39066 33028 39066 0 gpo[5]
rlabel metal1 4784 39066 4784 39066 0 gpo[6]
rlabel metal1 11408 39066 11408 39066 0 gpo[7]
rlabel metal2 26450 1520 26450 1520 0 gpo[8]
rlabel metal3 820 13668 820 13668 0 gpo[9]
rlabel metal1 16560 9554 16560 9554 0 net1
rlabel metal1 11730 20910 11730 20910 0 net10
rlabel metal1 20470 38318 20470 38318 0 net100
rlabel metal1 24288 26350 24288 26350 0 net101
rlabel metal1 30130 35700 30130 35700 0 net102
rlabel metal1 26956 28594 26956 28594 0 net103
rlabel metal1 34776 30770 34776 30770 0 net104
rlabel metal1 34086 28084 34086 28084 0 net105
rlabel metal2 32890 33830 32890 33830 0 net106
rlabel metal1 24840 38386 24840 38386 0 net107
rlabel metal2 31970 38080 31970 38080 0 net108
rlabel metal2 7866 24922 7866 24922 0 net109
rlabel metal1 2714 20332 2714 20332 0 net11
rlabel metal1 6992 36210 6992 36210 0 net110
rlabel metal1 11546 28084 11546 28084 0 net111
rlabel metal2 9430 31450 9430 31450 0 net112
rlabel metal1 6762 28084 6762 28084 0 net113
rlabel metal1 7038 33524 7038 33524 0 net114
rlabel metal1 10074 38318 10074 38318 0 net115
rlabel metal1 8418 37876 8418 37876 0 net116
rlabel metal1 28060 23698 28060 23698 0 net117
rlabel metal1 27002 34612 27002 34612 0 net118
rlabel metal1 27186 26010 27186 26010 0 net119
rlabel metal1 17710 38964 17710 38964 0 net12
rlabel metal2 29118 30362 29118 30362 0 net120
rlabel viali 29578 28524 29578 28524 0 net121
rlabel metal1 28198 33524 28198 33524 0 net122
rlabel metal1 26910 38318 26910 38318 0 net123
rlabel metal1 29440 38318 29440 38318 0 net124
rlabel metal2 29118 26010 29118 26010 0 net125
rlabel metal1 8832 4250 8832 4250 0 net126
rlabel metal1 8234 5746 8234 5746 0 net127
rlabel metal2 11454 6970 11454 6970 0 net128
rlabel metal1 8832 6426 8832 6426 0 net129
rlabel metal1 2070 4590 2070 4590 0 net13
rlabel metal1 9936 5270 9936 5270 0 net130
rlabel metal1 13156 4250 13156 4250 0 net131
rlabel metal2 10074 32674 10074 32674 0 net132
rlabel metal1 14674 5780 14674 5780 0 net133
rlabel metal1 15732 5134 15732 5134 0 net134
rlabel metal1 8326 30294 8326 30294 0 net135
rlabel metal1 8234 28458 8234 28458 0 net136
rlabel metal2 10442 28730 10442 28730 0 net137
rlabel metal1 7498 30736 7498 30736 0 net138
rlabel metal1 10925 5338 10925 5338 0 net139
rlabel via2 19274 11611 19274 11611 0 net14
rlabel metal2 1518 9418 1518 9418 0 net15
rlabel metal2 37674 16031 37674 16031 0 net16
rlabel metal1 2668 38930 2668 38930 0 net17
rlabel metal3 25553 38692 25553 38692 0 net18
rlabel metal1 17526 2414 17526 2414 0 net19
rlabel metal1 1702 11288 1702 11288 0 net2
rlabel metal2 1564 4556 1564 4556 0 net20
rlabel metal1 1840 22746 1840 22746 0 net21
rlabel metal1 22862 21318 22862 21318 0 net22
rlabel metal1 1794 20230 1794 20230 0 net23
rlabel metal1 34684 38250 34684 38250 0 net24
rlabel metal2 13018 38811 13018 38811 0 net25
rlabel metal2 4094 2587 4094 2587 0 net26
rlabel metal2 2162 4657 2162 4657 0 net27
rlabel via2 13386 21675 13386 21675 0 net28
rlabel metal1 1656 18734 1656 18734 0 net29
rlabel metal2 8970 20434 8970 20434 0 net3
rlabel metal1 15640 2414 15640 2414 0 net30
rlabel metal1 37490 33626 37490 33626 0 net31
rlabel metal1 37582 2992 37582 2992 0 net32
rlabel metal2 9338 38726 9338 38726 0 net33
rlabel metal1 37398 20842 37398 20842 0 net34
rlabel metal1 7452 2414 7452 2414 0 net35
rlabel metal1 13064 2414 13064 2414 0 net36
rlabel metal2 1840 23188 1840 23188 0 net37
rlabel metal1 37536 22610 37536 22610 0 net38
rlabel metal1 20746 2414 20746 2414 0 net39
rlabel metal2 11914 20927 11914 20927 0 net4
rlabel metal1 35190 38522 35190 38522 0 net40
rlabel metal1 32614 38522 32614 38522 0 net41
rlabel metal1 4922 38522 4922 38522 0 net42
rlabel metal1 11592 37978 11592 37978 0 net43
rlabel metal1 10442 2414 10442 2414 0 net44
rlabel metal1 1518 13192 1518 13192 0 net45
rlabel metal1 2254 21556 2254 21556 0 net46
rlabel metal1 4554 8976 4554 8976 0 net47
rlabel metal1 35420 18802 35420 18802 0 net48
rlabel metal2 14766 35020 14766 35020 0 net49
rlabel metal1 9706 20502 9706 20502 0 net5
rlabel metal1 22310 27438 22310 27438 0 net50
rlabel metal1 20746 27336 20746 27336 0 net51
rlabel metal1 18906 24650 18906 24650 0 net52
rlabel metal2 21390 23902 21390 23902 0 net53
rlabel viali 22402 21976 22402 21976 0 net54
rlabel metal1 17059 8534 17059 8534 0 net55
rlabel metal1 14083 8874 14083 8874 0 net56
rlabel metal1 2507 12818 2507 12818 0 net57
rlabel metal1 9069 29206 9069 29206 0 net58
rlabel metal1 8609 36074 8609 36074 0 net59
rlabel metal1 9384 20910 9384 20910 0 net6
rlabel metal2 32706 35938 32706 35938 0 net60
rlabel metal1 35965 32402 35965 32402 0 net61
rlabel metal1 27002 32436 27002 32436 0 net62
rlabel metal1 34776 26418 34776 26418 0 net63
rlabel metal1 34362 29172 34362 29172 0 net64
rlabel metal2 34362 26010 34362 26010 0 net65
rlabel metal1 31832 31450 31832 31450 0 net66
rlabel metal2 27002 30362 27002 30362 0 net67
rlabel metal1 34638 32436 34638 32436 0 net68
rlabel metal1 9798 23086 9798 23086 0 net69
rlabel metal1 15778 38760 15778 38760 0 net7
rlabel metal1 9522 33524 9522 33524 0 net70
rlabel metal1 9614 25262 9614 25262 0 net71
rlabel metal2 6394 30362 6394 30362 0 net72
rlabel metal1 7498 29172 7498 29172 0 net73
rlabel metal1 5934 31450 5934 31450 0 net74
rlabel metal1 9522 29172 9522 29172 0 net75
rlabel metal1 7866 34612 7866 34612 0 net76
rlabel metal1 5198 25262 5198 25262 0 net77
rlabel metal1 4370 34612 4370 34612 0 net78
rlabel metal1 8142 26996 8142 26996 0 net79
rlabel metal1 9476 13838 9476 13838 0 net8
rlabel metal1 10258 31790 10258 31790 0 net80
rlabel metal1 4186 29172 4186 29172 0 net81
rlabel metal1 4370 33524 4370 33524 0 net82
rlabel metal1 9062 35802 9062 35802 0 net83
rlabel metal1 10166 35054 10166 35054 0 net84
rlabel metal1 24242 23698 24242 23698 0 net85
rlabel metal1 30958 33966 30958 33966 0 net86
rlabel metal1 31510 26010 31510 26010 0 net87
rlabel metal1 32154 30260 32154 30260 0 net88
rlabel metal2 31510 28730 31510 28730 0 net89
rlabel metal1 18239 2482 18239 2482 0 net9
rlabel metal1 32706 32470 32706 32470 0 net90
rlabel metal1 27508 36210 27508 36210 0 net91
rlabel metal1 32430 36142 32430 36142 0 net92
rlabel metal1 5014 26350 5014 26350 0 net93
rlabel metal1 4922 36142 4922 36142 0 net94
rlabel metal1 10166 26350 10166 26350 0 net95
rlabel metal1 7682 32198 7682 32198 0 net96
rlabel metal1 4186 28084 4186 28084 0 net97
rlabel metal1 4002 31450 4002 31450 0 net98
rlabel metal1 12236 38386 12236 38386 0 net99
rlabel metal3 820 36788 820 36788 0 nrst
rlabel metal1 38134 18054 38134 18054 0 store_en
<< properties >>
string FIXED_BBOX 0 0 39418 41562
<< end >>
