* NGSPICE file created from Synthia.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

.subckt Synthia PWM_o clk modes octaves pb[0] pb[10] pb[11] pb[12] pb[1] pb[2] pb[3]
+ pb[4] pb[5] pb[6] pb[7] pb[8] pb[9] reset vccd1 vssd1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3155_ _0301_ _0721_ _0307_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a21oi_4
X_2106_ d2.count\[3\] _1733_ _1772_ _1712_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__a2bb2o_1
X_3086_ _0646_ _0647_ _0651_ _0652_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2037_ _1712_ _1713_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__nand2_4
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3988_ _1546_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2939_ _1735_ d8.count\[5\] _1988_ _1986_ _0537_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_72_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire18 net19 vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3911_ _1385_ _1389_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3842_ d1.saw_temp\[6\] _0330_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3773_ _1710_ net61 _0782_ em0.u1.R\[13\] _1334_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ _0363_ _0367_ _0382_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__o21a_1
X_2655_ p0.count\[1\] vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2586_ d13.count\[0\] d13.count\[1\] vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__nand2_1
X_4325_ clknet_leaf_6_clk _0048_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_4
X_4256_ clknet_leaf_33_clk _0019_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_4
X_4187_ _1705_ _1706_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__and2_1
X_3207_ _0760_ _0768_ _0772_ _0773_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__a31o_1
X_3138_ d8.saw_temp\[7\] _0301_ _0337_ _0307_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__a31o_2
XFILLER_0_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3069_ d13.saw_temp\[4\] d13.saw_temp\[2\] d13.saw_temp\[1\] _0344_ vssd1 vssd1 vccd1
+ vccd1 _0636_ sky130_fd_sc_hd__o31a_1
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold170 d5.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 d3.count\[4\] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 d3.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2440_ _0152_ _0153_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2371_ _1720_ _1981_ d8.count\[3\] vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__a21oi_1
X_4110_ net128 _0782_ _1662_ _1710_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4041_ _1598_ _1599_ _1596_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3825_ d10.saw_temp\[7\] _0672_ _0674_ d10.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1
+ _1386_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3756_ _1206_ _1208_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__and2_1
X_2707_ _0366_ _0332_ _0331_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3687_ _1247_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__nor2_1
X_2638_ m0.edgo.delay m0.edgo.in vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2569_ _0253_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_4308_ clknet_leaf_19_clk _0041_ net39 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
X_4239_ clknet_leaf_32_clk _0012_ net27 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_92_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3610_ _0681_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3541_ _1102_ _1104_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3472_ _1034_ _1035_ _0646_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__mux2_1
X_2423_ d9.count\[0\] d9.count\[1\] vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__or2_1
X_2354_ net181 _1966_ _1959_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2285_ d6.count\[5\] _1910_ _1724_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__a21oi_1
X_4024_ _1536_ _1538_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3808_ _1368_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3739_ _1189_ _1191_ _1300_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2070_ d1.count\[0\] d1.count\[1\] vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2972_ _0560_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3524_ _0750_ _1087_ _0875_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__a21oi_2
X_3455_ _0920_ _0924_ _0931_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__o21a_1
X_2406_ d8.count\[8\] _2006_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__xnor2_1
X_3386_ d9.saw_temp\[2\] _0335_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nand2_1
X_2337_ _1721_ d7.count\[7\] d7.count\[8\] _1805_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2268_ net194 _1898_ _1888_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4007_ _1565_ _1522_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__or2_1
X_2199_ d4.count\[2\] _1724_ _1843_ d4.count\[7\] _1845_ vssd1 vssd1 vccd1 vccd1 _1846_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold30 p0.count\[7\] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 em0.u1.Q\[1\] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 d9.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold63 d3.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 em0.u1.Q\[3\] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 d11.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 em0.u1.D\[8\] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ d8.saw_temp\[7\] _0337_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__or2b_1
X_3171_ _0723_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__buf_6
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ d2.count\[1\] d2.count\[0\] d2.count\[2\] vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2053_ d1.count\[2\] _1729_ d1.count\[3\] vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2955_ _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__and2_1
X_2886_ _0497_ _0500_ d6.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3507_ d1.saw_temp\[2\] _0623_ _0627_ _1070_ _0618_ vssd1 vssd1 vccd1 vccd1 _1071_
+ sky130_fd_sc_hd__o311a_1
X_4487_ clknet_leaf_25_clk p0.pwm net34 vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3438_ _1000_ _1001_ _0760_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__mux2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _0916_ _0845_ _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__a21o_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _0395_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2671_ _0329_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__nand2_1
X_4410_ clknet_leaf_0_clk d12.nxt_count\[1\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4341_ clknet_leaf_29_clk d8.nxt_count\[8\] net24 vssd1 vssd1 vccd1 vccd1 d8.count\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4272_ clknet_leaf_24_clk _0025_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_4
X_3223_ d4.saw_temp\[7\] _0752_ _0759_ d4.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0789_
+ sky130_fd_sc_hd__o22a_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ d6.saw_temp\[7\] _0346_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__and2_2
X_2105_ _1727_ d2.count\[5\] d2.count\[4\] vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3085_ d12.saw_temp\[0\] _0340_ _0640_ _0309_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2036_ d1.oct_dwn\[0\] vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__buf_6
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _1434_ _1447_ _1545_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2938_ d8.count\[0\] vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2869_ _0487_ _0488_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__nor2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire19 _0580_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3910_ _0705_ _1362_ _1367_ _1374_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_80_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ d1.saw_temp\[5\] _0623_ _0627_ _1292_ d1.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1
+ _1402_ sky130_fd_sc_hd__o32a_1
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3772_ _1331_ _1333_ _0893_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2723_ _0380_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2654_ p0.count\[2\] vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
X_2585_ d13.count\[0\] d13.count\[1\] vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4324_ clknet_leaf_31_clk net48 net31 vssd1 vssd1 vccd1 vccd1 d7.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4255_ clknet_leaf_33_clk _0018_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
X_4186_ d9.saw_temp\[5\] _1703_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__or2_1
X_3206_ d3.saw_temp\[0\] _0348_ _0738_ _0310_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__a31o_1
X_3137_ d8.saw_temp\[0\] _0337_ _0682_ _0310_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3068_ d13.saw_temp\[7\] _0344_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__and2_2
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold160 d12.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _0485_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 d10.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 em0.u1.D\[10\] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2370_ _1727_ d8.count\[1\] d8.count\[2\] _1735_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4040_ em0.u1.R\[15\] em0.u1.D\[8\] vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3824_ _0750_ _1384_ _0659_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3755_ _1270_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__xnor2_1
X_3686_ _1155_ _1231_ _1246_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2706_ _0363_ _0364_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or2_1
X_2637_ _0300_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__buf_12
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2568_ _0236_ _0251_ _0252_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__and3_1
X_2499_ _1872_ d11.count\[3\] _0198_ _0199_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__a211o_1
X_4307_ clknet_leaf_22_clk _0040_ net33 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
X_4238_ clknet_leaf_32_clk _0011_ net27 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4169_ d9.count\[8\] _1715_ _1718_ d9.count\[7\] _2017_ vssd1 vssd1 vccd1 vccd1 _1694_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3540_ _0915_ _0988_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3471_ d6.saw_temp\[7\] _0926_ _0728_ d6.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _1035_
+ sky130_fd_sc_hd__o22a_1
X_2422_ net76 _2023_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
X_2353_ d7.count\[3\] d7.count\[4\] _1963_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__and3_1
X_4023_ _1469_ _1539_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__or2b_1
X_2284_ _1735_ _1912_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3807_ _1363_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3738_ _0620_ _1181_ _1188_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__nor3_1
X_3669_ _1157_ _1137_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__or2b_1
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2971_ d1.saw_temp\[4\] d1.saw_temp\[3\] d1.saw_temp\[0\] _0561_ vssd1 vssd1 vccd1
+ vccd1 _0562_ sky130_fd_sc_hd__nand4_1
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3523_ _1085_ _1086_ _0646_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__mux2_1
X_3454_ _0999_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__xnor2_1
X_2405_ _2008_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_3385_ _0945_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__xor2_2
X_2336_ d7.count\[6\] _1733_ _1954_ _1955_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__a211oi_1
X_2267_ d5.count\[5\] d5.count\[4\] _1895_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4006_ _1518_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__inv_2
X_2198_ _1712_ _1844_ d4.count\[4\] d4.count\[5\] d4.count\[3\] vssd1 vssd1 vccd1
+ vccd1 _1845_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold31 d5.count\[0\] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 d13.count\[0\] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 d4.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 d13.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0128_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 d12.count\[6\] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 d6.count\[6\] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 p0.count\[2\] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _0695_ _0696_ _0734_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__o21a_1
X_2121_ _1786_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2052_ _1712_ _1727_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2954_ d8.saw_temp\[5\] _0545_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2885_ d6.saw_temp\[7\] _0499_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3506_ _0560_ d1.saw_temp\[2\] _0330_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand3_1
X_4486_ clknet_leaf_8_clk _0145_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_2
X_3437_ d5.saw_temp\[7\] _0897_ _0744_ d5.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _1001_
+ sky130_fd_sc_hd__o22a_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__nand2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _1940_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_3299_ _0861_ _0864_ _0634_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2670_ net3 vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__clkbuf_8
X_4340_ clknet_leaf_29_clk d8.nxt_count\[7\] net28 vssd1 vssd1 vccd1 vccd1 d8.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4271_ clknet_leaf_21_clk _0024_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
X_3222_ d4.saw_temp\[1\] _0347_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__nand2_1
X_3153_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__inv_2
X_2104_ d2.count\[3\] _1733_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3084_ d12.saw_temp\[6\] _0648_ _0649_ _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or4b_2
X_2035_ d1.oct_dwn\[1\] vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3986_ _1434_ _1447_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__a21o_1
X_2937_ _0534_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2868_ d5.saw_temp\[3\] _0481_ _0484_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2799_ d3.count\[0\] _1732_ _1812_ _1815_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4469_ clknet_leaf_18_clk net93 net38 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _0622_ _1400_ _0620_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3771_ _1327_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2722_ _0358_ _0361_ _0379_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2653_ p0.count\[3\] vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2584_ net71 _0266_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4323_ clknet_leaf_31_clk d7.nxt_count\[8\] net31 vssd1 vssd1 vccd1 vccd1 d7.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_4254_ clknet_leaf_33_clk _0017_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_4
X_4185_ d9.saw_temp\[5\] _1703_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3205_ d3.saw_temp\[6\] _0769_ _0770_ _0771_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__or4b_2
X_3136_ _0683_ _0702_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nor2_1
X_3067_ _0618_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__buf_8
XFILLER_0_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3969_ _1411_ _1415_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold161 d4.count\[6\] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 d12.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 d10.count\[4\] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 d11.count\[4\] vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 em0.u1.state\[2\] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3823_ _1382_ _1383_ _0683_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3754_ _1313_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__xnor2_2
X_3685_ _1155_ _1231_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__a21oi_1
X_2705_ _0331_ _0332_ _0363_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__o2bb2a_1
X_2636_ s0.type_switch\[0\] vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2567_ d12.count\[6\] _0247_ d12.count\[7\] vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2498_ _1872_ d11.count\[3\] d11.count\[2\] vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__o21a_1
X_4306_ clknet_leaf_3_clk net49 net26 vssd1 vssd1 vccd1 vccd1 d6.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4237_ clknet_leaf_32_clk _0010_ net27 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_4168_ _1727_ d9.count\[6\] d9.count\[3\] vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__a21boi_1
X_3119_ d9.saw_temp\[5\] _0335_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__nand2_1
X_4099_ _1592_ _1593_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3470_ d6.saw_temp\[3\] _0346_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nand2_1
X_2421_ d9.count\[8\] _1805_ _2022_ d9.count\[9\] vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__a211oi_4
X_2352_ _1968_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_2283_ _1872_ d6.count\[5\] d6.count\[4\] vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__a21o_1
X_4022_ _1558_ _1580_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3806_ _0749_ _1366_ _0708_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3737_ _1297_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3668_ _1125_ _1130_ _1124_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__a21bo_1
X_3599_ _0622_ _1160_ _1161_ _0659_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__a31o_1
X_2619_ net132 _0287_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2970_ d1.saw_temp\[6\] d1.saw_temp\[5\] d1.saw_temp\[2\] d1.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3522_ d12.saw_temp\[7\] _0977_ _0871_ d12.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1
+ _1086_ sky130_fd_sc_hd__o22a_1
X_3453_ _1015_ _1016_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__nor2_1
X_2404_ _1990_ _2006_ _2007_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__and3_1
X_3384_ _0622_ _0948_ _0669_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__a21o_1
X_2335_ _1721_ d7.count\[7\] vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2266_ _1898_ _1899_ vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
X_4005_ _1562_ _1563_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__and2_1
X_2197_ d4.count\[7\] vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold32 d5.nxt_count\[0\] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 d13.nxt_count\[0\] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 em0.u1.R\[12\] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 d7.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 d5.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 em0.u1.D\[9\] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 d6.count\[4\] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 d12.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _0288_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2120_ _1783_ _1784_ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__and3_1
X_2051_ _1727_ d1.count\[4\] _1718_ d1.count\[5\] vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2953_ d8.saw_temp\[5\] _0545_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2884_ d6.saw_temp\[4\] d6.saw_temp\[3\] d6.saw_temp\[0\] _0498_ vssd1 vssd1 vccd1
+ vccd1 _0499_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3505_ d1.saw_temp\[3\] _0330_ _0300_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__a21oi_1
X_4485_ clknet_leaf_8_clk _0144_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_1
X_3436_ d5.saw_temp\[3\] _0328_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__nand2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _0925_ _0930_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__or2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _1922_ _1938_ _1939_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3298_ _0862_ _0863_ d13.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__mux2_1
X_2249_ d5.count\[8\] _1805_ _1871_ _1886_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ clknet_leaf_27_clk net51 net28 vssd1 vssd1 vccd1 vccd1 d4.count\[9\] sky130_fd_sc_hd__dfrtp_2
X_3221_ _0751_ _0786_ _0747_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__a21boi_1
X_3152_ _0717_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__nor2_1
X_2103_ _1735_ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__nor2_1
X_3083_ d12.saw_temp\[5\] _0340_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__nand2_1
X_2034_ _1710_ _1711_ net245 vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _1448_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2936_ d8.count\[3\] _1718_ _1777_ d8.count\[1\] vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__a2bb2o_1
X_2867_ d5.saw_temp\[3\] _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2798_ _1735_ d3.count\[1\] d3.count\[5\] _1810_ _1813_ vssd1 vssd1 vccd1 vccd1 _0437_
+ sky130_fd_sc_hd__a2111o_1
X_4468_ clknet_leaf_17_clk _0127_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[0\] sky130_fd_sc_hd__dfrtp_1
X_3419_ _0880_ _0882_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__and2b_1
X_4399_ clknet_leaf_2_clk d11.nxt_count\[8\] net26 vssd1 vssd1 vccd1 vccd1 d11.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3770_ _1222_ _1224_ _1328_ _1329_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2721_ _0358_ _0361_ _0379_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2652_ p0.count\[5\] vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__inv_2
X_2583_ d13.count\[8\] _1805_ _0255_ _0265_ d13.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _0266_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ clknet_leaf_31_clk d7.nxt_count\[7\] net31 vssd1 vssd1 vccd1 vccd1 d7.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4253_ clknet_leaf_33_clk _0016_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
X_3204_ d3.saw_temp\[5\] _0348_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__nand2_1
X_4184_ _1703_ net166 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__nor2_1
X_3135_ _0697_ _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__nand2_2
X_3066_ d13.saw_temp\[7\] _0301_ _0344_ _0307_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__a31o_2
XFILLER_0_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3968_ _1523_ _1527_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__xnor2_2
X_2919_ d7.saw_temp\[3\] _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__nand2_1
X_3899_ d3.saw_temp\[6\] _0348_ _0772_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold162 d1.count\[3\] vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 d13.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 d6.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 d4.count\[7\] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 d2.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 d3.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3822_ d11.saw_temp\[6\] _0334_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3753_ _1175_ _1176_ _1205_ _1314_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3684_ _1242_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__xnor2_1
X_2704_ _0333_ _0362_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__and2_1
X_2635_ _1724_ _0297_ _0298_ _1726_ vssd1 vssd1 vccd1 vccd1 e0.next_q\[1\] sky130_fd_sc_hd__a22o_1
X_2566_ d12.count\[7\] d12.count\[6\] _0247_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__nand3_1
X_4305_ clknet_leaf_3_clk d6.nxt_count\[8\] net26 vssd1 vssd1 vccd1 vccd1 d6.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2497_ _0195_ _1729_ _0196_ _0197_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4236_ clknet_leaf_33_clk _0009_ net27 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_4167_ _1735_ d9.count\[1\] d9.count\[8\] _1715_ d9.count\[9\] vssd1 vssd1 vccd1
+ vccd1 _1692_ sky130_fd_sc_hd__a221o_1
X_3118_ d9.saw_temp\[0\] d9.saw_temp\[3\] _0335_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__o21a_1
X_4098_ _0893_ _1647_ _1649_ _1653_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__o31a_1
X_3049_ _0610_ _0611_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2420_ d9.count\[8\] _1805_ _1720_ d9.count\[7\] _2021_ vssd1 vssd1 vccd1 vccd1 _2022_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_51_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2351_ _1966_ _1967_ _1959_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2282_ _1721_ d6.count\[7\] d6.count\[6\] vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__o21ai_1
X_4021_ _1578_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3805_ _1364_ _1365_ _0682_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3736_ _1063_ _1291_ _1296_ _1064_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3667_ _1114_ _1134_ _1132_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21o_1
X_3598_ d11.saw_temp\[4\] _0334_ _0682_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__nand3_1
X_2618_ p0.count\[3\] _0287_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__and2_1
X_2549_ _0239_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_4219_ clknet_leaf_34_clk d1.nxt_count\[9\] net25 vssd1 vssd1 vccd1 vccd1 d1.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3521_ d12.saw_temp\[3\] _0340_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3452_ _0934_ _0940_ _1014_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__and3_1
X_3383_ _0946_ _0947_ _0618_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__mux2_1
X_2403_ d8.count\[7\] _2004_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__or2_1
X_2334_ d7.count\[6\] _1733_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__o21a_1
X_2265_ d5.count\[4\] _1895_ _1888_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4004_ _1559_ _1503_ _1561_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__nand3_1
X_2196_ _1713_ d4.count\[0\] d4.count\[1\] _1721_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3719_ _0686_ _1280_ _0646_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold22 d3.count\[0\] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 _0101_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 em0.u1.count\[1\] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 d12.count\[0\] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 em0.u1.R\[9\] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 d10.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 em0.u1.R\[22\] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 d3.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 d6.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2050_ _1716_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__buf_6
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2952_ _0545_ _0546_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__nor2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2883_ d6.saw_temp\[6\] d6.saw_temp\[5\] d6.saw_temp\[2\] d6.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4484_ clknet_leaf_8_clk _0143_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3504_ _1065_ _1067_ _0306_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3435_ _0905_ _0910_ _0904_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__a21bo_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _0925_ _0930_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__nand2_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ d6.count\[7\] _1936_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__or2_1
X_3297_ d13.saw_temp\[7\] _0345_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__or2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _1873_ _1883_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2179_ d3.count\[4\] d3.count\[5\] _1827_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3220_ _0783_ _0785_ _0760_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__mux2_1
X_3151_ _0706_ _0716_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__and2_1
X_2102_ _1713_ d2.count\[1\] d2.count\[2\] vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3082_ d12.saw_temp\[3\] d12.saw_temp\[0\] _0340_ vssd1 vssd1 vccd1 vccd1 _0649_
+ sky130_fd_sc_hd__o21a_1
X_2033_ net102 em0.u1.count\[1\] net60 vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__nand3_1
X_3984_ _1540_ _1543_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2935_ d8.count\[3\] _1718_ _1723_ d8.count\[2\] vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2866_ net222 _0486_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__nor2_1
X_2797_ d3.count\[2\] _1733_ _1807_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4467_ clknet_leaf_23_clk _0126_ net33 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4398_ clknet_leaf_2_clk d11.nxt_count\[7\] net26 vssd1 vssd1 vccd1 vccd1 d11.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3418_ _0955_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__xor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ _0912_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__nor2_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2720_ _0377_ _0378_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__or2_1
X_2651_ _0312_ em0.mixed_sample\[6\] vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2582_ _0256_ _0264_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4321_ clknet_leaf_30_clk d7.nxt_count\[6\] net29 vssd1 vssd1 vccd1 vccd1 d7.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4252_ clknet_leaf_24_clk d3.nxt_count\[9\] net32 vssd1 vssd1 vccd1 vccd1 d3.count\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3203_ d3.saw_temp\[3\] d3.saw_temp\[0\] _0348_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__o21a_1
X_4183_ d9.saw_temp\[3\] _1701_ net165 vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3134_ d8.saw_temp\[6\] _0698_ _0699_ _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__or4b_2
X_3065_ _0621_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__xor2_2
XFILLER_0_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3967_ _0310_ _1526_ _0645_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__o21a_1
X_2918_ net180 _0520_ _0522_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_30_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3898_ _1453_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2849_ _0456_ _0461_ d4.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__a21oi_1
Xhold141 d7.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 d7.count\[4\] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 d3.count\[3\] vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 d10.count\[5\] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 d8.count\[4\] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 p0.count\[4\] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 d11.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ d11.saw_temp\[7\] _0662_ _0664_ d11.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1
+ _1382_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3752_ _1204_ _1202_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__and2b_1
X_3683_ _0751_ _1244_ _0767_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2703_ _0333_ _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__nor2_1
X_2634_ _0298_ _0299_ vssd1 vssd1 vccd1 vccd1 e0.next_q\[0\] sky130_fd_sc_hd__nand2_1
X_2565_ net137 _0247_ _0250_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[6\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4304_ clknet_leaf_3_clk d6.nxt_count\[7\] net26 vssd1 vssd1 vccd1 vccd1 d6.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2496_ d11.count\[2\] _1723_ _1777_ d11.count\[1\] vssd1 vssd1 vccd1 vccd1 _0197_
+ sky130_fd_sc_hd__o22a_1
X_4235_ clknet_leaf_31_clk _0008_ net31 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_4166_ d9.saw_temp\[7\] _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3117_ d9.saw_temp\[4\] d9.saw_temp\[1\] d9.saw_temp\[2\] _0335_ vssd1 vssd1 vccd1
+ vccd1 _0684_ sky130_fd_sc_hd__o31a_1
X_4097_ em0.u1.R\[19\] _1633_ _1652_ _0326_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__o22a_1
X_3048_ d2.saw_temp\[6\] _0612_ _0613_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4382__45 vssd1 vssd1 vccd1 vccd1 _4382__45/HI net45 sky130_fd_sc_hd__conb_1
XFILLER_0_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2350_ d7.count\[3\] _1963_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__or2_1
X_2281_ _1721_ _1909_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__nand2_1
X_4020_ _1575_ _1577_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3804_ d7.saw_temp\[6\] net12 vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__nand2_1
X_3735_ _1063_ _1064_ _1291_ _1296_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3666_ _1111_ _1217_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__nand2_1
X_3597_ _0682_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2617_ _0287_ net127 vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2548_ _0236_ _0237_ _0238_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2479_ d10.count\[5\] d10.count\[4\] _0179_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__and3_1
X_4218_ clknet_leaf_33_clk net110 net25 vssd1 vssd1 vccd1 vccd1 d1.count\[8\] sky130_fd_sc_hd__dfrtp_4
X_4149_ net188 net63 em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3520_ _1078_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__xor2_2
X_3451_ _0934_ _0940_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__a21oi_1
X_3382_ d10.saw_temp\[7\] _0833_ _0674_ d10.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1
+ _0947_ sky130_fd_sc_hd__o22a_1
X_2402_ d8.count\[7\] _2004_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__nand2_1
X_2333_ d7.count\[5\] _1944_ _1947_ _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__a22o_1
X_2264_ d5.count\[3\] d5.count\[4\] _1892_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4003_ _1559_ _1503_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__a21o_1
X_2195_ d4.count\[6\] _1725_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3718_ _0688_ _0840_ d9.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__mux2_1
X_3649_ _1043_ _1097_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold23 d4.count\[0\] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 em0.u1.Q\[7\] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _0136_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 d7.count\[0\] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 em0.u1.R\[10\] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 d8.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 d5.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 d6.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2951_ d8.saw_temp\[3\] _0543_ net167 vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__a21oi_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2882_ _1918_ _1921_ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and3b_1
XFILLER_0_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4483_ clknet_leaf_8_clk _0142_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
X_3503_ d2.saw_temp\[2\] _0611_ _0615_ _1066_ _0618_ vssd1 vssd1 vccd1 vccd1 _1067_
+ sky130_fd_sc_hd__o311a_1
X_3434_ _0896_ _0914_ _0912_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__a21oi_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__inv_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ d6.count\[7\] _1936_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__nand2_1
X_3296_ _0635_ _0639_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__nand2_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _1725_ _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2178_ _1829_ _1830_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_0_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3150_ _0706_ _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nor2_1
X_2101_ d2.count\[7\] _1722_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__nand2_1
X_3081_ d12.saw_temp\[4\] d12.saw_temp\[2\] d12.saw_temp\[1\] _0340_ vssd1 vssd1 vccd1
+ vccd1 _0648_ sky130_fd_sc_hd__o31a_1
X_2032_ em0.u1.state\[1\] vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3983_ _1357_ _1541_ _1542_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2934_ d8.count\[6\] _1733_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a21oi_1
X_2865_ _0481_ _0484_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__and2_1
X_2796_ net239 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4466_ clknet_leaf_22_clk _0125_ net33 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4397_ clknet_leaf_2_clk d11.nxt_count\[6\] net26 vssd1 vssd1 vccd1 vccd1 d11.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3417_ _0980_ _0981_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__xor2_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3348_ _0823_ _0826_ _0911_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__and3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _0838_ _0844_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4400__44 vssd1 vssd1 vccd1 vccd1 _4400__44/HI net44 sky130_fd_sc_hd__conb_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2650_ p0.count\[6\] vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2581_ d13.count\[6\] _1723_ _1726_ d13.count\[5\] _0263_ vssd1 vssd1 vccd1 vccd1
+ _0264_ sky130_fd_sc_hd__o221a_1
X_4320_ clknet_leaf_35_clk d7.nxt_count\[5\] net25 vssd1 vssd1 vccd1 vccd1 d7.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4251_ clknet_leaf_24_clk d3.nxt_count\[8\] net32 vssd1 vssd1 vccd1 vccd1 d3.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3202_ d3.saw_temp\[4\] d3.saw_temp\[2\] d3.saw_temp\[1\] _0348_ vssd1 vssd1 vccd1
+ vccd1 _0769_ sky130_fd_sc_hd__o31a_1
X_4182_ d9.saw_temp\[4\] d9.saw_temp\[3\] _1701_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__and3_1
X_3133_ d8.saw_temp\[5\] _0337_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__nand2_1
X_3064_ _0622_ _0628_ _0629_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3966_ _0738_ _0647_ _1418_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__o31ai_1
X_2917_ _0514_ _0517_ d7.saw_temp\[2\] d7.saw_temp\[1\] d7.saw_temp\[0\] vssd1 vssd1
+ vccd1 vccd1 _0522_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3897_ _0310_ _1455_ _1456_ _0762_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2848_ net130 _0470_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__xnor2_1
X_2779_ net235 _0421_ _0425_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__o21a_1
Xhold153 d9.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 d10.count\[6\] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 d4.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 d6.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ clknet_leaf_27_clk d13.nxt_count\[7\] net29 vssd1 vssd1 vccd1 vccd1 d13.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold186 d7.count\[5\] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 d13.count\[4\] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 p0.nxt_count\[4\] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 d2.count\[3\] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3820_ _1379_ _1380_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__and2_1
X_3751_ _1286_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__xor2_2
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2702_ _0360_ _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3682_ _0771_ _1243_ _0760_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__mux2_1
X_2633_ _1872_ _0297_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__or2_1
X_2564_ d12.count\[6\] _0247_ _0236_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4303_ clknet_leaf_1_clk d6.nxt_count\[6\] net22 vssd1 vssd1 vccd1 vccd1 d6.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2495_ _1872_ d11.count\[3\] vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__xor2_1
X_4234_ clknet_leaf_26_clk d2.nxt_count\[9\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4165_ d9.saw_temp\[6\] d9.saw_temp\[0\] d9.saw_temp\[3\] _1689_ vssd1 vssd1 vccd1
+ vccd1 _1690_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3116_ _0682_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__buf_6
X_4096_ em0.u1.R\[18\] _1651_ _1609_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3047_ d2.saw_temp\[2\] d2.saw_temp\[1\] _0329_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3949_ _0749_ _1507_ _1508_ _0620_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4288__50 vssd1 vssd1 vccd1 vccd1 _4288__50/HI net50 sky130_fd_sc_hd__conb_1
XFILLER_0_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2280_ _1727_ d6.count\[6\] d6.count\[7\] vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3803_ d7.saw_temp\[7\] _0711_ _0713_ d7.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 _1364_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3734_ _0622_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3665_ _0779_ _1225_ _1226_ _1227_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__a31o_1
X_2616_ p0.count\[1\] p0.count\[0\] net126 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a21oi_1
X_3596_ d11.saw_temp\[7\] _1044_ _0664_ d11.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1
+ _1159_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2547_ d12.count\[1\] d12.count\[0\] vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__or2_1
X_2478_ _0182_ _0183_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4217_ clknet_leaf_35_clk d1.nxt_count\[7\] net25 vssd1 vssd1 vccd1 vccd1 d1.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_4148_ _1685_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _1620_ _1621_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3450_ _1009_ _1013_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__xnor2_1
X_3381_ d10.saw_temp\[2\] _0336_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__nand2_1
X_2401_ _2004_ _2005_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
X_2332_ _1948_ _1951_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__nand2_1
X_4002_ _0722_ _1480_ _1483_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__o31a_1
X_2263_ _1897_ vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_2194_ d4.count\[6\] _1725_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3717_ _1277_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3648_ _1096_ _1094_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__and2b_1
X_3579_ d7.saw_temp\[7\] _1027_ _0713_ d7.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 _1142_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold13 _0134_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 d10.count\[0\] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 d4.nxt_count\[0\] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _0099_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 d9.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 d4.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 d1.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ d8.saw_temp\[4\] d8.saw_temp\[3\] _0543_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__and3_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ d6.count\[3\] _1777_ _1919_ _1923_ d6.count\[2\] vssd1 vssd1 vccd1 vccd1 _0496_
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4482_ clknet_leaf_8_clk _0141_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3502_ d2.saw_temp\[7\] d2.saw_temp\[2\] _0329_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__nand3b_1
X_3433_ _0779_ _0995_ _0996_ _0997_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _0749_ _0928_ _0722_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__a21o_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _1936_ _1937_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
X_3295_ d13.saw_temp\[1\] _0344_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__nand2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _1721_ d5.count\[7\] d5.count\[6\] vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2177_ net232 _1827_ _1819_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2100_ d2.count\[9\] _1714_ _1718_ d2.count\[8\] vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__a22o_1
X_3080_ d12.saw_temp\[7\] _0340_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__and2_2
X_2031_ _1709_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _1429_ _1431_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__nor2_1
X_2933_ d8.count\[8\] _1715_ _1980_ d8.count\[9\] vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2864_ d5.saw_temp\[1\] _0484_ net221 vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__a21oi_1
X_2795_ _0424_ _0434_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ clknet_leaf_22_clk _0124_ net33 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4396_ clknet_leaf_34_clk d11.nxt_count\[5\] net34 vssd1 vssd1 vccd1 vccd1 d11.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3416_ _0868_ _0877_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__and2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ _0823_ _0826_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__a21oi_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3278_ _0843_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2229_ _1868_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2580_ d13.count\[4\] _1720_ _1726_ d13.count\[5\] _0262_ vssd1 vssd1 vccd1 vccd1
+ _0263_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4250_ clknet_leaf_24_clk d3.nxt_count\[7\] net32 vssd1 vssd1 vccd1 vccd1 d3.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4181_ net125 _1701_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__xor2_1
X_3201_ d3.saw_temp\[7\] _0348_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__and2_1
X_3132_ d8.saw_temp\[0\] d8.saw_temp\[3\] _0337_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3063_ d1.saw_temp\[7\] _0300_ _0330_ _0306_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _0647_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__nand2_1
X_2916_ _0520_ _0521_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__nor2_1
X_3896_ d4.saw_temp\[7\] d4.saw_temp\[6\] _0347_ _0760_ vssd1 vssd1 vccd1 vccd1 _1456_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2847_ _0472_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2778_ _0424_ _0421_ d2.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__o21ai_2
Xhold110 d4.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 d10.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 d5.count\[5\] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 d1.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 d8.count\[6\] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 d9.count\[5\] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ clknet_leaf_27_clk d13.nxt_count\[6\] net29 vssd1 vssd1 vccd1 vccd1 d13.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold165 d8.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 d1.count\[6\] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 d3.count\[6\] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlygate4sd3_1
X_4379_ clknet_leaf_1_clk d10.nxt_count\[6\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3750_ _1310_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__xnor2_2
X_2701_ _0334_ _0359_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3681_ _0793_ _0794_ d3.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2632_ _1872_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2563_ _0249_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4302_ clknet_leaf_1_clk d6.nxt_count\[5\] net22 vssd1 vssd1 vccd1 vccd1 d6.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4233_ clknet_leaf_26_clk d2.nxt_count\[8\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2494_ d11.count\[2\] vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4164_ d9.saw_temp\[5\] d9.saw_temp\[4\] d9.saw_temp\[1\] d9.saw_temp\[2\] vssd1
+ vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__and4_1
XFILLER_0_65_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3115_ _0640_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__clkbuf_8
X_4095_ _1602_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3046_ d2.saw_temp\[0\] _0329_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3948_ d2.saw_temp\[7\] _0682_ _1399_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__or3_1
X_3879_ _1437_ _1439_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3802_ _0705_ _1362_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__nand2_1
X_3733_ _0640_ _1292_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3664_ em0.u1.state\[1\] em0.u1.R\[11\] net61 _0781_ vssd1 vssd1 vccd1 vccd1 _1227_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2615_ p0.count\[2\] p0.count\[1\] p0.count\[0\] vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__and3_1
X_3595_ _1137_ _1157_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2546_ d12.count\[1\] d12.count\[0\] vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__nand2_1
X_2477_ net223 _0179_ _0172_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__o21ai_1
X_4216_ clknet_leaf_35_clk d1.nxt_count\[6\] net25 vssd1 vssd1 vccd1 vccd1 d1.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4147_ net187 net88 em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__mux2_1
X_4078_ _1562_ _1619_ _1616_ _1569_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3029_ _0600_ _0601_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2400_ net227 _2002_ _1990_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__o21ai_1
X_3380_ _0622_ _0944_ _0659_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2331_ d7.count\[1\] _1949_ _1950_ d7.count\[3\] _1948_ vssd1 vssd1 vccd1 vccd1 _1951_
+ sky130_fd_sc_hd__o221ai_1
X_2262_ _1895_ _1896_ _1888_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__and3b_1
X_4001_ _1475_ _1479_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__or2b_1
X_2193_ _1840_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3716_ _1273_ _1276_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3647_ _1158_ _1209_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__xnor2_2
X_3578_ _1139_ _1140_ _0705_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2529_ _0222_ _0223_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
Xhold14 d11.count\[0\] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 d2.count\[8\] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 d9.count\[0\] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 d3.count\[8\] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 d10.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 d1.count\[8\] vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ _0495_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4481_ clknet_leaf_8_clk _0140_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3501_ d2.saw_temp\[3\] _0329_ _0300_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3432_ em0.u1.state\[1\] net95 net96 _0781_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__a22o_1
X_3363_ _0926_ _0927_ _0634_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__mux2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ net148 _1933_ _1922_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__o21ai_1
X_3294_ _0857_ _0858_ _0848_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__a21o_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _1876_ _1877_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__a21oi_1
X_2176_ d3.count\[3\] d3.count\[4\] _1823_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2030_ em0.u1.state\[3\] em0.u1.state\[0\] vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__or2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3981_ _1429_ _1431_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__nand2_1
X_2932_ d8.saw_temp\[7\] _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2863_ net118 _0484_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__xor2_1
X_2794_ _0423_ _0421_ d2.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4464_ clknet_leaf_19_clk _0123_ net39 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4395_ clknet_leaf_34_clk d11.nxt_count\[4\] net34 vssd1 vssd1 vccd1 vccd1 d11.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3415_ _0974_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__xor2_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _0906_ _0910_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__xnor2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _0622_ _0842_ _0681_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _1850_ _1866_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__and3_1
X_2159_ d3.count\[5\] _1814_ _1815_ _1777_ d3.count\[6\] vssd1 vssd1 vccd1 vccd1 _1816_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4180_ _1701_ _1702_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__nor2_1
X_3200_ d3.saw_temp\[7\] _0301_ _0348_ _0307_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__a31o_2
X_3131_ d8.saw_temp\[4\] d8.saw_temp\[1\] d8.saw_temp\[2\] _0337_ vssd1 vssd1 vccd1
+ vccd1 _0698_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3062_ _0618_ _0625_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3964_ _0651_ _1418_ _0723_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__a21o_1
X_2915_ _0519_ _0518_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3895_ _0738_ _1454_ _0753_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__o21a_1
X_2846_ _0470_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold100 d9.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dlygate4sd3_1
X_2777_ d2.saw_temp\[7\] _0423_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__and2_1
Xhold122 d7.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold111 d5.count\[6\] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _1901_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold133 d3.count\[5\] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 d5.count\[9\] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_1
X_4447_ clknet_leaf_30_clk d13.nxt_count\[5\] net29 vssd1 vssd1 vccd1 vccd1 d13.count\[5\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold155 d6.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _0544_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 d1.count\[4\] vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold188 d3.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__dlygate4sd3_1
X_4378_ clknet_leaf_37_clk d10.nxt_count\[5\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _1710_ net66 _0782_ net95 vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2700_ _0334_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or2_1
X_3680_ _1240_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ net220 m0.edgy.in vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__or2b_1
X_2562_ _0247_ _0248_ _0236_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__and3b_1
X_4301_ clknet_leaf_1_clk d6.nxt_count\[4\] net22 vssd1 vssd1 vccd1 vccd1 d6.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_4232_ clknet_leaf_26_clk d2.nxt_count\[7\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2493_ _1713_ d11.count\[4\] d11.count\[5\] vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_4_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4163_ _0326_ _1711_ _1687_ net60 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__o22a_1
X_4094_ em0.u1.D\[11\] em0.u1.R\[18\] vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__xor2_1
X_3114_ _0301_ _0680_ _0307_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__a21oi_4
X_3045_ d2.saw_temp\[5\] d2.saw_temp\[4\] d2.saw_temp\[3\] net7 vssd1 vssd1 vccd1
+ vccd1 _0612_ sky130_fd_sc_hd__o31a_1
XFILLER_0_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3947_ _0634_ _0615_ _1506_ _0611_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3878_ _1229_ _1325_ _1438_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__a21boi_1
X_2829_ _1735_ d4.count\[1\] _1869_ _1724_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3801_ _0682_ _1359_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3732_ d1.saw_temp\[4\] _0623_ _0627_ _1293_ _0618_ vssd1 vssd1 vccd1 vccd1 _1294_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3663_ _1222_ _1224_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2614_ net134 net90 vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[1\] sky130_fd_sc_hd__xor2_1
X_3594_ _1155_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2545_ net84 _0236_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2476_ d10.count\[3\] d10.count\[4\] _0176_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__and3_1
X_4215_ clknet_leaf_35_clk d1.nxt_count\[5\] net25 vssd1 vssd1 vccd1 vccd1 d1.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4146_ _1684_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
X_4077_ _1634_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
X_3028_ d11.saw_temp\[2\] d11.saw_temp\[1\] _0599_ vssd1 vssd1 vccd1 vccd1 _0601_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2330_ _1727_ d7.count\[2\] vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__and2_1
X_2261_ d5.count\[3\] _1892_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__or2_1
X_4000_ _1493_ _1497_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__or2b_1
X_2192_ _1819_ _1838_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3715_ _1273_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3646_ _1206_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__xor2_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3577_ d8.saw_temp\[4\] _0337_ _0682_ _0310_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2528_ net159 _0220_ _0208_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__o21ai_1
X_2459_ _1872_ _0163_ _0165_ _0168_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__o211a_1
Xhold26 d9.nxt_count\[0\] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 em0.u1.Q\[6\] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 em0.u1.R\[8\] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 d11.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 d1.nxt_count\[8\] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dlygate4sd3_1
X_4129_ _1675_ _1676_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3500_ d1.saw_temp\[7\] _0300_ _0330_ _0306_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a31o_2
X_4480_ clknet_leaf_8_clk _0139_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3431_ _0892_ _0994_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3362_ d6.saw_temp\[7\] _0817_ _0728_ d6.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0927_
+ sky130_fd_sc_hd__o22a_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ d6.count\[6\] _1933_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__and2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _0848_ _0857_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__nand3_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _1881_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__inv_2
X_2175_ _1827_ _1828_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_79_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3629_ _1189_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__xor2_4
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _1469_ _1539_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__xnor2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2931_ d8.saw_temp\[6\] d8.saw_temp\[0\] d8.saw_temp\[3\] _0529_ vssd1 vssd1 vccd1
+ vccd1 _0530_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2862_ net196 _0479_ _0484_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2793_ net123 _0432_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4463_ clknet_leaf_19_clk _0122_ net39 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3414_ _0976_ _0978_ _0645_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__o21ai_1
X_4394_ clknet_leaf_34_clk d11.nxt_count\[3\] net25 vssd1 vssd1 vccd1 vccd1 d11.count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3345_ _0751_ _0909_ _0767_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__a21boi_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3276_ _0839_ _0841_ _0634_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__mux2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ d4.count\[7\] _1864_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__or2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2158_ d3.count\[4\] _1714_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__and2_1
X_2089_ net238 _1757_ _1745_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3130_ d8.saw_temp\[7\] _0337_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__and2_1
X_3061_ _0610_ _0623_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3963_ _1518_ _1522_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__xor2_2
X_2914_ _0519_ _0518_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nor2_1
X_3894_ d4.saw_temp\[6\] _0347_ _0758_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2845_ d4.saw_temp\[5\] _0468_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__or2_1
Xhold101 d4.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ d2.saw_temp\[4\] d2.saw_temp\[3\] d2.saw_temp\[0\] _0422_ vssd1 vssd1 vccd1
+ vccd1 _0423_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 _1903_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 d12.count\[8\] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 d2.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ clknet_leaf_30_clk d13.nxt_count\[4\] net29 vssd1 vssd1 vccd1 vccd1 d13.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold156 d2.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 d2.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 d5.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ clknet_leaf_37_clk d10.nxt_count\[4\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold189 d9.count\[6\] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 d5.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _0780_ _0891_ _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__a21o_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _0823_ _0824_ _0717_ _0732_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2630_ net81 _0294_ vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[7\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2561_ d12.count\[4\] _0243_ d12.count\[5\] vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4300_ clknet_leaf_3_clk d6.nxt_count\[3\] net26 vssd1 vssd1 vccd1 vccd1 d6.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2492_ _1727_ d11.count\[6\] _1718_ d11.count\[7\] vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ clknet_leaf_26_clk d2.nxt_count\[6\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _1687_ _1688_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__nor2_1
X_3113_ d9.saw_temp\[7\] _0335_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__and2_2
X_4093_ _1648_ _1641_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3044_ d2.saw_temp\[7\] _0329_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3946_ _0640_ _1399_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3877_ _1324_ _1321_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2828_ d4.count\[2\] _1724_ _1777_ d4.count\[0\] vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2759_ d13.saw_temp\[3\] _0409_ net210 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__a21oi_1
X_4429_ clknet_leaf_20_clk _0098_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout40 net16 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_6
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _0634_ _1360_ _0622_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__o21a_1
X_4451__42 vssd1 vssd1 vccd1 vccd1 _4451__42/HI net42 sky130_fd_sc_hd__conb_1
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3731_ d1.saw_temp\[4\] _1183_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3662_ _1222_ _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__nand2_1
X_3593_ _1052_ _1060_ _1154_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__nand3_1
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2613_ net90 vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[0\] sky130_fd_sc_hd__inv_2
X_2544_ _0229_ _0235_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__nor2_2
X_2475_ _0181_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4214_ clknet_leaf_35_clk d1.nxt_count\[4\] net24 vssd1 vssd1 vccd1 vccd1 d1.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4145_ em0.mixed_sample\[5\] net208 em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1 _1684_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ em0.u1.R\[17\] _1632_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3027_ d11.saw_temp\[1\] _0599_ d11.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _0600_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3929_ _1470_ _1488_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2260_ d5.count\[3\] _1892_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__and2_1
X_2191_ d3.count\[9\] d3.count\[8\] _1835_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3714_ _0749_ _1275_ _0669_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3645_ _1062_ _1093_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3576_ _0683_ _1138_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nor2_1
X_2527_ d11.count\[6\] _0220_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__and2_1
X_2458_ d10.count\[5\] _1729_ _0164_ _0167_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold16 em0.u1.R\[21\] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 _0133_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 em0.u1.Q\[2\] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold49 d12.count\[4\] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ d8.count\[3\] _1994_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__and2_1
X_4128_ d12.saw_temp\[3\] _1673_ net176 vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__a21oi_1
X_4059_ _1569_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3430_ _0892_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3361_ d6.saw_temp\[2\] _0346_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2312_ _1935_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _0620_ _0852_ _0856_ _0630_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _1878_ _1879_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__a21oi_1
X_2174_ net203 _1823_ _1819_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3628_ _0956_ _0967_ _1075_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__a31o_2
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 PWM_o sky130_fd_sc_hd__clkbuf_4
X_3559_ d4.saw_temp\[4\] _0347_ _0683_ _0310_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__a31o_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2930_ d8.saw_temp\[5\] d8.saw_temp\[4\] d8.saw_temp\[1\] d8.saw_temp\[2\] vssd1
+ vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2861_ _0483_ _0478_ d5.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2792_ _0433_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4462_ clknet_leaf_19_clk _0121_ net39 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3413_ _0760_ _0977_ _0750_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__o21ai_1
X_4393_ clknet_leaf_37_clk d11.nxt_count\[2\] net23 vssd1 vssd1 vccd1 vccd1 d11.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3344_ _0907_ _0908_ _0760_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _0688_ _0840_ d9.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2226_ net246 _1864_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__nand2_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2157_ _1809_ _1811_ _1812_ _1813_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__a211oi_1
X_2088_ d1.count\[6\] _1757_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3060_ d1.saw_temp\[6\] _0624_ _0625_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3962_ _0751_ _1520_ _1521_ _0866_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__a31o_1
X_2913_ d7.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3893_ _1451_ _1452_ _0747_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__o21a_1
X_2844_ d4.saw_temp\[5\] _0468_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2775_ d2.saw_temp\[6\] d2.saw_temp\[5\] d2.saw_temp\[2\] d2.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and4_1
Xhold113 d8.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 d2.count\[7\] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 d11.count\[5\] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 d13.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 d2.count\[5\] vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ clknet_leaf_31_clk d13.nxt_count\[3\] net31 vssd1 vssd1 vccd1 vccd1 d13.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold168 d13.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 em0.u1.Q\[5\] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 d1.count\[5\] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlygate4sd3_1
X_4376_ clknet_leaf_0_clk d10.nxt_count\[3\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3327_ em0.u1.state\[2\] _0326_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__nand2_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _0804_ _0692_ _0822_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__or3_1
X_2209_ d4.count\[0\] d4.count\[1\] d4.count\[2\] vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__and3_1
X_3189_ d4.saw_temp\[2\] _0347_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ d12.count\[5\] d12.count\[4\] _0243_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__and3_1
X_2491_ _0192_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_4230_ clknet_leaf_28_clk d2.nxt_count\[5\] net28 vssd1 vssd1 vccd1 vccd1 d2.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4161_ _1710_ net102 net106 vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__a21oi_1
X_4092_ _1639_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__inv_2
X_3112_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__inv_2
X_3043_ _0300_ _0306_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_77_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3945_ _1503_ _1504_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ _1335_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2827_ _1847_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__inv_2
X_2758_ net145 _0409_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2689_ _0347_ _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__or2_1
X_4428_ clknet_leaf_20_clk _0097_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[9\] sky130_fd_sc_hd__dfrtp_1
X_4359_ clknet_leaf_37_clk d9.nxt_count\[8\] net22 vssd1 vssd1 vccd1 vccd1 d9.count\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout30 net34 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_6
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3730_ d1.saw_temp\[5\] _0330_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3661_ _0995_ _1108_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__o21ai_2
X_3592_ _1052_ _1060_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__a21o_1
X_2612_ _0286_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_2543_ d12.count\[8\] _1805_ _1720_ d12.count\[7\] _0234_ vssd1 vssd1 vccd1 vccd1
+ _0235_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2474_ _0179_ _0180_ _0172_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__and3b_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4213_ clknet_leaf_37_clk d1.nxt_count\[3\] net24 vssd1 vssd1 vccd1 vccd1 d1.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4144_ _1683_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ em0.u1.state\[2\] em0.u1.state\[1\] vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3026_ net135 _0598_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3928_ _1486_ _1487_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3859_ _0751_ _1419_ _0875_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2190_ d3.count\[8\] _1835_ d3.count\[9\] vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3713_ _0672_ _1274_ _0646_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3644_ _1089_ _1092_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3575_ d8.saw_temp\[7\] _1023_ _0702_ d8.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 _1138_
+ sky130_fd_sc_hd__o22a_1
X_2526_ _0220_ _0221_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
X_2457_ d10.count\[4\] _1733_ _0166_ _1735_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__o22a_1
Xhold17 d8.count\[0\] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold28 _0130_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _1996_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
Xhold39 p0.count\[0\] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_1
X_4127_ d12.saw_temp\[4\] d12.saw_temp\[3\] _1673_ vssd1 vssd1 vccd1 vccd1 _1675_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4058_ _1564_ _1574_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__and2_1
X_3009_ net142 _0585_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3360_ _0920_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__xor2_1
X_2311_ _1933_ _1934_ _1922_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__and3b_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _0620_ _0630_ _0852_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__or4_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ d5.count\[4\] _1718_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__xor2_1
X_2173_ d3.count\[3\] _1823_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3627_ net21 _1073_ _1074_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__o21a_1
X_3558_ _0723_ _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nor2_1
X_2509_ d11.count\[1\] d11.count\[0\] vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__or2_1
X_3489_ _1047_ _1051_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2860_ d5.saw_temp\[7\] _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2791_ _0431_ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ clknet_leaf_17_clk _0120_ net38 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3412_ d12.saw_temp\[2\] _0340_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__nand2_1
X_4392_ clknet_leaf_2_clk d11.nxt_count\[1\] net23 vssd1 vssd1 vccd1 vccd1 d11.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3343_ d3.saw_temp\[7\] _0796_ _0793_ d3.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0908_
+ sky130_fd_sc_hd__o22a_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ d9.saw_temp\[7\] _0335_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__or2b_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2225_ _1864_ _1865_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2156_ _1721_ d3.count\[3\] vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__nor2_1
X_2087_ _1757_ _1758_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ d1.saw_temp\[7\] _0572_ _0563_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3961_ _0723_ _0635_ _1413_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__or3_1
X_2912_ net189 _0514_ _0518_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3892_ d5.saw_temp\[6\] _0328_ _0739_ _0760_ _0310_ vssd1 vssd1 vccd1 vccd1 _1452_
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2843_ _0468_ _0469_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__nor2_1
X_2774_ _0416_ _0420_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold114 d9.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold103 d12.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 d12.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 d10.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 d3.count\[7\] vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ clknet_leaf_31_clk d13.nxt_count\[2\] net31 vssd1 vssd1 vccd1 vccd1 d13.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold136 em0.mixed_sample\[6\] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4375_ clknet_leaf_0_clk d10.nxt_count\[2\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold169 m0.edgy.delay vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _0780_ _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nor2_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _0804_ _0692_ _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__o21ai_2
X_2208_ _1853_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_3188_ d4.saw_temp\[3\] _0347_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__nand2_1
X_2139_ d2.count\[7\] d2.count\[6\] _1795_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2490_ _0172_ _0191_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4160_ em0.u1.state\[1\] em0.u1.count\[0\] em0.u1.count\[1\] vssd1 vssd1 vccd1 vccd1
+ _1687_ sky130_fd_sc_hd__and3_1
X_3111_ _0667_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__xor2_1
X_4091_ _1636_ _1637_ _1635_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__o21a_1
X_3042_ _0306_ _0300_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3944_ _1498_ _1502_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3875_ _1434_ _1435_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2826_ d4.saw_temp\[7\] _0456_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2757_ _0408_ _0409_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2688_ net8 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__buf_4
X_4427_ clknet_leaf_20_clk _0096_ net39 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[8\] sky130_fd_sc_hd__dfrtp_1
X_4358_ clknet_leaf_37_clk d9.nxt_count\[7\] net22 vssd1 vssd1 vccd1 vccd1 d9.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ clknet_leaf_31_clk _0032_ net31 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
X_3309_ _0301_ _0647_ _0307_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout31 net33 vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3660_ _1107_ _1106_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3591_ _1152_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__nand2_1
X_2611_ _0266_ _0285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2542_ d12.count\[7\] _1720_ _0230_ _0232_ _0233_ vssd1 vssd1 vccd1 vccd1 _0234_
+ sky130_fd_sc_hd__a221o_1
X_4212_ clknet_leaf_37_clk d1.nxt_count\[2\] net24 vssd1 vssd1 vccd1 vccd1 d1.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2473_ d10.count\[3\] _0176_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__or2_1
X_4143_ em0.mixed_sample\[4\] net251 em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1 _1683_
+ sky130_fd_sc_hd__mux2_1
X_4074_ _0326_ _1627_ _1628_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__a31o_1
X_3025_ _0597_ _0599_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3927_ _1471_ _1395_ _1485_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3858_ _1417_ _1418_ _0683_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__mux2_1
X_2809_ net160 _0446_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__xor2_1
X_3789_ _0738_ _1349_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3712_ _0674_ _0834_ d10.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3643_ _1177_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__xnor2_2
X_3574_ _1136_ _1037_ _1031_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2525_ net175 _0218_ _0208_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__o21ai_1
X_2456_ _1872_ d10.count\[2\] d10.count\[3\] vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__o21a_1
Xhold29 d1.count\[0\] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 d8.nxt_count\[0\] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ _1994_ _1995_ _1990_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__and3b_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4126_ net149 _1673_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__xor2_1
X_4057_ _1584_ _1553_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__or2b_1
X_3008_ _0585_ _0586_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2310_ d6.count\[4\] _1929_ d6.count\[5\] vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__a21o_1
X_3290_ _0853_ _0855_ _0306_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__o21a_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ d5.count\[5\] _1715_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__or2_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2172_ _1826_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3626_ _1182_ _1188_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__xnor2_4
X_3557_ d4.saw_temp\[7\] _0755_ _0759_ d4.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 _1120_
+ sky130_fd_sc_hd__o22a_1
X_2508_ net65 _0208_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
X_3488_ _1047_ _1051_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__or2_1
X_2439_ net205 _0150_ _2023_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__o21ai_1
X_4109_ _1660_ _1607_ _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2790_ d2.saw_temp\[5\] _0430_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4460_ clknet_leaf_18_clk _0119_ net38 vssd1 vssd1 vccd1 vccd1 em0.mixed_sample\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4391_ clknet_leaf_1_clk d11.nxt_count\[0\] net23 vssd1 vssd1 vccd1 vccd1 d11.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3411_ _0683_ _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3342_ d3.saw_temp\[2\] _0348_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ d9.saw_temp\[1\] _0335_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__nand2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ net212 _1862_ _1850_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__o21ai_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2155_ d3.count\[4\] _1714_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2086_ net230 _1755_ _1745_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2988_ _0562_ _0559_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3609_ _0683_ _1170_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3960_ _0635_ _1519_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2911_ _0514_ _0517_ d7.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3891_ _0739_ _1450_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2842_ net104 _0466_ net161 vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2773_ _1779_ _1773_ _0417_ _0419_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold104 d7.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _1704_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold126 d1.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _0584_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4443_ clknet_leaf_21_clk d13.nxt_count\[1\] net32 vssd1 vssd1 vccd1 vccd1 d13.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold159 d13.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 em0.mixed_sample\[7\] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dlygate4sd3_1
X_4374_ clknet_leaf_0_clk d10.nxt_count\[1\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _0803_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__xnor2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _0816_ _0821_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__xnor2_1
X_2207_ _1850_ _1851_ _1852_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__and3_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3187_ d4.saw_temp\[5\] d4.saw_temp\[4\] d4.saw_temp\[1\] _0347_ vssd1 vssd1 vccd1
+ vccd1 _0754_ sky130_fd_sc_hd__o31a_1
X_2138_ _1797_ _1798_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
X_2069_ net80 _1745_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_48_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3110_ _0669_ _0676_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ em0.u1.R\[18\] _1633_ _0893_ _1642_ _1646_ vssd1 vssd1 vccd1 vccd1 _0106_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3041_ _0608_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
X_3943_ _1498_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3874_ _1336_ _1337_ _1433_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__or3_1
X_2825_ d4.saw_temp\[6\] d4.saw_temp\[0\] d4.saw_temp\[3\] _0455_ vssd1 vssd1 vccd1
+ vccd1 _0456_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2756_ d13.saw_temp\[2\] d13.saw_temp\[1\] _0407_ vssd1 vssd1 vccd1 vccd1 _0409_
+ sky130_fd_sc_hd__and3_1
X_2687_ net9 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4426_ clknet_leaf_5_clk _0095_ net26 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4357_ clknet_leaf_37_clk d9.nxt_count\[6\] net22 vssd1 vssd1 vccd1 vccd1 d9.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ clknet_leaf_35_clk net50 net25 vssd1 vssd1 vccd1 vccd1 d5.count\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _0870_ _0873_ _0646_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__mux2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ d8.saw_temp\[1\] _0337_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout32 net33 vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_6
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3590_ _1146_ _1151_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__or2_1
X_2610_ d13.count\[8\] _0282_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2541_ _1727_ d12.count\[6\] vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2472_ d10.count\[3\] _0176_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__and2_1
X_4211_ clknet_leaf_37_clk d1.nxt_count\[1\] net24 vssd1 vssd1 vccd1 vccd1 d1.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_4142_ _1682_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
X_4073_ em0.u1.R\[16\] _1609_ _1630_ em0.u1.state\[1\] vssd1 vssd1 vccd1 vccd1 _1631_
+ sky130_fd_sc_hd__o211a_1
X_3024_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3926_ _1471_ _1395_ _1485_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_18_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3857_ d12.saw_temp\[6\] _0340_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__nand2_1
X_2808_ _0435_ _0441_ _0446_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a21oi_1
X_3788_ d3.saw_temp\[7\] _0771_ _0793_ d3.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 _1349_
+ sky130_fd_sc_hd__o22a_1
X_2739_ _0327_ em0.u1.D\[12\] vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__and2_1
X_4409_ clknet_leaf_38_clk d12.nxt_count\[0\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3711_ _0749_ _1272_ _0659_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3642_ _1202_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__xnor2_2
X_3573_ _1033_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2524_ d11.count\[5\] d11.count\[4\] _0215_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__and3_1
X_2455_ _1723_ _0164_ d10.count\[5\] vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__a21bo_1
X_2386_ d8.count\[1\] d8.count\[0\] d8.count\[2\] vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__a21o_1
Xhold19 d6.count\[0\] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlygate4sd3_1
X_4125_ _1673_ _1674_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__nor2_1
X_4056_ _1581_ _1583_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__or2_1
X_3007_ net120 _0583_ net144 vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3909_ _1449_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ d5.count\[5\] _1715_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2171_ _1819_ _1824_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3625_ _1186_ _1187_ _1064_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3556_ _1117_ _1118_ _0747_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2507_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_2
X_3487_ _0749_ _1050_ _0669_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2438_ d9.count\[5\] d9.count\[4\] _0147_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__and3_1
X_2369_ d8.count\[4\] _1726_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__nor2_1
X_4108_ em0.u1.R\[21\] _1606_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__nand2_1
X_4039_ _1596_ _1597_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4390_ clknet_leaf_5_clk _0079_ net27 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3410_ d12.saw_temp\[7\] _0870_ _0871_ d12.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1
+ _0975_ sky130_fd_sc_hd__o22a_1
X_3341_ _0904_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _0832_ _0837_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__xor2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ d4.count\[6\] _1862_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__and2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ d3.count\[2\] _1733_ _1810_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__a21oi_1
X_2085_ d1.count\[5\] d1.count\[4\] _1753_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2987_ net108 _0569_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3608_ d9.saw_temp\[4\] _0335_ _0682_ _0309_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3539_ _0986_ _0987_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2910_ d7.saw_temp\[7\] _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3890_ _0743_ _1340_ _0738_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__a21oi_1
X_2841_ d4.saw_temp\[4\] d4.saw_temp\[3\] _0466_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__and3_1
X_2772_ _1712_ d2.count\[2\] _1782_ _0418_ d2.count\[0\] vssd1 vssd1 vccd1 vccd1 _0419_
+ sky130_fd_sc_hd__a2111o_1
Xhold105 d9.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 d8.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ clknet_leaf_21_clk net72 net32 vssd1 vssd1 vccd1 vccd1 d13.count\[0\] sky130_fd_sc_hd__dfrtp_2
Xhold138 d7.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 d2.count\[4\] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 d1.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dlygate4sd3_1
X_4373_ clknet_leaf_0_clk d10.nxt_count\[0\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _0888_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__nand2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _0750_ _0820_ _0722_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__a21o_1
X_2206_ d4.count\[0\] d4.count\[1\] vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__or2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ d4.saw_temp\[7\] _0347_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2137_ d2.count\[6\] _1795_ _1783_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__o21ai_1
X_2068_ _1719_ _1743_ _1744_ _1724_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_76_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3040_ _0595_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3942_ _1500_ _1501_ _0681_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3873_ _1336_ _1337_ _1433_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2824_ d4.saw_temp\[5\] d4.saw_temp\[4\] d4.saw_temp\[1\] d4.saw_temp\[2\] vssd1
+ vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2755_ d13.saw_temp\[1\] _0407_ net219 vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__a21oi_1
X_2686_ net11 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__clkbuf_4
X_4425_ clknet_leaf_10_clk _0094_ net37 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4356_ clknet_leaf_38_clk d9.nxt_count\[5\] net22 vssd1 vssd1 vccd1 vccd1 d9.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3307_ _0871_ _0872_ d12.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__mux2_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ clknet_leaf_30_clk d5.nxt_count\[8\] net29 vssd1 vssd1 vccd1 vccd1 d5.count\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3238_ _0667_ _0677_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__nor2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__inv_2
Xfanout22 net34 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_6
XFILLER_0_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout33 net34 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_4
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2540_ _1872_ d12.count\[5\] d12.count\[4\] _1723_ _0231_ vssd1 vssd1 vccd1 vccd1
+ _0232_ sky130_fd_sc_hd__a221o_1
X_2471_ _0178_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4210_ clknet_leaf_37_clk d1.nxt_count\[0\] net24 vssd1 vssd1 vccd1 vccd1 d1.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4141_ em0.mixed_sample\[3\] em0.u1.Q\[3\] em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _1682_ sky130_fd_sc_hd__mux2_1
X_4072_ _1609_ _1629_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__nand2_1
X_3023_ d11.saw_temp\[0\] _0596_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__nand2_1
X_3925_ _1480_ _1484_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3856_ d12.saw_temp\[7\] _0650_ _0871_ d12.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1
+ _1417_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2807_ d3.saw_temp\[0\] _0445_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__and2_1
X_3787_ _1343_ _1347_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2738_ em0.u1.state\[2\] net158 _0393_ _0394_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__o22a_1
X_4408_ clknet_leaf_10_clk _0087_ net37 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_2669_ net7 vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4339_ clknet_leaf_36_clk d8.nxt_count\[6\] net24 vssd1 vssd1 vccd1 vccd1 d8.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4418__43 vssd1 vssd1 vccd1 vccd1 _4418__43/HI net43 sky130_fd_sc_hd__conb_1
XFILLER_0_37_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3710_ _0662_ _1271_ _0646_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3641_ _1084_ _1088_ _1203_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__a21boi_2
X_3572_ _1114_ _1134_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2523_ _0218_ _0219_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
X_2454_ d10.count\[4\] _1733_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__nand2_1
X_2385_ d8.count\[1\] d8.count\[0\] d8.count\[2\] vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__and3_1
X_4124_ d12.saw_temp\[1\] _1672_ net211 vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__a21oi_1
Xinput1 modes vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_4055_ _1585_ _1587_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__or2_1
X_3006_ d10.saw_temp\[4\] d10.saw_temp\[3\] _0583_ vssd1 vssd1 vccd1 vccd1 _0585_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3908_ _1466_ _1467_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__nor2_1
X_3839_ _1398_ _1399_ _0640_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ d3.count\[0\] d3.count\[1\] d3.count\[2\] vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3624_ d1.saw_temp\[4\] _0330_ _0640_ _0309_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3555_ d5.saw_temp\[4\] _0328_ _0683_ _0310_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a31o_1
X_3486_ _1048_ _1049_ _0634_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__mux2_1
X_2506_ _0205_ _0206_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__and2_1
X_2437_ _0150_ _0151_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2368_ _1979_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_4107_ em0.u1.R\[22\] vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__inv_2
X_2299_ d6.count\[1\] d6.count\[0\] d6.count\[2\] vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__nand3_1
X_4038_ em0.u1.R\[16\] em0.u1.D\[9\] vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3340_ _0900_ _0903_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__or2_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _0622_ _0836_ _0669_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__a21o_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _1862_ _1863_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _1721_ d3.count\[3\] vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ _1755_ _1756_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_0_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2986_ _0571_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_1
X_3607_ d9.saw_temp\[7\] _1055_ _0688_ d9.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 _1170_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ _1018_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__xor2_1
X_3469_ _1031_ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2840_ net104 _0466_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2771_ d2.count\[8\] _1717_ _1768_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4441_ clknet_leaf_16_clk _0110_ net16 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[22\] sky130_fd_sc_hd__dfrtp_1
Xhold106 d4.count\[4\] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 d6.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 em0.mixed_sample\[1\] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 em0.mixed_sample\[0\] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ clknet_leaf_17_clk _0000_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _0886_ _0887_ _0735_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__o21ai_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _0817_ _0819_ _0646_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__mux2_1
X_2205_ d4.count\[0\] d4.count\[1\] vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ d4.saw_temp\[0\] _0347_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__nand2_1
X_2136_ d2.count\[6\] _1795_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2067_ d1.count\[9\] vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2969_ d1.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3941_ _0738_ _0680_ _1392_ _0751_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3872_ _1357_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2823_ _0444_ _0454_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__nor2_1
X_2754_ net153 _0407_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2685_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
X_4424_ clknet_leaf_9_clk _0093_ net36 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4355_ clknet_leaf_38_clk d9.nxt_count\[4\] net22 vssd1 vssd1 vccd1 vccd1 d9.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3306_ d12.saw_temp\[7\] _0340_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__or2b_1
X_4286_ clknet_leaf_27_clk d5.nxt_count\[7\] net29 vssd1 vssd1 vccd1 vccd1 d5.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _0801_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__nand2_1
X_3168_ _0695_ _0696_ _0734_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__or3_2
X_2119_ d2.count\[1\] d2.count\[0\] vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__or2_1
X_3099_ _0640_ _0664_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout23 net34 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_8
Xfanout34 net16 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2470_ _0176_ _0177_ _0172_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4140_ _1681_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
X_4071_ _1598_ _1599_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__xnor2_1
X_3022_ net247 _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3924_ _0722_ _1483_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3855_ _1411_ _1415_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__xor2_2
X_2806_ _0444_ _0441_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__or2b_1
X_3786_ _1345_ _1346_ _0762_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__o21a_1
X_2737_ _0372_ _0377_ _0380_ _0389_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2668_ net10 vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__buf_4
X_4407_ clknet_leaf_13_clk _0086_ net40 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2599_ _0276_ _0277_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
X_4338_ clknet_leaf_36_clk d8.nxt_count\[5\] net24 vssd1 vssd1 vccd1 vccd1 d8.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4269_ clknet_leaf_28_clk d4.nxt_count\[8\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3640_ _1078_ _1083_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3571_ _1132_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__nor2_1
X_2522_ net234 _0215_ _0208_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2453_ d10.count\[6\] vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__inv_2
X_4360__46 vssd1 vssd1 vccd1 vccd1 _4360__46/HI net46 sky130_fd_sc_hd__conb_1
X_2384_ _1993_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_4123_ d12.saw_temp\[2\] d12.saw_temp\[1\] _1672_ vssd1 vssd1 vccd1 vccd1 _1673_
+ sky130_fd_sc_hd__and3_1
X_4054_ _1589_ _1591_ _1612_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__a21o_1
Xinput2 octaves vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_3005_ net120 _0583_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3907_ _1377_ _1379_ _1465_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3838_ d2.saw_temp\[6\] _0329_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3769_ _1327_ _1328_ _1330_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__o21ai_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3623_ _0640_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3554_ _0723_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__nor2_1
X_3485_ d10.saw_temp\[7\] _0946_ _0674_ d10.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1
+ _1049_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2505_ d11.count\[8\] _1715_ d11.count\[9\] vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a21oi_1
X_2436_ d9.count\[4\] _0147_ _2023_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__o21ai_1
X_2367_ _1959_ _1978_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4106_ _1710_ _1609_ _1659_ net67 _0782_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__a32o_1
X_2298_ _1925_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4037_ em0.u1.D\[9\] em0.u1.R\[16\] vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap20 net21 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3270_ _0833_ _0835_ _0634_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__mux2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ net141 _1860_ _1850_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__o21ai_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ d3.count\[2\] _1733_ _1808_ _1721_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__a2bb2o_1
X_2083_ net250 _1753_ _1745_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2985_ _0569_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3606_ _1167_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3537_ _1098_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3468_ _1026_ _1030_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2419_ d9.count\[7\] _1720_ _2011_ _2020_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__a22o_1
X_3399_ d1.saw_temp\[1\] _0623_ _0627_ _0963_ _0618_ vssd1 vssd1 vccd1 vccd1 _0964_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2770_ d2.count\[1\] d2.count\[6\] _1732_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4440_ clknet_leaf_16_clk _0109_ net16 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[21\] sky130_fd_sc_hd__dfrtp_1
Xhold107 em0.u1.D\[11\] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 d7.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 d1.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dlygate4sd3_1
X_4371_ clknet_leaf_17_clk _0002_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _0735_ _0886_ _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__or3_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _0728_ _0818_ d6.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__mux2_1
X_3184_ _0750_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__buf_6
X_2204_ net74 _1850_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _1795_ _1796_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
X_2066_ d1.count\[8\] _1720_ _1723_ d1.count\[7\] _1742_ vssd1 vssd1 vccd1 vccd1 _1743_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2968_ _1737_ _0552_ _0554_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__or4_2
XFILLER_0_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2899_ net112 _0507_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3940_ _0680_ _1499_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3871_ _1429_ _1431_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__xnor2_1
X_2822_ _0453_ _0441_ d3.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2753_ net191 _0403_ _0407_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2684_ net6 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__clkbuf_4
X_4423_ clknet_leaf_9_clk _0092_ net37 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
X_4354_ clknet_leaf_36_clk d9.nxt_count\[3\] net24 vssd1 vssd1 vccd1 vccd1 d9.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _0647_ _0651_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand2_2
X_4285_ clknet_leaf_27_clk d5.nxt_count\[6\] net28 vssd1 vssd1 vccd1 vccd1 d5.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _0764_ _0775_ _0800_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__or3_1
X_3167_ _0732_ _0733_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__or2_1
X_3098_ d11.saw_temp\[0\] _0334_ _0640_ _0309_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__a31o_1
X_2118_ d2.count\[1\] d2.count\[0\] vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__nand2_1
X_2049_ _1724_ _1725_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__nor2_4
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout24 net34 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_6
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout35 net37 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_6
XFILLER_0_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _1613_ _1589_ _1626_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__nand3_1
X_3021_ _0198_ _0589_ _0592_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__a31o_2
XFILLER_0_46_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3923_ _0738_ _0721_ _1371_ _1482_ _0751_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__o311a_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3854_ _0750_ _1414_ _0866_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2805_ d3.saw_temp\[7\] _0442_ _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__and3_1
X_3785_ d4.saw_temp\[6\] _0347_ _0738_ _0310_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__a31o_1
X_2736_ em0.u1.state\[2\] _0391_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__nand2_1
X_2667_ em0.u1.state\[2\] vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__inv_2
X_4406_ clknet_leaf_11_clk _0085_ net40 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2598_ net215 _0273_ _0266_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ clknet_leaf_36_clk d8.nxt_count\[4\] net24 vssd1 vssd1 vccd1 vccd1 d8.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4268_ clknet_leaf_29_clk d4.nxt_count\[7\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3219_ _0744_ _0784_ d5.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__mux2_1
X_4199_ clknet_leaf_24_clk p0.nxt_count\[7\] net32 vssd1 vssd1 vccd1 vccd1 p0.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _1039_ _1115_ _1131_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2521_ d11.count\[3\] d11.count\[4\] _0212_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2452_ _1727_ d10.count\[6\] vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2383_ _1990_ _1991_ _1992_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__and3_1
X_4122_ net154 _1672_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__xor2_1
X_4053_ _1610_ _1611_ em0.u1.R\[16\] _0782_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__a2bb2o_1
X_3004_ _0583_ net199 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__nor2_1
Xinput3 pb[0] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
X_3906_ _1377_ _1379_ _1465_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3837_ d2.saw_temp\[5\] _0611_ _0615_ _1287_ d2.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1
+ _1398_ sky130_fd_sc_hd__o32a_1
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3768_ _1222_ _1224_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2719_ _0339_ _0342_ _0376_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__and3_1
X_3699_ _0726_ _1260_ _0646_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__mux2_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4342__47 vssd1 vssd1 vccd1 vccd1 _4342__47/HI net47 sky130_fd_sc_hd__conb_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3622_ d1.saw_temp\[3\] _0623_ _0627_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3553_ d5.saw_temp\[7\] _1000_ _0744_ d5.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 _1116_
+ sky130_fd_sc_hd__o22a_1
X_3484_ d10.saw_temp\[3\] _0336_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__nand2_1
X_2504_ d11.count\[8\] _1805_ _0204_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__o21ai_1
X_2435_ d9.count\[3\] d9.count\[4\] _2027_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__and3_1
X_4105_ _1606_ _1658_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__nand2_1
X_2366_ d7.count\[8\] _1975_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__xnor2_1
X_2297_ _1922_ _1923_ _1924_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__and3_1
X_4036_ em0.u1.D\[10\] vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ d4.count\[4\] d4.count\[5\] _1857_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__and3_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2151_ _1713_ d3.count\[0\] d3.count\[1\] vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__o21ai_1
X_2082_ d1.count\[3\] d1.count\[4\] _1749_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2984_ d1.saw_temp\[5\] _0567_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3605_ _1162_ _1166_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3536_ _0941_ _0985_ _1099_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__a21o_1
X_3467_ _1026_ _1030_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__nor2_1
X_2418_ _1727_ d9.count\[6\] _2018_ _2019_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__a211o_1
X_3398_ _0560_ d1.saw_temp\[1\] _0330_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__nand3_1
X_2349_ d7.count\[3\] _1963_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__and2_1
X_4019_ _1575_ _1577_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 d11.count\[6\] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 d2.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ clknet_leaf_17_clk _0001_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3321_ _0884_ _0885_ _0827_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__o21a_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ d6.saw_temp\[7\] _0346_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__or2b_1
X_2203_ d4.count\[8\] _1805_ _1849_ d4.count\[9\] vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__a211oi_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _0749_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__buf_6
X_2134_ net197 _1793_ _1783_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2065_ d1.count\[7\] _1723_ _1726_ d1.count\[6\] _1741_ vssd1 vssd1 vccd1 vccd1 _1742_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2967_ _1945_ _1730_ _0555_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2898_ d6.saw_temp\[5\] _0505_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__and2_1
X_3519_ _0310_ _1080_ _1082_ _0633_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__o31a_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3870_ _1270_ _1316_ _1430_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2821_ _0442_ _0443_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2752_ _0406_ _0403_ d13.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__o21a_1
X_4422_ clknet_leaf_9_clk _0091_ net36 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_2
X_2683_ _0341_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__nand2_1
X_4353_ clknet_leaf_36_clk d9.nxt_count\[2\] net24 vssd1 vssd1 vccd1 vccd1 d9.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4284_ clknet_leaf_29_clk d5.nxt_count\[5\] net28 vssd1 vssd1 vccd1 vccd1 d5.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ d12.saw_temp\[1\] _0340_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nand2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _0764_ _0775_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__o21ai_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _0720_ _0731_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__and2_1
X_3097_ _0658_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__nand2_2
X_2117_ net111 _1783_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2048_ _1712_ _1713_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__nor2_4
Xfanout36 net37 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_6
Xfanout25 net34 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3999_ _1556_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3020_ d11.saw_temp\[7\] _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__and2_1
X_3922_ _0721_ _1481_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3853_ _1412_ _1413_ _0683_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2804_ d3.saw_temp\[6\] d3.saw_temp\[5\] d3.saw_temp\[2\] d3.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3784_ _0738_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__nor2_1
X_2735_ _0327_ net244 _0391_ _0392_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a22o_1
X_2666_ _0326_ _1711_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__nor2_1
X_4405_ clknet_leaf_11_clk _0084_ net37 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_4336_ clknet_leaf_36_clk d8.nxt_count\[3\] net24 vssd1 vssd1 vccd1 vccd1 d8.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2597_ d13.count\[3\] d13.count\[4\] _0270_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__and3_1
X_4267_ clknet_leaf_29_clk d4.nxt_count\[6\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4198_ clknet_leaf_24_clk p0.nxt_count\[6\] net32 vssd1 vssd1 vccd1 vccd1 p0.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3218_ d5.saw_temp\[7\] _0328_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__or2b_1
X_3149_ _0708_ _0715_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2520_ _0217_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2451_ d10.count\[8\] _1715_ _1718_ d10.count\[7\] vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__o22a_1
X_2382_ d8.count\[1\] d8.count\[0\] vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__nand2_1
X_4121_ net201 _1668_ _1672_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__o21ba_1
X_4052_ em0.u1.D\[8\] em0.u1.R\[15\] _1609_ _0326_ vssd1 vssd1 vccd1 vccd1 _1611_
+ sky130_fd_sc_hd__a31o_1
Xinput4 pb[10] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_3003_ d10.saw_temp\[1\] _0581_ net198 vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3905_ _1463_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__or2_1
X_3836_ _1395_ _1396_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__or2b_2
XFILLER_0_6_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3767_ _1218_ _1221_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2718_ _0339_ _0342_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3698_ _0728_ _0818_ d6.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__mux2_1
X_2649_ p0.count\[7\] vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4319_ clknet_leaf_35_clk d7.nxt_count\[4\] net25 vssd1 vssd1 vccd1 vccd1 d7.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3621_ d1.saw_temp\[3\] _1183_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3552_ _1019_ _1040_ _1041_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2503_ d11.count\[7\] _1720_ _0193_ _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__a22o_1
X_3483_ _0749_ _1046_ _0659_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__a21o_1
X_2434_ _0149_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_2365_ _1977_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_4104_ _1657_ _1605_ em0.u1.R\[20\] vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__a21bo_1
X_2296_ d6.count\[1\] d6.count\[0\] vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__nand2_1
X_4035_ em0.u1.D\[11\] vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__inv_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3819_ _1377_ _1378_ _1257_ _1358_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4324__48 vssd1 vssd1 vccd1 vccd1 _4324__48/HI net48 sky130_fd_sc_hd__conb_1
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2150_ d3.count\[7\] _1723_ _1732_ d3.count\[6\] vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2081_ _1753_ _1754_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_88_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2983_ d1.saw_temp\[5\] _0567_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3604_ _1162_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3535_ _0984_ _0983_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__and2b_1
X_3466_ _0622_ _1029_ _0708_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a21o_1
X_2417_ _1872_ d9.count\[4\] d9.count\[5\] _1721_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3397_ d1.saw_temp\[2\] _0330_ _0301_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2348_ _1965_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_2279_ _1908_ vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4018_ _1489_ _1535_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_79_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold109 d3.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3320_ _0827_ _0884_ _0885_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__nor3_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ d6.saw_temp\[1\] _0346_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__nand2_1
X_2202_ d4.count\[8\] _1805_ _1847_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__o22a_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _0622_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__clkbuf_8
X_2133_ d2.count\[5\] d2.count\[4\] _1791_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__and3_1
X_2064_ d1.count\[5\] _1720_ _1728_ _1739_ _1740_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2966_ d1.count\[8\] _1720_ _1723_ d1.count\[7\] _0556_ vssd1 vssd1 vccd1 vccd1 _0557_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2897_ net140 _0505_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3518_ _0646_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__nor2_1
X_3449_ _0751_ _1012_ _0767_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__a21boi_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2820_ net114 _0452_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2751_ d13.saw_temp\[7\] _0405_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2682_ _0340_ _0338_ _0339_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__nand3_1
X_4421_ clknet_leaf_9_clk _0090_ net36 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
X_4352_ clknet_leaf_36_clk d9.nxt_count\[1\] net24 vssd1 vssd1 vccd1 vccd1 d9.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_4283_ clknet_leaf_29_clk d5.nxt_count\[4\] net29 vssd1 vssd1 vccd1 vccd1 d5.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _0859_ _0860_ _0867_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__a21o_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _0792_ _0799_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__xnor2_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3165_ _0720_ _0731_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__nor2_1
X_3096_ d11.saw_temp\[6\] _0660_ _0661_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__or4b_1
X_2116_ _1767_ _1781_ _1782_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2047_ _1721_ _1716_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__nor2_8
XFILLER_0_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout26 net27 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_6
Xfanout37 net16 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
XFILLER_0_76_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ _1486_ _1554_ _1555_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__nand3_1
X_2949_ net164 _0543_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3921_ _0727_ _1371_ _0723_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3852_ d13.saw_temp\[6\] _0344_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2803_ d3.saw_temp\[4\] d3.saw_temp\[3\] d3.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1
+ _0442_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3783_ _0759_ _1235_ d4.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2734_ _0383_ _0387_ _0390_ em0.u1.state\[2\] vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__o31a_1
X_2665_ em0.u1.state\[1\] vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4404_ clknet_leaf_11_clk _0083_ net37 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2596_ _0275_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4335_ clknet_leaf_36_clk d8.nxt_count\[2\] net24 vssd1 vssd1 vccd1 vccd1 d8.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4266_ clknet_leaf_29_clk d4.nxt_count\[5\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4197_ clknet_leaf_22_clk p0.nxt_count\[5\] net32 vssd1 vssd1 vccd1 vccd1 p0.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3217_ d5.saw_temp\[1\] _0328_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3148_ _0682_ _0713_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3079_ _0634_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__buf_8
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2450_ _0160_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_2381_ d8.count\[1\] d8.count\[0\] vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__or2_1
X_4120_ _1671_ _1668_ d12.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__o21a_1
X_4051_ em0.u1.D\[8\] _1609_ em0.u1.R\[15\] vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__a21oi_1
X_3002_ d10.saw_temp\[2\] d10.saw_temp\[1\] _0581_ vssd1 vssd1 vccd1 vccd1 _0583_
+ sky130_fd_sc_hd__and3_1
Xinput5 pb[11] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3904_ _1458_ _1462_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3835_ _1390_ _1394_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3766_ _1215_ _1228_ _1326_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2717_ _0374_ _0375_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__xnor2_1
X_3697_ _1257_ _1258_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2648_ _0307_ _0303_ _0310_ _0302_ vssd1 vssd1 vccd1 vccd1 s0.next_q\[1\] sky130_fd_sc_hd__a22o_1
XFILLER_0_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2579_ d13.count\[4\] _1720_ _0261_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__o21a_1
X_4318_ clknet_leaf_33_clk d7.nxt_count\[3\] net34 vssd1 vssd1 vccd1 vccd1 d7.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4249_ clknet_leaf_24_clk d3.nxt_count\[6\] net32 vssd1 vssd1 vccd1 vccd1 d3.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3620_ d1.saw_temp\[7\] _0330_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__and2b_1
X_3551_ _1008_ _1013_ _1007_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2502_ _0194_ _0200_ _0201_ _0202_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3482_ _1044_ _1045_ _0634_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2433_ _0147_ _0148_ _2023_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__and3b_1
X_2364_ _1959_ _1975_ _1976_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__and3_1
X_4103_ em0.u1.D\[12\] em0.u1.R\[19\] vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__or2b_1
X_2295_ d6.count\[1\] d6.count\[0\] vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__or2_1
X_4034_ em0.u1.R\[19\] em0.u1.D\[12\] vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3818_ _1257_ _1358_ _1377_ _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3749_ _0633_ _1192_ _1195_ _1197_ _1201_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_30_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ net213 _1749_ _1745_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2982_ _0567_ _0568_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3603_ _0622_ _1164_ _1165_ _0669_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3534_ _1043_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__xnor2_1
X_3465_ _1027_ _1028_ _0634_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__mux2_1
X_2416_ d9.count\[2\] _1724_ _2015_ _2017_ d9.count\[3\] vssd1 vssd1 vccd1 vccd1 _2018_
+ sky130_fd_sc_hd__o2111a_1
X_4306__49 vssd1 vssd1 vccd1 vccd1 _4306__49/HI net49 sky130_fd_sc_hd__conb_1
X_3396_ _0307_ _0960_ _0620_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__a21o_1
X_2347_ _1963_ _1964_ _1959_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2278_ _1888_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4017_ _1534_ _1532_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _0810_ _0815_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__xor2_2
X_2201_ _1721_ d4.count\[7\] d4.count\[6\] _1725_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__a22o_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _0745_ _0746_ _0747_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__o21ai_1
X_2132_ _1793_ _1794_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_0_28_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2063_ d1.count\[6\] _1726_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2965_ d1.count\[6\] _1726_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2896_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3517_ d13.saw_temp\[3\] _0344_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__nand2_1
X_3448_ _1010_ _1011_ _0760_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__mux2_1
X_3379_ _0942_ _0943_ _0618_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__mux2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4369__41 vssd1 vssd1 vccd1 vccd1 _4369__41/HI net41 sky130_fd_sc_hd__conb_1
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2750_ d13.saw_temp\[4\] d13.saw_temp\[3\] d13.saw_temp\[0\] _0404_ vssd1 vssd1 vccd1
+ vccd1 _0405_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2681_ _0338_ _0339_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__a21o_1
X_4420_ clknet_leaf_9_clk _0089_ net36 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4351_ clknet_leaf_36_clk net77 net24 vssd1 vssd1 vccd1 vccd1 d9.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_4282_ clknet_leaf_35_clk d5.nxt_count\[3\] net29 vssd1 vssd1 vccd1 vccd1 d5.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _0859_ _0860_ _0867_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__nand3_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _0767_ _0798_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nand2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _0722_ _0730_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__or2_1
X_3095_ d11.saw_temp\[5\] _0334_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__nand2_1
X_2115_ d2.count\[9\] _1714_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__nor2_1
X_2046_ _1722_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__buf_6
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout27 net34 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_6
Xfanout38 net39 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_6
XFILLER_0_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3997_ _1486_ _1554_ _1555_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2948_ _0543_ net217 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2879_ _0483_ _0494_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__and2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _1475_ _1479_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3851_ d13.saw_temp\[7\] _0638_ _0862_ d13.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1
+ _1412_ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2802_ _1806_ _0436_ _0437_ _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or4_2
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3782_ _0747_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nand2_1
X_2733_ _0383_ _0387_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2664_ _0311_ net113 _0325_ vssd1 vssd1 vccd1 vccd1 p0.pwm sky130_fd_sc_hd__o21a_1
XFILLER_0_41_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4403_ clknet_leaf_10_clk _0082_ net37 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_2595_ _0273_ _0274_ _0266_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__and3b_1
X_4334_ clknet_leaf_36_clk d8.nxt_count\[1\] net24 vssd1 vssd1 vccd1 vccd1 d8.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4265_ clknet_leaf_29_clk d4.nxt_count\[4\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4196_ clknet_leaf_22_clk net226 net32 vssd1 vssd1 vccd1 vccd1 p0.count\[4\] sky130_fd_sc_hd__dfrtp_1
X_3216_ _0778_ _0779_ _0780_ _0782_ net66 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__a32o_1
X_3147_ d7.saw_temp\[0\] net12 _0640_ _0309_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ d12.saw_temp\[7\] _0301_ _0340_ _0307_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a31o_2
XFILLER_0_77_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2380_ net68 _1990_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
X_4050_ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__clkbuf_4
Xinput6 pb[12] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
X_3001_ net124 _0581_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3903_ _1458_ _1462_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__and2_1
X_3834_ _1390_ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3765_ _1215_ _1228_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__and3_1
X_3696_ _1253_ _1256_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__and2_1
X_2716_ _0345_ _0352_ _0355_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2647_ _0309_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_8
X_2578_ _0258_ _0259_ _0260_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4317_ clknet_leaf_33_clk d7.nxt_count\[2\] net27 vssd1 vssd1 vccd1 vccd1 d7.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4248_ clknet_leaf_24_clk d3.nxt_count\[5\] net30 vssd1 vssd1 vccd1 vccd1 d3.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4179_ d9.saw_temp\[1\] _1699_ net156 vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3550_ _1018_ _1101_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nor2_1
X_2501_ _1872_ d11.count\[4\] d11.count\[5\] vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__o21a_1
X_3481_ d11.saw_temp\[7\] _0942_ _0664_ d11.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1
+ _1045_ sky130_fd_sc_hd__o22a_1
X_2432_ d9.count\[3\] _2027_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__or2_1
X_2363_ d7.count\[7\] _1973_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__or2_1
X_4102_ net91 _0782_ _1656_ _1710_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__a22o_1
X_4033_ em0.u1.D\[12\] em0.u1.R\[19\] vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__and2b_1
X_2294_ net70 _1922_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3817_ _1277_ _1284_ _1376_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__nand3_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3748_ _1306_ _1309_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3679_ _1234_ _1239_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2981_ d1.saw_temp\[3\] _0565_ net172 vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3602_ d10.saw_temp\[4\] _0336_ _0682_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nand3_1
XFILLER_0_71_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3533_ _1094_ _1096_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__xnor2_2
X_3464_ d7.saw_temp\[7\] _0921_ _0713_ d7.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _1028_
+ sky130_fd_sc_hd__o22a_1
X_2415_ _1721_ _2016_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__nand2_1
X_3395_ _0618_ _0957_ _0958_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__a31o_1
X_2346_ d7.count\[0\] d7.count\[1\] d7.count\[2\] vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__a21o_1
X_2277_ d5.count\[8\] _1904_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__xnor2_1
X_4016_ _1564_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_32_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _1841_ _1842_ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__and3_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3180_ d5.saw_temp\[7\] _0301_ _0328_ _0307_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__a31o_2
X_2131_ net200 _1791_ _1783_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__o21ai_1
X_2062_ _1730_ _1737_ _1738_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2964_ d1.count\[6\] _1726_ _1728_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2895_ d6.saw_temp\[3\] _0503_ net168 vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__a21oi_1
X_3516_ _0682_ _1079_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3447_ d3.saw_temp\[7\] _0907_ _0793_ d3.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _1011_
+ sky130_fd_sc_hd__o22a_1
X_3378_ d11.saw_temp\[7\] _0828_ _0664_ d11.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1
+ _0943_ sky130_fd_sc_hd__o22a_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ d7.count\[1\] _1723_ _1777_ d7.count\[0\] vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2680_ net5 vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ clknet_leaf_13_clk _0063_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
X_3301_ _0622_ _0865_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__a21oi_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ clknet_leaf_30_clk d5.nxt_count\[2\] net29 vssd1 vssd1 vccd1 vccd1 d5.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3232_ _0738_ _0795_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__o21ai_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _0723_ _0728_ _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__o21ba_1
X_2114_ _1768_ _1780_ d2.count\[8\] _1720_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3094_ d11.saw_temp\[3\] d11.saw_temp\[0\] _0334_ vssd1 vssd1 vccd1 vccd1 _0661_
+ sky130_fd_sc_hd__o21a_1
X_2045_ _1721_ _1713_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout28 net30 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_6
XFILLER_0_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout39 net16 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_6
X_3996_ _1453_ _1457_ _1463_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2947_ d8.saw_temp\[1\] _0541_ net216 vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2878_ _0482_ _0479_ d5.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4479_ clknet_leaf_8_clk _0138_ net36 vssd1 vssd1 vccd1 vccd1 d9.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3850_ _1408_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__xnor2_2
X_2801_ _1809_ _1817_ _0438_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or4b_1
X_3781_ _0738_ _1339_ _1341_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2732_ _0380_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__xor2_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2663_ _0311_ em0.mixed_sample\[7\] _0313_ _0324_ vssd1 vssd1 vccd1 vccd1 _0325_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4402_ clknet_leaf_10_clk _0081_ net37 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2594_ d13.count\[3\] _0270_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4333_ clknet_leaf_36_clk net69 net24 vssd1 vssd1 vccd1 vccd1 d8.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_4264_ clknet_leaf_29_clk d4.nxt_count\[3\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3215_ _0781_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4195_ clknet_leaf_19_clk p0.nxt_count\[3\] net39 vssd1 vssd1 vccd1 vccd1 p0.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3146_ _0707_ _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__nand2_2
X_3077_ _0632_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3979_ _1536_ _1538_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3000_ _0581_ _0582_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__nor2_1
Xinput7 pb[1] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3902_ _0310_ _1460_ _1461_ _0767_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__o31a_1
XFILLER_0_86_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3833_ _0751_ _1393_ _0681_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3764_ _1229_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__xnor2_1
X_3695_ _1253_ _1256_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2715_ _0372_ _0373_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__or2_1
X_2646_ _0308_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2577_ _1727_ d13.count\[2\] d13.count\[3\] vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4316_ clknet_leaf_33_clk d7.nxt_count\[1\] net27 vssd1 vssd1 vccd1 vccd1 d7.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_4247_ clknet_leaf_24_clk d3.nxt_count\[4\] net30 vssd1 vssd1 vccd1 vccd1 d3.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4178_ d9.saw_temp\[1\] d9.saw_temp\[2\] _1699_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__and3_1
X_3129_ _0657_ _0694_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__and2_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3480_ d11.saw_temp\[3\] _0334_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2500_ _1727_ d11.count\[6\] vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2431_ d9.count\[3\] _2027_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__and2_1
X_2362_ d7.count\[7\] _1973_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__nand2_1
X_4101_ em0.u1.R\[19\] _1655_ _1609_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__mux2_1
X_2293_ _1920_ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__and2_2
X_4032_ _1588_ _1590_ _0893_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3816_ _1277_ _1284_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3747_ _0751_ _1308_ _0875_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3678_ _1234_ _1239_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2629_ _0296_ vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2980_ d1.saw_temp\[4\] d1.saw_temp\[3\] _0565_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3601_ _0640_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 pb[4] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3532_ _0955_ _0982_ _1095_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__a21oi_2
X_3463_ d7.saw_temp\[3\] net12 vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2414_ _1713_ d9.count\[0\] d9.count\[1\] vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__o21ai_1
X_3394_ d2.saw_temp\[2\] _0329_ _0300_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a21oi_1
X_2345_ d7.count\[0\] d7.count\[1\] d7.count\[2\] vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2276_ _1906_ vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4015_ _1571_ _1573_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ d2.count\[3\] d2.count\[4\] _1787_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__and3_1
X_2061_ _1727_ d1.count\[4\] vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ d1.count\[0\] _1777_ _0553_ _1719_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2894_ d6.saw_temp\[4\] d6.saw_temp\[3\] _0503_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3515_ d13.saw_temp\[7\] _0971_ _0862_ d13.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1
+ _1079_ sky130_fd_sc_hd__o22a_1
X_3446_ d3.saw_temp\[3\] _0348_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__nand2_1
X_3377_ d11.saw_temp\[2\] _0334_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _1727_ d7.count\[2\] d7.count\[3\] vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2259_ _1894_ vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3300_ _0301_ _0635_ _0307_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__a21oi_2
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ clknet_leaf_30_clk d5.nxt_count\[1\] net29 vssd1 vssd1 vccd1 vccd1 d5.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _0760_ _0796_ _0751_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__o21a_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ d6.saw_temp\[0\] _0346_ _0683_ _0310_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a31o_1
X_2113_ _1774_ _1776_ _1778_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__a31o_1
X_3093_ d11.saw_temp\[4\] d11.saw_temp\[2\] d11.saw_temp\[1\] _0334_ vssd1 vssd1 vccd1
+ vccd1 _0660_ sky130_fd_sc_hd__o31a_1
XFILLER_0_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2044_ _1712_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__inv_6
Xfanout29 net30 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_4
X_3995_ _1470_ _1488_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__or2b_1
X_2946_ d8.saw_temp\[1\] d8.saw_temp\[2\] _0541_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and3_1
X_2877_ net105 _0492_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4478_ clknet_leaf_17_clk _0137_ net39 vssd1 vssd1 vccd1 vccd1 em0.u1.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3429_ _0801_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__xor2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2800_ d3.count\[9\] _1714_ _1732_ d3.count\[6\] vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__o22a_1
X_3780_ _0760_ _1340_ _0751_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2731_ _0374_ _0375_ _0388_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_54_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4401_ clknet_leaf_10_clk _0080_ net36 vssd1 vssd1 vccd1 vccd1 d10.saw_temp\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2662_ _0312_ em0.mixed_sample\[6\] em0.mixed_sample\[5\] _0314_ _0323_ vssd1 vssd1
+ vccd1 vccd1 _0324_ sky130_fd_sc_hd__a221o_1
X_2593_ d13.count\[3\] _0270_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4332_ clknet_leaf_6_clk _0055_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
X_4263_ clknet_leaf_28_clk d4.nxt_count\[2\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3214_ em0.u1.state\[2\] em0.u1.state\[1\] vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4194_ clknet_leaf_19_clk p0.nxt_count\[2\] net39 vssd1 vssd1 vccd1 vccd1 p0.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3145_ d7.saw_temp\[6\] _0709_ _0710_ _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__or4b_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3076_ _0633_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _1381_ _1428_ _1537_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__a21boi_2
X_2929_ _0517_ _0528_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 pb[2] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3901_ d3.saw_temp\[7\] d3.saw_temp\[6\] _0348_ _0760_ vssd1 vssd1 vccd1 vccd1 _1461_
+ sky130_fd_sc_hd__and4b_1
X_3832_ _1391_ _1392_ _0723_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3763_ _1321_ _1324_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__xnor2_1
X_3694_ _0749_ _1255_ _0708_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__a21o_1
X_2714_ _0371_ _0331_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2645_ _0306_ _0300_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2576_ _1727_ d13.count\[2\] d13.count\[3\] vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__a21o_1
X_4315_ clknet_leaf_33_clk d7.nxt_count\[0\] net27 vssd1 vssd1 vccd1 vccd1 d7.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4246_ clknet_leaf_25_clk d3.nxt_count\[3\] net30 vssd1 vssd1 vccd1 vccd1 d3.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4177_ net151 _1699_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3128_ _0657_ _0694_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__nor2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ d1.saw_temp\[2\] d1.saw_temp\[1\] _0330_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2430_ _0146_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_2361_ _1973_ _1974_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
X_4100_ _1654_ _1604_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__xnor2_1
X_2292_ d6.count\[8\] _1715_ d6.count\[9\] vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__a21oi_1
X_4031_ _1446_ _1441_ _1546_ _1552_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3815_ _1374_ _1375_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3746_ _0650_ _1307_ _0760_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3677_ _1237_ _1238_ _0762_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__o21a_1
X_2628_ _0294_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__and2_1
X_2559_ net100 _0243_ _0246_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[4\] sky130_fd_sc_hd__a21oi_1
X_4229_ clknet_leaf_28_clk d2.nxt_count\[4\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3600_ d10.saw_temp\[7\] _1048_ _0674_ d10.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1
+ _1163_ sky130_fd_sc_hd__o22a_1
Xinput11 pb[5] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_1
X_3531_ _0980_ _0981_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3462_ _0622_ _1025_ _0809_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__a21o_1
X_2413_ _2012_ _2013_ _2014_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3393_ d2.saw_temp\[7\] d2.saw_temp\[1\] _0329_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2344_ _1962_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2275_ _1888_ _1904_ _1905_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__and3_1
X_4014_ _1505_ _1531_ _1572_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3729_ _0622_ _1290_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ d1.count\[2\] _1733_ _1736_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2962_ _1735_ d1.count\[1\] _1744_ _1724_ _1738_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2893_ net146 _0503_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3514_ _1075_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__xnor2_2
X_3445_ _1007_ _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__and2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _0939_ _0940_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__and2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ d7.count\[5\] _1945_ _1946_ _1872_ _1943_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__o221a_1
X_2258_ _1892_ _1893_ _1888_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__and3b_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2189_ net87 _1835_ _1837_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[8\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ d3.saw_temp\[1\] _0348_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__nand2_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _0721_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__nand2_2
X_2112_ d2.count\[7\] _1723_ _1777_ d2.count\[6\] vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__o22ai_1
X_3092_ _0301_ _0658_ _0307_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ _1718_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3994_ _1449_ _1468_ _1466_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2945_ net129 _0541_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2876_ _0493_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_1
X_4477_ clknet_leaf_17_clk net107 net39 vssd1 vssd1 vccd1 vccd1 em0.u1.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3428_ _0991_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nand2_1
X_3359_ _0749_ _0923_ _0708_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__a21o_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2730_ _0372_ _0377_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2661_ _0314_ em0.mixed_sample\[5\] em0.mixed_sample\[4\] _0291_ _0322_ vssd1 vssd1
+ vccd1 vccd1 _0323_ sky130_fd_sc_hd__o221a_1
X_4400_ clknet_leaf_2_clk net44 net26 vssd1 vssd1 vccd1 vccd1 d11.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2592_ _0272_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4331_ clknet_leaf_6_clk _0054_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4262_ clknet_leaf_28_clk d4.nxt_count\[1\] net28 vssd1 vssd1 vccd1 vccd1 d4.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3213_ _0777_ _0736_ _0737_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__or3_1
X_4193_ clknet_leaf_18_clk p0.nxt_count\[1\] net38 vssd1 vssd1 vccd1 vccd1 p0.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3144_ d7.saw_temp\[5\] net12 vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__nand2_1
X_3075_ _0634_ _0635_ _0639_ _0641_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3977_ _1427_ _1425_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__or2b_1
X_2928_ _0514_ _0516_ net192 vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2859_ d5.saw_temp\[6\] d5.saw_temp\[5\] _0480_ _0481_ vssd1 vssd1 vccd1 vccd1 _0482_
+ sky130_fd_sc_hd__and4_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 pb[3] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ _0738_ _1459_ _0768_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__o21a_1
X_3831_ d9.saw_temp\[6\] _0335_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3762_ _1135_ _1322_ _1323_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3693_ _0711_ _1254_ _0634_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2713_ _0329_ _0330_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__and3_1
X_2644_ _0306_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__clkbuf_16
X_2575_ d13.count\[1\] _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4314_ clknet_leaf_22_clk _0047_ net33 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4245_ clknet_leaf_25_clk d3.nxt_count\[2\] net30 vssd1 vssd1 vccd1 vccd1 d3.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4176_ _1699_ _1700_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3127_ _0692_ _0693_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ d1.saw_temp\[0\] _0330_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2360_ d7.count\[6\] _1971_ _1959_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__o21ai_1
X_2291_ _1910_ _1915_ _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__a31o_1
X_4030_ _1446_ _1441_ _1546_ _1552_ _1588_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__a311o_1
XFILLER_0_63_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3814_ _1369_ _1373_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__and2_1
X_3745_ _0871_ _0872_ d12.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3676_ d4.saw_temp\[5\] _0347_ _0723_ _0310_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2627_ p0.count\[6\] _0292_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2558_ net100 _0243_ _0236_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__o21ai_1
X_2489_ d10.count\[8\] _0188_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__xnor2_1
X_4228_ clknet_leaf_28_clk d2.nxt_count\[3\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4159_ _1710_ net102 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_35_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 pb[6] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
X_3530_ _1062_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__xor2_2
X_3461_ _1023_ _1024_ _0634_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__mux2_1
X_2412_ d9.count\[4\] _1725_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__or2_1
X_3392_ d2.saw_temp\[1\] _0611_ _0615_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2343_ _1959_ _1960_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__and3_1
X_2274_ d5.count\[7\] _1902_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__or2_1
X_4013_ _1530_ _1528_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3728_ _0610_ _1287_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__a21o_1
X_3659_ _1218_ _1221_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2961_ d1.count\[5\] _1720_ _1723_ d1.count\[7\] vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2892_ _0503_ _0504_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3513_ _0956_ _0967_ net20 vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__a21oi_1
X_3444_ _1003_ _1006_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _0936_ _0938_ _0934_ _0935_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__o211ai_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _1735_ d7.count\[5\] d7.count\[4\] vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__a21boi_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ d5.count\[0\] d5.count\[1\] d5.count\[2\] vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2188_ net87 _1835_ _1819_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ d6.saw_temp\[6\] _0724_ _0725_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__or4b_1
Xhold1 m0.synco.delay vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ d11.saw_temp\[7\] _0334_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__and2_2
X_2111_ d2.count\[6\] _1777_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__nand2_1
X_2042_ d1.count\[9\] _1715_ _1718_ d1.count\[8\] vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3993_ _1547_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2944_ _0541_ _0542_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2875_ _0491_ _0492_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4476_ clknet_leaf_18_clk _0135_ net16 vssd1 vssd1 vccd1 vccd1 em0.u1.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3427_ _0989_ _0990_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__nand2_1
X_3358_ _0921_ _0922_ _0634_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__mux2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ d6.count\[4\] d6.count\[5\] _1929_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__and3_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ d1.saw_temp\[0\] _0623_ _0627_ _0854_ _0618_ vssd1 vssd1 vccd1 vccd1 _0855_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2660_ _0291_ em0.mixed_sample\[4\] em0.mixed_sample\[3\] _0315_ _0321_ vssd1 vssd1
+ vccd1 vccd1 _0322_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2591_ _0270_ _0271_ _0266_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__and3b_1
X_4330_ clknet_leaf_7_clk _0053_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_1
X_4261_ clknet_leaf_28_clk net75 net28 vssd1 vssd1 vccd1 vccd1 d4.count\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3212_ _0327_ em0.u1.state\[1\] vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__nor2_2
X_4192_ clknet_leaf_19_clk p0.nxt_count\[0\] net39 vssd1 vssd1 vccd1 vccd1 p0.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3143_ d7.saw_temp\[3\] d7.saw_temp\[0\] net12 vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__o21a_1
X_3074_ d13.saw_temp\[0\] _0344_ _0640_ _0309_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3976_ _1489_ _1535_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2927_ net94 _0526_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2858_ d5.saw_temp\[2\] d5.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__and2_1
X_2789_ d2.saw_temp\[5\] _0430_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4459_ clknet_leaf_4_clk _0118_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3830_ d9.saw_temp\[7\] _0686_ _0688_ d9.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 _1391_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3761_ _1210_ _1212_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__nor2_1
X_2712_ _0346_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a21bo_1
X_3692_ _0713_ _0812_ d7.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2643_ s0.type_switch\[1\] vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__buf_4
X_2574_ d13.count\[1\] _1723_ _1777_ d13.count\[0\] vssd1 vssd1 vccd1 vccd1 _0257_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4313_ clknet_leaf_20_clk _0046_ net39 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4244_ clknet_leaf_25_clk d3.nxt_count\[1\] net30 vssd1 vssd1 vccd1 vccd1 d3.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_4175_ net242 _1691_ _1698_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__nor3_1
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3126_ _0679_ _0691_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ d1.saw_temp\[5\] d1.saw_temp\[4\] d1.saw_temp\[3\] _0330_ vssd1 vssd1 vccd1
+ vccd1 _0624_ sky130_fd_sc_hd__o31a_1
XFILLER_0_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3959_ _0639_ _1413_ _0723_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2290_ d6.count\[8\] _1715_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3813_ _1369_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3744_ _1302_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__xor2_2
X_3675_ _0738_ _1236_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2626_ p0.count\[6\] _0292_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2557_ _0245_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2488_ _0190_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_4227_ clknet_leaf_26_clk d2.nxt_count\[2\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _1710_ em0.u1.Q\[6\] net63 _0782_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__a22o_1
X_3109_ _0640_ _0674_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__o21ba_1
X_4089_ _0326_ _1645_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 pb[7] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3460_ d8.saw_temp\[7\] _0917_ _0702_ d8.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _1024_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2411_ d9.count\[4\] _1725_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__nand2_1
X_3391_ _0848_ _0858_ _0857_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a21bo_1
X_2342_ d7.count\[0\] d7.count\[1\] vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__nand2_1
X_4012_ _1569_ _1570_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__or2_1
X_2273_ d5.count\[7\] _1902_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3727_ d2.saw_temp\[4\] _0611_ _0615_ _1288_ _0618_ vssd1 vssd1 vccd1 vccd1 _1289_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3658_ _1219_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__and2_1
X_3589_ _1146_ _1151_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__nand2_1
X_2609_ _0284_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2960_ d1.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2891_ d6.saw_temp\[1\] _0502_ net171 vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3512_ _0307_ _0960_ _0965_ _0620_ _0630_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__a2111oi_1
X_3443_ _1003_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__nand2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _0934_ _0935_ _0936_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__a211o_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _1718_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__inv_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ d5.count\[0\] d5.count\[1\] d5.count\[2\] vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2187_ _1835_ _1836_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[7\] sky130_fd_sc_hd__nor2_1
XFILLER_0_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2110_ _1732_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__buf_6
Xhold2 m0.syncy.delay vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _0655_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__or2_1
X_2041_ _1717_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__buf_6
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3992_ _1710_ net56 _0782_ em0.u1.R\[15\] _1551_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2943_ d8.saw_temp\[0\] _0531_ _0540_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__nor3_1
X_2874_ d5.saw_temp\[5\] _0490_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4475_ clknet_leaf_23_clk net64 net33 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3426_ _0989_ _0990_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__or2_1
X_3357_ d7.saw_temp\[7\] _0811_ _0713_ d7.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0922_
+ sky130_fd_sc_hd__o22a_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ net138 _1929_ _1932_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[4\] sky130_fd_sc_hd__a21oi_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ d1.saw_temp\[7\] _0625_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__or2_1
X_2239_ d5.count\[2\] _1729_ d5.count\[3\] vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2590_ d13.count\[0\] d13.count\[1\] d13.count\[2\] vssd1 vssd1 vccd1 vccd1 _0271_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4260_ clknet_leaf_33_clk _0023_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
X_4191_ _1691_ _1708_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__nor2_1
X_3211_ _0736_ _0737_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o21ai_1
X_3142_ d7.saw_temp\[4\] d7.saw_temp\[2\] d7.saw_temp\[1\] net12 vssd1 vssd1 vccd1
+ vccd1 _0709_ sky130_fd_sc_hd__o31a_1
X_3073_ _0610_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3975_ _1532_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2926_ _0526_ _0527_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2857_ d5.saw_temp\[4\] d5.saw_temp\[3\] d5.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1
+ _0480_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2788_ _0429_ _0430_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__nor2_1
X_4458_ clknet_leaf_6_clk _0117_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_1
X_3409_ _0968_ _0973_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__xnor2_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ clknet_leaf_4_clk _0078_ net27 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3760_ _1210_ _1212_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2711_ _0327_ net147 _0369_ _0370_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
X_3691_ _0749_ _1252_ _0809_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2642_ _0305_ vssd1 vssd1 vccd1 vccd1 s0.next_q\[0\] sky130_fd_sc_hd__clkbuf_1
X_2573_ d13.count\[7\] _1717_ _1722_ d13.count\[6\] vssd1 vssd1 vccd1 vccd1 _0256_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4312_ clknet_leaf_20_clk _0045_ net39 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4243_ clknet_leaf_27_clk d3.nxt_count\[0\] net30 vssd1 vssd1 vccd1 vccd1 d3.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_4174_ _1691_ _1698_ d9.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__o21a_1
X_3125_ _0679_ _0691_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__nor2_1
X_3056_ d1.saw_temp\[7\] _0330_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3958_ _1516_ _1517_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__xnor2_2
X_2909_ d7.saw_temp\[4\] d7.saw_temp\[3\] d7.saw_temp\[0\] _0515_ vssd1 vssd1 vccd1
+ vccd1 _0516_ sky130_fd_sc_hd__and4_1
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3889_ _0747_ _1342_ _1347_ _1348_ _1352_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3812_ _0750_ _1372_ _0722_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__a21o_1
X_3743_ _0750_ _1304_ _0866_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__a21o_1
X_3674_ _0759_ _1235_ d4.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2625_ _0292_ net122 vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2556_ _0243_ _0244_ _0236_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__and3b_1
X_2487_ _0172_ _0188_ _0189_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4226_ clknet_leaf_26_clk d2.nxt_count\[1\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4157_ _1710_ em0.u1.Q\[5\] net88 _0782_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__a22o_1
X_3108_ d10.saw_temp\[0\] _0336_ _0640_ _0309_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__a31o_1
X_4088_ em0.u1.R\[17\] _1644_ _1609_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__mux2_1
X_3039_ _0198_ _0594_ _0589_ _0592_ d11.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0607_
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 pb[8] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_1
XFILLER_0_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2410_ d9.count\[5\] _1723_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__xnor2_1
X_3390_ _0950_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__xnor2_2
X_2341_ d7.count\[0\] d7.count\[1\] vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__or2_1
X_2272_ _1902_ net163 vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
X_4011_ _1566_ _1567_ _1568_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3726_ d2.saw_temp\[7\] d2.saw_temp\[4\] _0329_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3657_ _0998_ _1105_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__or2b_1
X_2608_ _0266_ _0282_ _0283_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3588_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__inv_2
X_2539_ d12.count\[4\] _1723_ _1777_ d12.count\[3\] vssd1 vssd1 vccd1 vccd1 _0231_
+ sky130_fd_sc_hd__o22a_1
X_4209_ clknet_leaf_32_clk s0.next_q\[1\] net31 vssd1 vssd1 vccd1 vccd1 s0.type_switch\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2890_ d6.saw_temp\[2\] d6.saw_temp\[1\] _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3511_ _1073_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__and2b_1
X_3442_ _0750_ _1005_ _0762_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_69_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _0937_ _0821_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__nor2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _1720_ _1943_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _1891_ vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2186_ net209 _1833_ _1819_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3709_ _0664_ _0829_ d11.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 m0.edgy.in vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _1712_ _1716_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3991_ _1549_ _1550_ _0779_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2942_ _0531_ _0540_ d8.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__o21a_1
X_2873_ d5.saw_temp\[5\] _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4474_ clknet_leaf_23_clk net89 net33 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3425_ _0803_ _0890_ _0888_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__o21a_1
X_3356_ d7.saw_temp\[2\] net12 vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__nand2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ d6.count\[4\] _1929_ _1922_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__o21ai_1
X_3287_ d1.saw_temp\[1\] _0330_ _0300_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__a21oi_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ d5.count\[2\] _1733_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ _1690_ _1698_ net204 vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__a21oi_1
X_3210_ _0775_ _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__or2_1
X_3141_ _0301_ _0707_ _0307_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__a21oi_4
X_3072_ d13.saw_temp\[6\] _0636_ _0637_ _0638_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__or4b_2
XFILLER_0_89_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _1421_ _1423_ _1533_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__o21a_1
X_2925_ d7.saw_temp\[4\] d7.saw_temp\[3\] _0522_ net155 vssd1 vssd1 vccd1 vccd1 _0527_
+ sky130_fd_sc_hd__a31oi_1
X_2856_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2787_ d2.saw_temp\[4\] d2.saw_temp\[3\] _0428_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__and3_1
Xhold200 em0.u1.Q\[4\] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ clknet_leaf_6_clk _0116_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3408_ _0970_ _0972_ _0633_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__o21ai_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4388_ clknet_leaf_4_clk _0077_ net26 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _0900_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2710_ _0328_ _0368_ em0.u1.state\[2\] vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__o21a_1
X_3690_ _0700_ _1251_ _0646_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2641_ _0303_ _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__and2_1
X_2572_ d13.count\[8\] _1714_ _1718_ d13.count\[7\] vssd1 vssd1 vccd1 vccd1 _0255_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4311_ clknet_leaf_20_clk _0044_ net39 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
X_4242_ clknet_leaf_31_clk _0015_ net31 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_4173_ _2015_ _1695_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__and3_2
X_3124_ _0681_ _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3055_ _0609_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ _1408_ _1410_ _1406_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__a21bo_1
X_2908_ d7.saw_temp\[6\] d7.saw_temp\[5\] d7.saw_temp\[2\] d7.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3888_ _1338_ _1356_ _1354_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2839_ _0466_ _0467_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__nor2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3811_ _1370_ _1371_ _0683_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3742_ _0638_ _1303_ _0646_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ d4.saw_temp\[7\] _0347_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2624_ p0.count\[4\] _0289_ net121 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2555_ d12.count\[1\] d12.count\[0\] d12.count\[2\] d12.count\[3\] vssd1 vssd1 vccd1
+ vccd1 _0244_ sky130_fd_sc_hd__a31o_1
X_2486_ d10.count\[7\] _0186_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__or2_1
X_4225_ clknet_leaf_26_clk d2.nxt_count\[0\] net30 vssd1 vssd1 vccd1 vccd1 d2.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_4156_ _1710_ net58 em0.u1.Q\[5\] _0782_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__a22o_1
X_3107_ _0668_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4087_ _1600_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__xnor2_1
X_3038_ net99 _0605_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput15 pb[9] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
XFILLER_0_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2340_ net85 _1959_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_58_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2271_ net162 _1900_ _1888_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__o21ai_1
X_4010_ _1566_ _1567_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3725_ d2.saw_temp\[5\] _0329_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3656_ _1104_ _1102_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__or2b_1
X_2607_ d13.count\[7\] _0280_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3587_ _0722_ _1149_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2538_ d12.count\[5\] d12.count\[6\] _1872_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__mux2_1
X_2469_ d10.count\[1\] d10.count\[0\] d10.count\[2\] vssd1 vssd1 vccd1 vccd1 _0177_
+ sky130_fd_sc_hd__a21o_1
X_4208_ clknet_leaf_32_clk s0.next_q\[0\] net31 vssd1 vssd1 vccd1 vccd1 s0.type_switch\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ em0.mixed_sample\[2\] net78 em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1 _1681_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ _1063_ _1068_ _1072_ _1064_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3441_ _0755_ _1004_ _0760_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__mux2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _0816_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__inv_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _1872_ d7.count\[4\] vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _1888_ _1889_ _1890_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__and3_1
X_2185_ d3.count\[7\] d3.count\[6\] _1831_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3708_ _1268_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3639_ _1197_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__xor2_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 m0.edgo.in vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ _1446_ _1441_ _1548_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2941_ d8.count\[6\] _1733_ _1983_ _0533_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2872_ _0489_ _0490_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4473_ clknet_leaf_23_clk net59 net33 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[5\] sky130_fd_sc_hd__dfrtp_1
X_3424_ _0915_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__xnor2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _0749_ _0919_ _0809_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__a21o_1
X_2306_ _1931_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_3286_ _0849_ _0851_ _0306_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__o21a_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ d5.count\[3\] _1729_ _1874_ _1712_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__o22a_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2168_ d3.count\[0\] d3.count\[1\] d3.count\[2\] vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2099_ _1766_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3140_ d7.saw_temp\[7\] net12 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__and2_2
XFILLER_0_89_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3071_ d13.saw_temp\[5\] _0344_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3973_ _1397_ _1424_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__or2_1
X_2924_ d7.saw_temp\[5\] d7.saw_temp\[4\] d7.saw_temp\[3\] _0522_ vssd1 vssd1 vccd1
+ vccd1 _0526_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2855_ d5.count\[0\] _1777_ _1882_ _0474_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_60_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold201 d10.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlygate4sd3_1
X_2786_ d2.saw_temp\[3\] _0428_ net218 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__a21oi_1
X_4456_ clknet_leaf_6_clk _0115_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
X_4387_ clknet_leaf_4_clk _0076_ net26 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
X_3407_ _0646_ _0971_ _0622_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _0750_ _0902_ _0762_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__a21boi_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _0674_ _0834_ d10.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ _0301_ _0302_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2571_ _0254_ _0251_ _0236_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[8\] sky130_fd_sc_hd__a21boi_1
XFILLER_0_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4310_ clknet_leaf_19_clk _0043_ net39 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4241_ clknet_leaf_32_clk _0014_ net31 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4172_ d9.count\[2\] _1724_ _1777_ d9.count\[0\] _1696_ vssd1 vssd1 vccd1 vccd1 _1697_
+ sky130_fd_sc_hd__a221oi_1
X_3123_ _0683_ _0688_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__o21ba_1
X_3054_ _0609_ _0616_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3956_ _1514_ _1515_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2907_ _1947_ _0511_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__and3_2
XFILLER_0_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3887_ _1335_ _1436_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2838_ net182 _0463_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__nor2_1
X_2769_ _1767_ _1770_ _1771_ _1776_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4439_ clknet_leaf_16_clk _0108_ net16 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[20\] sky130_fd_sc_hd__dfrtp_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3810_ d6.saw_temp\[6\] _0346_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__nand2_1
X_3741_ _0862_ _0863_ d13.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _0751_ _1233_ _0747_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__a21boi_1
X_2623_ p0.count\[4\] p0.count\[5\] _0289_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__and3_1
X_2554_ d12.count\[1\] d12.count\[0\] d12.count\[3\] d12.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _0243_ sky130_fd_sc_hd__and4_1
X_2485_ d10.count\[7\] _0186_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4224_ clknet_leaf_16_clk _0007_ net40 vssd1 vssd1 vccd1 vccd1 em0.u1.D\[12\] sky130_fd_sc_hd__dfrtp_1
X_4155_ _1710_ net103 net58 _0782_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__a22o_1
X_3106_ d10.saw_temp\[6\] _0670_ _0671_ _0672_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__or4b_1
X_4086_ em0.u1.D\[10\] em0.u1.R\[17\] vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__xor2_1
X_3037_ _0606_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3939_ _0687_ _1392_ _0738_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput16 reset vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_4
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2270_ d5.count\[6\] _1900_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3724_ _1284_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3655_ _1111_ _1217_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__xnor2_2
X_2606_ d13.count\[7\] _0280_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3586_ _0682_ _1147_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2537_ d12.count\[8\] _1715_ d12.count\[9\] vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__a21o_1
X_2468_ d10.count\[1\] d10.count\[0\] d10.count\[2\] vssd1 vssd1 vccd1 vccd1 _0176_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ clknet_leaf_28_clk e0.next_q\[1\] net28 vssd1 vssd1 vccd1 vccd1 d1.oct_dwn\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2399_ d8.count\[6\] _2002_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__and2_1
X_4138_ _1680_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
X_4069_ _1613_ _1589_ _1626_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3440_ d4.saw_temp\[7\] _0756_ _0759_ d4.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _1004_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3371_ _0810_ _0815_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nor2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2322_ _1942_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ d5.count\[0\] d5.count\[1\] vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__nand2_1
X_2184_ _1833_ _1834_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_19_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3707_ _1267_ _1265_ _1266_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3638_ _1199_ _1200_ _0645_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__o21a_2
X_3569_ _1039_ _1115_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 em0.u1.R\[14\] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2940_ d8.count\[8\] _1805_ _1981_ _0536_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2871_ d5.saw_temp\[4\] _0488_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4472_ clknet_leaf_19_clk _0131_ net39 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[4\] sky130_fd_sc_hd__dfrtp_1
X_3423_ _0986_ _0987_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__xnor2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _0917_ _0918_ _0634_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__mux2_1
X_2305_ _1929_ _1930_ _1922_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__and3b_1
X_3285_ d2.saw_temp\[0\] _0611_ _0615_ _0850_ _0618_ vssd1 vssd1 vccd1 vccd1 _0851_
+ sky130_fd_sc_hd__o311a_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _1713_ d5.count\[0\] d5.count\[1\] vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__o21a_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2167_ _1822_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_2098_ _1745_ _1764_ _1765_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3070_ d13.saw_temp\[3\] d13.saw_temp\[0\] _0344_ vssd1 vssd1 vccd1 vccd1 _0637_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3972_ _1505_ _1531_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__xor2_2
X_2923_ net173 _0523_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2854_ d5.count\[9\] _1876_ _0475_ _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__or4_1
X_2785_ net174 _0428_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4455_ clknet_leaf_4_clk _0114_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_4
X_4386_ clknet_leaf_4_clk _0075_ net26 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_4
X_3406_ d13.saw_temp\[2\] _0344_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__nand2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _0756_ _0901_ _0646_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__mux2_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ d10.saw_temp\[7\] _0336_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__or2b_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _1860_ _1861_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
X_3199_ _0764_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2570_ net185 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4240_ clknet_leaf_32_clk _0013_ net31 vssd1 vssd1 vccd1 vccd1 d13.saw_temp\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4171_ d9.count\[2\] _1724_ _1720_ d9.count\[7\] vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__a2bb2o_1
X_3122_ d9.saw_temp\[0\] _0335_ _0682_ _0309_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3053_ d2.saw_temp\[7\] _0329_ _0300_ _0306_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_89_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ _1509_ _1513_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2906_ d7.count\[8\] _1805_ _1957_ _0512_ d7.count\[9\] vssd1 vssd1 vccd1 vccd1 _0513_
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3886_ _1445_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2837_ d4.saw_temp\[2\] _0463_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__and2_1
X_2768_ _0406_ _0415_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__nor2_1
X_2699_ _0357_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__and2_1
X_4438_ clknet_leaf_14_clk _0107_ net40 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[19\] sky130_fd_sc_hd__dfrtp_1
X_4369_ clknet_leaf_17_clk net41 net38 vssd1 vssd1 vccd1 vccd1 em0.u1.state\[0\] sky130_fd_sc_hd__dfstp_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3740_ _1299_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3671_ _0742_ _1232_ _0760_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__mux2_1
X_2622_ _0291_ _0289_ vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[4\] sky130_fd_sc_hd__xnor2_1
X_2553_ _0242_ vssd1 vssd1 vccd1 vccd1 d12.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2484_ _0186_ _0187_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
X_4223_ clknet_leaf_15_clk _0006_ net40 vssd1 vssd1 vccd1 vccd1 em0.u1.D\[11\] sky130_fd_sc_hd__dfrtp_1
X_4154_ _1710_ net78 em0.u1.Q\[3\] _0782_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__a22o_1
X_3105_ d10.saw_temp\[5\] _0336_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nand2_1
X_4085_ _1639_ _1641_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__xnor2_1
X_3036_ _0604_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3938_ _1493_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3869_ _1315_ _1313_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3723_ _1279_ _1283_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3654_ _1215_ _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2605_ _0280_ _0281_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3585_ d6.saw_temp\[4\] _0346_ _0640_ _0309_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a31o_1
X_2536_ _0228_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_2467_ _0175_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_4206_ clknet_leaf_28_clk e0.next_q\[0\] net28 vssd1 vssd1 vccd1 vccd1 d1.oct_dwn\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2398_ _2002_ _2003_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
X_4137_ net179 net92 em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__mux2_1
X_4068_ _1624_ _1625_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__or2_1
X_3019_ d11.saw_temp\[4\] d11.saw_temp\[3\] d11.saw_temp\[0\] _0593_ vssd1 vssd1 vccd1
+ vccd1 _0594_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3370_ _0916_ _0845_ _0933_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nand3_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _1920_ _1921_ _1941_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__and3_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ d5.count\[0\] d5.count\[1\] vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2183_ net249 _1831_ _1819_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3706_ _1265_ _1266_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3637_ d12.saw_temp\[4\] _0340_ _0683_ _0310_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3568_ _1126_ _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2519_ _0215_ _0216_ _0208_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__and3b_1
X_3499_ d2.saw_temp\[7\] _0329_ _0301_ _0306_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 _0103_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2870_ net229 _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4471_ clknet_leaf_19_clk net79 net39 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3422_ _0884_ _0886_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__nor2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ d8.saw_temp\[7\] _0805_ _0702_ d8.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0918_
+ sky130_fd_sc_hd__o22a_1
X_2304_ d6.count\[1\] d6.count\[0\] d6.count\[2\] d6.count\[3\] vssd1 vssd1 vccd1
+ vccd1 _1930_ sky130_fd_sc_hd__a31o_1
X_3284_ d2.saw_temp\[7\] _0613_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__or2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _1872_ d5.count\[4\] d5.count\[5\] _1735_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__o211a_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _1819_ _1820_ _1821_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__and3_1
X_2097_ d1.count\[9\] d1.count\[8\] _1761_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2999_ net233 _0575_ net18 vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__nor3_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3971_ _1528_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__xnor2_2
X_2922_ _0525_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2853_ d5.count\[8\] _1715_ _1871_ _1885_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2784_ _0427_ _0428_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4454_ clknet_leaf_6_clk _0113_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4385_ clknet_leaf_4_clk _0074_ net26 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
X_3405_ _0682_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__nor2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ d4.saw_temp\[7\] _0788_ _0759_ d4.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0901_
+ sky130_fd_sc_hd__o22a_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ d10.saw_temp\[1\] _0336_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__nand2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ net157 _1857_ _1850_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__o21ai_1
X_3198_ _0748_ _0763_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__and2_1
X_2149_ d3.count\[9\] _1715_ _1718_ d3.count\[8\] vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _1692_ _2011_ _1693_ _1694_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__and4b_1
X_3121_ _0680_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3052_ _0618_ _0613_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3954_ _1509_ _1513_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2905_ d7.count\[1\] _1723_ _1777_ d7.count\[0\] _1955_ vssd1 vssd1 vccd1 vccd1 _0512_
+ sky130_fd_sc_hd__a221o_1
X_3885_ _1437_ _1439_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__nor2_1
X_2836_ _0463_ _0465_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__nor2_1
X_2767_ _0405_ _0403_ d13.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2698_ _0335_ _0356_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__nand2_1
X_4437_ clknet_leaf_15_clk _0106_ net40 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[18\] sky130_fd_sc_hd__dfrtp_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ clknet_leaf_7_clk _0071_ net37 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ clknet_leaf_3_clk d6.nxt_count\[2\] net26 vssd1 vssd1 vccd1 vccd1 d6.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3319_ _0882_ _0883_ _0695_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3670_ _0744_ _0784_ d5.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2621_ net225 vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__inv_2
X_2552_ _0236_ _0240_ _0241_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4222_ clknet_leaf_17_clk _0005_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.D\[10\] sky130_fd_sc_hd__dfrtp_1
X_2483_ net193 _0184_ _0172_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__o21ai_1
X_4153_ _1710_ net92 net78 _0782_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__a22o_1
X_3104_ d10.saw_temp\[3\] d10.saw_temp\[0\] _0336_ vssd1 vssd1 vccd1 vccd1 _0671_
+ sky130_fd_sc_hd__o21a_1
X_4084_ _1613_ _1589_ _1640_ _1624_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__a31o_1
X_3035_ d11.saw_temp\[5\] _0603_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3937_ _1495_ _1496_ _0669_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3868_ _1381_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__xnor2_1
X_2819_ _0451_ _0452_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__nor2_1
X_3799_ d8.saw_temp\[6\] _0337_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__nand2_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3722_ _1279_ _1283_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3653_ _1112_ _1113_ _1214_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2604_ d13.count\[6\] _0278_ _0266_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3584_ d6.saw_temp\[7\] _1034_ _0728_ d6.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 _1147_
+ sky130_fd_sc_hd__o22a_1
X_2535_ _0208_ _0227_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__and2_1
X_2466_ _0172_ _0173_ _0174_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__and3_1
X_4205_ clknet_leaf_28_clk net53 vssd1 vssd1 vccd1 vccd1 m0.edgy.in sky130_fd_sc_hd__dfxtp_1
X_2397_ d8.count\[5\] _2000_ _1990_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__o21ai_1
X_4136_ _1679_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
X_4067_ _1614_ _1615_ _1623_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__a21oi_1
X_3018_ d11.saw_temp\[6\] d11.saw_temp\[5\] d11.saw_temp\[2\] d11.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ d6.count\[8\] _1938_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__xnor2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ net82 _1888_ vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
X_2182_ d3.count\[6\] _1831_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3705_ _1141_ _1145_ _1152_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3636_ _0683_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3567_ _1128_ _1129_ _0767_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__o21a_1
X_2518_ d11.count\[3\] _0212_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__or2_1
X_3498_ _1060_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nand2_2
X_2449_ _2023_ _0159_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__and2_1
X_4119_ d12.saw_temp\[7\] _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7 em0.u1.Q\[4\] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ clknet_leaf_18_clk _0129_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.Q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3421_ _0941_ _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__xnor2_1
X_3352_ d8.saw_temp\[2\] _0337_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2303_ d6.count\[1\] d6.count\[0\] d6.count\[3\] d6.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _1929_ sky130_fd_sc_hd__and4_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ d2.saw_temp\[1\] _0329_ _0300_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__a21oi_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _1713_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__buf_6
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ d3.count\[0\] d3.count\[1\] vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2096_ d1.count\[8\] _1761_ d1.count\[9\] vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2998_ _0575_ net18 d10.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3619_ _0620_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _1416_ _1420_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__a21oi_2
X_2921_ _0523_ _0524_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2852_ _1945_ _1877_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__nor2_1
X_2783_ d2.saw_temp\[2\] d2.saw_temp\[1\] _0426_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4453_ clknet_leaf_6_clk _0112_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3404_ d13.saw_temp\[7\] _0861_ _0862_ d13.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1
+ _0969_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4384_ clknet_leaf_5_clk _0073_ net26 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _0750_ _0899_ _0747_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__a21boi_1
X_3266_ _0622_ _0831_ _0659_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__a21o_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ d4.count\[3\] d4.count\[4\] _1854_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__and3_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3197_ _0748_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__nor2_1
X_2148_ _1715_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__clkbuf_16
X_2079_ d1.count\[3\] _1749_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3120_ d9.saw_temp\[6\] _0684_ _0685_ _0686_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__or4b_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3051_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3953_ _0749_ _1511_ _1512_ _0630_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__a31o_1
X_3884_ _1441_ _1443_ _1444_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__a21o_1
X_2904_ _0509_ _1726_ _1949_ _0510_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__o211a_1
X_2835_ _0464_ _0462_ d4.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2766_ net115 _0413_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__xnor2_1
X_2697_ _0335_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__or2_1
X_4436_ clknet_leaf_15_clk _0105_ net40 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4367_ clknet_leaf_7_clk _0070_ net37 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3318_ _0695_ _0882_ _0883_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ clknet_leaf_3_clk d6.nxt_count\[1\] net26 vssd1 vssd1 vccd1 vccd1 d6.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_3249_ _0749_ _0814_ _0708_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _0289_ _0290_ vssd1 vssd1 vccd1 vccd1 p0.nxt_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2551_ d12.count\[1\] d12.count\[0\] d12.count\[2\] vssd1 vssd1 vccd1 vccd1 _0241_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2482_ d10.count\[6\] _0184_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4221_ clknet_leaf_17_clk _0004_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.D\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4152_ _1710_ em0.u1.Q\[0\] net92 _0782_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a22o_1
X_3103_ d10.saw_temp\[4\] d10.saw_temp\[2\] d10.saw_temp\[1\] _0336_ vssd1 vssd1 vccd1
+ vccd1 _0670_ sky130_fd_sc_hd__o31a_1
X_4083_ _1625_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__inv_2
X_3034_ d11.saw_temp\[5\] _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3936_ _0723_ _0668_ _1387_ _0750_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__o31a_1
X_3867_ _1425_ _1427_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__xnor2_2
X_3798_ d8.saw_temp\[7\] _0700_ _0702_ d8.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 _1359_
+ sky130_fd_sc_hd__o22a_1
X_2818_ d3.saw_temp\[5\] d3.saw_temp\[4\] _0450_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2749_ d13.saw_temp\[6\] d13.saw_temp\[5\] d13.saw_temp\[2\] d13.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4419_ clknet_leaf_9_clk _0088_ net36 vssd1 vssd1 vccd1 vccd1 d11.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _1282_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3652_ _1112_ _1113_ _1214_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__o21ai_1
X_3583_ _1141_ _1145_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__xor2_1
X_2603_ d13.count\[6\] _0278_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2534_ d11.count\[8\] _0224_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__xnor2_1
X_2465_ d10.count\[1\] d10.count\[0\] vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__nand2_1
X_4204_ clknet_leaf_13_clk net52 vssd1 vssd1 vccd1 vccd1 m0.edgo.in sky130_fd_sc_hd__dfxtp_1
X_2396_ d8.count\[5\] d8.count\[4\] _1997_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__and3_1
X_4135_ net190 em0.u1.Q\[0\] em0.u1.state\[3\] vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__mux2_1
X_4066_ _1614_ _1615_ _1623_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__and3_1
X_3017_ d11.count\[8\] _1715_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__o21a_1
Xwire21 _1076_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3919_ _1477_ _1478_ _0708_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ d5.count\[8\] _1805_ _1887_ net228 vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__a211oi_4
X_2181_ _1831_ _1832_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_87_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3704_ _1167_ _1175_ _1263_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3635_ d12.saw_temp\[7\] _1085_ _0871_ d12.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1
+ _1198_ sky130_fd_sc_hd__o22a_1
X_3566_ d3.saw_temp\[4\] _0348_ _0738_ _0310_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__a31o_1
X_3497_ _1054_ _1059_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__or2_1
X_2517_ d11.count\[3\] _0212_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__and2_1
X_2448_ d9.count\[8\] _0156_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2379_ d8.count\[8\] _1805_ _1989_ d8.count\[9\] vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4118_ d12.saw_temp\[4\] d12.saw_temp\[3\] d12.saw_temp\[0\] _1669_ vssd1 vssd1 vccd1
+ vccd1 _1670_ sky130_fd_sc_hd__and4_1
X_4049_ em0.u1.R\[22\] _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 _0132_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3420_ _0983_ _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__xnor2_1
X_3351_ _0832_ _0837_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2302_ _1928_ vssd1 vssd1 vccd1 vccd1 d6.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _0621_ _0631_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__nor2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _1735_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__nor2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ d3.count\[0\] d3.count\[1\] vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__nand2_1
X_2095_ net109 _1761_ _1763_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[8\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2997_ d10.count\[5\] _1729_ _0168_ _0576_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3618_ _0640_ _1179_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__o21ba_1
X_3549_ _1098_ _1100_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2920_ d7.saw_temp\[3\] _0522_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__or2_1
X_2851_ d5.count\[8\] _1805_ _1735_ d5.count\[1\] vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__a2bb2o_1
X_2782_ d2.saw_temp\[1\] _0426_ net207 vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4452_ clknet_leaf_6_clk _0111_ net35 vssd1 vssd1 vccd1 vccd1 d12.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3403_ _0956_ _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__xor2_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4383_ clknet_leaf_5_clk _0072_ net26 vssd1 vssd1 vccd1 vccd1 d1.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _0897_ _0898_ _0760_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__mux2_1
X_3265_ _0828_ _0830_ _0634_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__mux2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _1859_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _0751_ _0761_ _0762_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__a21bo_1
X_2147_ _1804_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2078_ _1752_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _0300_ _0306_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3952_ _0560_ _1510_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__nand2_1
X_2903_ d7.count\[6\] _1733_ _1950_ d7.count\[3\] _1948_ vssd1 vssd1 vccd1 vccd1 _0510_
+ sky130_fd_sc_hd__o221a_1
X_3883_ em0.u1.state\[1\] em0.u1.R\[13\] net56 _0782_ vssd1 vssd1 vccd1 vccd1 _1444_
+ sky130_fd_sc_hd__a22o_1
X_2834_ d4.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2765_ _0414_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2696_ _0354_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__and2_1
X_4435_ clknet_leaf_14_clk _0104_ net40 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ clknet_leaf_7_clk _0069_ net35 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3317_ _0880_ _0881_ _0847_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__o21ai_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ clknet_leaf_3_clk d6.nxt_count\[0\] net26 vssd1 vssd1 vccd1 vccd1 d6.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_3248_ _0811_ _0813_ _0646_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__mux2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ d5.saw_temp\[0\] _0328_ _0723_ _0310_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__a31o_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2550_ d12.count\[1\] d12.count\[0\] d12.count\[2\] vssd1 vssd1 vccd1 vccd1 _0240_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_50_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2481_ _0184_ _0185_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
X_4220_ clknet_leaf_17_clk _0003_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.D\[8\] sky130_fd_sc_hd__dfrtp_1
X_4151_ net131 _0782_ _1609_ _1710_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__a22o_1
X_3102_ _0301_ _0668_ _0307_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__a21oi_4
X_4082_ _1635_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3033_ _0602_ _0603_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3935_ _0668_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3866_ _1286_ _1312_ _1426_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3797_ _1257_ _1258_ _1262_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nor3_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2817_ d3.saw_temp\[4\] _0450_ net241 vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__a21oi_1
X_2748_ _0260_ _0259_ _0402_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__and3_1
X_4418_ clknet_leaf_38_clk net43 net22 vssd1 vssd1 vccd1 vccd1 d12.count\[9\] sky130_fd_sc_hd__dfrtp_1
X_2679_ _0336_ _0337_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__nand2_1
X_4349_ clknet_leaf_14_clk _0062_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3720_ _0750_ _1281_ _0681_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ _1135_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__xnor2_1
X_3582_ _0749_ _1143_ _1144_ _0708_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__a31o_1
X_2602_ _0278_ _0279_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
X_2533_ _0226_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_2464_ d10.count\[1\] d10.count\[0\] vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4203_ clknet_leaf_28_clk net2 vssd1 vssd1 vccd1 vccd1 m0.syncy.delay sky130_fd_sc_hd__dfxtp_1
X_2395_ _2000_ _2001_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4134_ _1671_ _1678_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__nor2_1
X_4065_ _1556_ _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__xor2_1
X_3016_ d11.count\[7\] _1718_ _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3918_ _0723_ _0707_ _1365_ _0750_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_31_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3849_ _1189_ _1191_ _1299_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2180_ net184 _1829_ _1819_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3703_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3634_ _1192_ _1196_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3565_ _0738_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3496_ _1054_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__nand2_1
X_2516_ _0214_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_2447_ _0158_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2378_ d8.count\[8\] _1805_ _1985_ _1987_ _1988_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__o221a_1
X_4117_ d12.saw_temp\[6\] d12.saw_temp\[5\] d12.saw_temp\[2\] d12.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4048_ em0.u1.R\[21\] _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold9 em0.u1.count\[2\] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3350_ _0896_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__xnor2_1
X_2301_ _1922_ _1926_ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__and3_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _0845_ _0846_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__nand2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _1727_ d5.count\[6\] d5.count\[7\] vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ net73 _1819_ vssd1 vssd1 vccd1 vccd1 d3.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
X_2094_ d1.count\[8\] _1761_ _1745_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _0577_ _0171_ _0578_ _0161_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__or4b_1
XFILLER_0_28_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3617_ d2.saw_temp\[4\] _0329_ _0610_ _0309_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__a31o_1
X_3548_ _0999_ _1017_ _1015_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a21o_1
X_3479_ _1019_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2850_ _0457_ _0473_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2781_ _0425_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4451_ clknet_leaf_27_clk net42 net28 vssd1 vssd1 vccd1 vccd1 d13.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3402_ _0961_ _0966_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__xnor2_2
X_4382_ clknet_leaf_0_clk net45 net23 vssd1 vssd1 vccd1 vccd1 d10.count\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ d5.saw_temp\[7\] _0783_ _0744_ d5.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0898_
+ sky130_fd_sc_hd__o22a_1
X_3264_ _0664_ _0829_ d11.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__mux2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2215_ _1857_ _1858_ _1850_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__and3b_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3195_ d4.saw_temp\[7\] _0301_ _0347_ _0307_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__a31o_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2146_ _1783_ _1802_ _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__and3_1
X_2077_ _1745_ _1750_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2979_ net169 _0565_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3951_ _0634_ _0627_ _1510_ _0623_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ d7.count\[6\] vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3882_ _1442_ _1440_ _0779_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__o21a_1
X_2833_ _0457_ _0461_ d4.saw_temp\[1\] d4.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0463_
+ sky130_fd_sc_hd__o211a_1
X_2764_ _0412_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2695_ _0343_ _0353_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__or2_1
X_4434_ clknet_leaf_16_clk net57 net40 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4365_ clknet_leaf_7_clk _0068_ net36 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3316_ _0847_ _0880_ _0881_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ clknet_leaf_31_clk _0039_ net31 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
X_3247_ _0713_ _0812_ d7.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__mux2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _0738_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nor2_1
X_2129_ _1791_ _1792_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[3\] sky130_fd_sc_hd__nor2_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2480_ net214 _0182_ _0172_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4150_ _1686_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
X_3101_ d10.saw_temp\[7\] _0336_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__and2_2
X_4081_ _1636_ _1637_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__nor2_1
X_3032_ d11.saw_temp\[4\] d11.saw_temp\[3\] _0601_ vssd1 vssd1 vccd1 vccd1 _0603_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3934_ _0673_ _1387_ _0723_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3865_ _1310_ _1311_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__nor2_1
X_2816_ net150 _0450_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__xor2_1
X_3796_ _1338_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2747_ _0257_ _0396_ _0400_ _0401_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2678_ _0336_ _0337_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__or2_1
X_4417_ clknet_leaf_38_clk d12.nxt_count\[8\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4348_ clknet_leaf_14_clk _0061_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4279_ clknet_leaf_30_clk net83 net28 vssd1 vssd1 vccd1 vccd1 d5.count\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _1210_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__xnor2_1
X_3581_ d7.saw_temp\[4\] net12 _0683_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__nand3_1
X_2601_ d13.count\[5\] _0276_ _0266_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__o21ai_1
X_2532_ _0208_ _0224_ _0225_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__and3_1
X_4202_ clknet_leaf_13_clk net1 vssd1 vssd1 vccd1 vccd1 m0.synco.delay sky130_fd_sc_hd__dfxtp_1
X_2463_ net86 _0172_ vssd1 vssd1 vccd1 vccd1 d10.nxt_count\[0\] sky130_fd_sc_hd__nand2_1
X_2394_ net236 _1997_ _1990_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4133_ _1670_ _1668_ d12.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a21oi_1
X_4064_ _1620_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__xor2_1
X_3015_ d11.count\[1\] _1732_ _0201_ d11.count\[0\] vssd1 vssd1 vccd1 vccd1 _0590_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3917_ _0707_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__nand2_1
X_3848_ _1300_ _1297_ _1298_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__o21ba_1
X_3779_ d5.saw_temp\[6\] _0328_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3702_ _1167_ _1175_ _1263_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__a21o_1
X_3633_ _0633_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__nand2_1
X_3564_ d3.saw_temp\[7\] _1010_ _0793_ d3.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 _1127_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3495_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__inv_2
X_2515_ _0212_ _0213_ _0208_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__and3b_1
X_2446_ _2023_ _0156_ _0157_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__and3_1
X_4116_ d12.count\[7\] _1720_ _1667_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__a21oi_2
X_2377_ _1721_ d8.count\[7\] vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4047_ em0.u1.R\[20\] _1592_ _1605_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__or3b_1
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3280_ _0838_ _0844_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__or2_1
X_2300_ d6.count\[1\] d6.count\[0\] d6.count\[2\] vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__a21o_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _1869_ _1866_ _1850_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[8\] sky130_fd_sc_hd__a21boi_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2162_ d3.count\[9\] _1805_ _1806_ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__o22ai_4
X_2093_ _1761_ _1762_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[7\] sky130_fd_sc_hd__nor2_1
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2995_ _1735_ d10.count\[3\] _0162_ _0173_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3616_ d2.saw_temp\[3\] _0611_ _0615_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o31a_1
XFILLER_0_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3547_ _1710_ net96 _0782_ em0.u1.R\[11\] _1110_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3478_ _1040_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__nor2_1
X_2429_ _2027_ _2028_ _2023_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__and3b_1
XFILLER_0_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2780_ net170 _0425_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4450_ clknet_leaf_27_clk d13.nxt_count\[8\] net30 vssd1 vssd1 vccd1 vccd1 d13.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_4381_ clknet_leaf_0_clk d10.nxt_count\[8\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3401_ _0630_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3332_ d5.saw_temp\[2\] _0328_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ d11.saw_temp\[7\] _0334_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__or2b_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ d4.count\[3\] _1854_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__or2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _0752_ _0759_ _0760_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__mux2_1
X_2145_ d2.count\[9\] d2.count\[8\] _1799_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2076_ d1.count\[0\] d1.count\[1\] d1.count\[2\] vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2978_ _0565_ _0566_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 d4.count\[5\] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dlygate4sd3_1
X_3950_ _0640_ _1403_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__nor2_1
X_2901_ _0500_ _0508_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3881_ _1327_ _1332_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2832_ net152 _0462_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2763_ d13.saw_temp\[5\] _0411_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2694_ _0343_ _0353_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__nand2_1
X_4433_ clknet_2_3__leaf_clk _0102_ net40 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4364_ clknet_leaf_8_clk _0067_ net36 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ clknet_leaf_21_clk _0038_ net31 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_2
X_3315_ _0877_ _0878_ _0879_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__a21oi_1
X_3246_ d7.saw_temp\[7\] _0333_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__or2_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3177_ _0739_ _0743_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__nand2b_2
X_2128_ net248 _1787_ _1783_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2059_ d1.count\[3\] _1729_ _1734_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__o22a_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3100_ _0659_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__or2_1
X_4080_ _1556_ _1622_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__and2b_1
X_3031_ d11.saw_temp\[3\] _0601_ net231 vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3933_ _0751_ _1491_ _1492_ _0659_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3864_ _1397_ _1424_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__xor2_2
X_2815_ _0449_ _0450_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3795_ _1354_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2746_ d13.count\[5\] _1733_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2677_ net13 vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4416_ clknet_leaf_38_clk d12.nxt_count\[7\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4347_ clknet_leaf_14_clk _0060_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_4
X_4278_ clknet_leaf_21_clk _0031_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[7\] sky130_fd_sc_hd__dfrtp_4
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _0793_ _0794_ d3.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3580_ _0682_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__or2_1
X_2600_ d13.count\[5\] d13.count\[4\] _0273_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__and3_1
X_2531_ d11.count\[7\] _0222_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__or2_1
X_4201_ clknet_leaf_28_clk net54 vssd1 vssd1 vccd1 vccd1 m0.edgy.delay sky130_fd_sc_hd__dfxtp_1
X_2462_ _0161_ _0170_ _0171_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__a21oi_4
X_2393_ d8.count\[3\] d8.count\[4\] _1994_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__and3_1
X_4132_ net101 _1677_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__xor2_1
X_4063_ _1558_ _1579_ _1578_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__a21oi_1
X_3014_ _0202_ _0194_ _0206_ _0193_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__and4b_1
XFILLER_0_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3916_ _0712_ _1365_ _0723_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3847_ _1406_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__and2_1
X_3778_ d5.saw_temp\[7\] _0742_ _0744_ d5.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 _1339_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2729_ _0386_ _0387_ net116 _0327_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_14_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3701_ _1259_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3632_ d13.saw_temp\[4\] _0344_ _0682_ _1194_ _0309_ vssd1 vssd1 vccd1 vccd1 _1195_
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_70_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3563_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__and2_1
X_3494_ _0750_ _1057_ _0681_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__a21o_1
X_2514_ _0195_ _0210_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__nand2_1
X_2445_ d9.count\[7\] _0154_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__or2_1
X_2376_ d8.count\[6\] _1733_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__a21bo_1
X_4115_ d12.count\[4\] _1723_ _1777_ d12.count\[3\] _1666_ vssd1 vssd1 vccd1 vccd1
+ _1667_ sky130_fd_sc_hd__a221o_1
X_4046_ _1592_ _1593_ _1604_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__or3_1
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ d4.count\[8\] vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2161_ _1807_ _1816_ _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__o21ba_1
X_2092_ d1.count\[7\] _1759_ _1745_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2994_ _1872_ _0163_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3615_ d2.saw_temp\[7\] d2.saw_temp\[3\] _0329_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__nand3b_1
X_3546_ _0995_ _1108_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__o21a_1
X_3477_ _1020_ _1022_ _1038_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2428_ d9.count\[0\] d9.count\[1\] d9.count\[2\] vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__a21o_1
X_2359_ d7.count\[6\] _1971_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__and2_1
X_4029_ _1585_ _1587_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4380_ clknet_leaf_0_clk d10.nxt_count\[7\] net23 vssd1 vssd1 vccd1 vccd1 d10.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3400_ _0962_ _0964_ _0307_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3331_ _0767_ _0792_ _0798_ _0787_ _0791_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__a32o_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ d11.saw_temp\[1\] _0334_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__nand2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ d4.count\[3\] _1854_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__and2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _0646_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__clkbuf_8
X_2144_ d2.count\[8\] _1799_ d2.count\[9\] vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2977_ d1.saw_temp\[1\] _0564_ net178 vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3529_ _1089_ _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold91 d10.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 em0.u1.Q\[0\] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2900_ _0497_ _0499_ net202 vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3880_ _1327_ _1332_ _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2831_ _0457_ _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2762_ d13.saw_temp\[5\] _0411_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__or2_1
X_2693_ _0345_ _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__xnor2_1
X_4432_ clknet_leaf_17_clk net62 net38 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[13\] sky130_fd_sc_hd__dfrtp_1
X_4363_ clknet_leaf_8_clk _0066_ net36 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ clknet_leaf_21_clk _0037_ net31 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_2
X_3314_ _0877_ _0878_ _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__and3_1
X_3245_ d7.saw_temp\[1\] net12 vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__nand2_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ d5.saw_temp\[6\] _0740_ _0741_ _0742_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__or4b_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2127_ d2.count\[3\] _1787_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__and2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _1712_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__buf_6
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3030_ net136 _0601_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _0723_ _0658_ _1383_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2814_ d3.saw_temp\[3\] _0448_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__and2_1
X_3794_ _1264_ _1269_ _1353_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2745_ _0255_ _0397_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__and3_1
X_2676_ net15 vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4415_ clknet_leaf_38_clk d12.nxt_count\[6\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4346_ clknet_leaf_13_clk _0059_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4277_ clknet_leaf_22_clk _0030_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ d3.saw_temp\[7\] _0348_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__or2b_1
X_3159_ d6.saw_temp\[5\] _0346_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_34_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2530_ d11.count\[7\] _0222_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__nand2_1
X_2461_ d10.count\[8\] _1715_ d10.count\[9\] vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__a21o_1
X_4200_ clknet_leaf_13_clk net55 vssd1 vssd1 vccd1 vccd1 m0.edgo.delay sky130_fd_sc_hd__dfxtp_1
X_2392_ _1999_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_4131_ d12.saw_temp\[5\] _1675_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__and2_1
X_4062_ _1562_ _1619_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__xnor2_2
X_3013_ _0575_ _0588_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3915_ _0751_ _1473_ _1474_ _0809_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3846_ _1401_ _1405_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3777_ _1241_ _1245_ _1240_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__a21bo_1
X_2728_ _0369_ _0385_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2659_ _0315_ em0.mixed_sample\[3\] em0.mixed_sample\[2\] _0316_ _0320_ vssd1 vssd1
+ vccd1 vccd1 _0321_ sky130_fd_sc_hd__o221a_1
X_4329_ clknet_leaf_7_clk _0052_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3700_ _0750_ _1261_ _0722_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3631_ _0682_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3562_ _1119_ _1123_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__or2_1
X_2513_ _0195_ _0210_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3493_ _1055_ _1056_ _0646_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2444_ d9.count\[7\] _0154_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_5_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2375_ _1721_ d8.count\[7\] vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__nand2_1
X_4114_ _0230_ _1663_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__nand3_1
X_4045_ _1594_ em0.u1.R\[18\] _1603_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3829_ _1385_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ d3.count\[8\] _1718_ _1722_ d3.count\[7\] vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__o22ai_1
X_2091_ d1.count\[7\] d1.count\[6\] _1757_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2993_ d10.count\[7\] _1720_ _1777_ d10.count\[2\] vssd1 vssd1 vccd1 vccd1 _0576_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3614_ _1175_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3545_ _0995_ _1108_ _0893_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__a21oi_1
X_3476_ _1039_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2427_ d9.count\[0\] d9.count\[1\] d9.count\[2\] vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2358_ _1971_ _1972_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2289_ _1735_ _1916_ _1913_ _1917_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__o211ai_1
X_4028_ _1448_ _1544_ _1586_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3330_ _0892_ _0894_ _0895_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__o21ai_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _0825_ _0826_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__nand2_1
X_2212_ _1856_ vssd1 vssd1 vccd1 vccd1 d4.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _0753_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__nand2_2
X_2143_ net98 _1799_ _1801_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[8\] sky130_fd_sc_hd__a21oi_1
X_2074_ d1.count\[0\] d1.count\[1\] d1.count\[2\] vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2976_ d1.saw_temp\[2\] d1.saw_temp\[1\] _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3528_ _1090_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__nor2_1
X_3459_ d8.saw_temp\[3\] _0337_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold70 p0.count\[5\] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 p0.count\[3\] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 d12.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ d4.count\[8\] _1805_ _0458_ _0460_ d4.count\[9\] vssd1 vssd1 vccd1 vccd1 _0461_
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2761_ _0410_ _0411_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2692_ _0346_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__xor2_1
XANTENNA_1 _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4431_ clknet_leaf_20_clk _0100_ net38 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[12\] sky130_fd_sc_hd__dfrtp_1
X_4362_ clknet_leaf_8_clk _0065_ net36 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ clknet_leaf_21_clk _0036_ net33 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_2
X_3313_ _0632_ _0633_ _0642_ _0655_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__a31o_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _0749_ _0808_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__a21o_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ d5.saw_temp\[5\] _0328_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__nand2_1
X_2126_ _1790_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_2057_ _1713_ d1.count\[0\] d1.count\[1\] vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__o21a_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2959_ _0531_ _0550_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ _0658_ _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3862_ _1306_ _1309_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__a21oi_2
X_2813_ net243 _0448_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__nor2_1
X_3793_ _1264_ _1269_ _1353_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2744_ d13.count\[0\] _1732_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__a21oi_1
X_2675_ net14 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__clkbuf_4
X_4414_ clknet_leaf_38_clk d12.nxt_count\[5\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4345_ clknet_leaf_13_clk _0058_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
X_4276_ clknet_leaf_22_clk _0029_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _0768_ _0772_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__nand2_2
X_3158_ d6.saw_temp\[3\] d6.saw_temp\[0\] _0346_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__o21a_1
X_2109_ _1715_ _1775_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__nand2_1
X_3089_ _0644_ _0654_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2460_ _0162_ _0169_ d10.count\[7\] _1720_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2391_ _1997_ _1998_ _1990_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__and3b_1
X_4130_ net143 _1675_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__xor2_1
X_4061_ _1617_ _1618_ _1571_ _1573_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__o2bb2a_1
X_3012_ _0574_ net18 net183 vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3914_ _0683_ _0697_ _1360_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3845_ _1401_ _1405_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__or2_1
X_3776_ _1250_ _1320_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__nor2_1
X_2727_ _0369_ _0385_ _0327_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2658_ p0.nxt_count\[0\] em0.mixed_sample\[0\] _0318_ _0319_ vssd1 vssd1 vccd1 vccd1
+ _0320_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2589_ d13.count\[0\] d13.count\[1\] d13.count\[2\] vssd1 vssd1 vccd1 vccd1 _0270_
+ sky130_fd_sc_hd__and3_1
X_4328_ clknet_leaf_7_clk _0051_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_2
X_4259_ clknet_leaf_5_clk _0022_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3630_ d13.saw_temp\[7\] _1081_ _0862_ d13.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1
+ _1193_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3561_ _1119_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2512_ _0211_ vssd1 vssd1 vccd1 vccd1 d11.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3492_ d9.saw_temp\[7\] _0951_ _0688_ d9.saw_temp\[2\] vssd1 vssd1 vccd1 vccd1 _1056_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2443_ _0154_ _0155_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_59_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2374_ _1735_ d8.count\[5\] _1733_ d8.count\[6\] _1984_ vssd1 vssd1 vccd1 vccd1 _1985_
+ sky130_fd_sc_hd__o221a_1
X_4113_ d12.count\[2\] _0229_ _0233_ _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nor4_1
X_4044_ _1594_ em0.u1.R\[18\] _1602_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3828_ _0750_ _1388_ _0669_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3759_ _1250_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2090_ _1759_ _1760_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2992_ d10.saw_temp\[7\] _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3613_ _1169_ _1174_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3544_ _1106_ _1107_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__xor2_2
X_3475_ _1020_ _1022_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2426_ _2026_ vssd1 vssd1 vccd1 vccd1 d9.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2357_ net237 _1969_ _1959_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2288_ _1777_ _1911_ _1914_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__a21oi_1
X_4027_ _1543_ _1540_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__or2b_1
XFILLER_0_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _0717_ _0732_ _0823_ _0824_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__o211ai_2
X_2211_ _1854_ _1855_ _1850_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__and3b_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ d4.saw_temp\[6\] _0754_ _0757_ _0752_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__or4b_1
X_2142_ net98 _1799_ _1783_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__o21ai_1
X_2073_ _1748_ vssd1 vssd1 vccd1 vccd1 d1.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2975_ net177 _0564_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3527_ _0976_ _0978_ _0645_ _0974_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3458_ _1021_ _0954_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__or2_1
X_3389_ _0749_ _0953_ _0681_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__a21o_1
X_2409_ _1727_ d9.count\[6\] vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 d2.count\[0\] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold71 _0293_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 d8.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 d10.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2760_ d13.saw_temp\[4\] d13.saw_temp\[3\] _0409_ vssd1 vssd1 vccd1 vccd1 _0411_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2691_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__nand2_1
X_4430_ clknet_leaf_20_clk net97 net38 vssd1 vssd1 vccd1 vccd1 em0.u1.R\[11\] sky130_fd_sc_hd__dfrtp_1
X_4361_ clknet_leaf_7_clk _0064_ net35 vssd1 vssd1 vccd1 vccd1 d8.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4292_ clknet_leaf_21_clk _0035_ net31 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_1
X_3312_ _0868_ _0869_ _0876_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3243_ _0301_ _0697_ _0307_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a21oi_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ d5.saw_temp\[3\] d5.saw_temp\[0\] _0328_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__o21a_1
X_2125_ _1783_ _1788_ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__and3_1
X_2056_ _1714_ _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__nand2_8
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2958_ _0530_ _0540_ d8.saw_temp\[7\] vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2889_ _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4270__51 vssd1 vssd1 vccd1 vccd1 _4270__51/HI net51 sky130_fd_sc_hd__conb_1
XFILLER_0_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3930_ _0663_ _1383_ _0723_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3861_ _1302_ _1305_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2812_ _0447_ _0448_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__nor2_1
X_3792_ _1348_ _1352_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__xnor2_1
X_2743_ d13.count\[8\] _1714_ _0256_ d13.count\[9\] vssd1 vssd1 vccd1 vccd1 _0398_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2674_ net4 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__clkbuf_4
X_4413_ clknet_leaf_38_clk d12.nxt_count\[4\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_4344_ clknet_leaf_13_clk _0057_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
X_4275_ clknet_leaf_22_clk _0028_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _0787_ _0791_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3157_ d6.saw_temp\[4\] d6.saw_temp\[2\] d6.saw_temp\[1\] _0346_ vssd1 vssd1 vccd1
+ vccd1 _0724_ sky130_fd_sc_hd__o31a_1
X_2108_ _1721_ d2.count\[4\] d2.count\[5\] vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__a21o_1
X_3088_ _0644_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__nor2_1
X_2039_ _1713_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2390_ d8.count\[3\] _1994_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__or2_1
X_4060_ _1569_ _1616_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3011_ net117 _0587_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3913_ _0697_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__nand2_1
X_3844_ _0622_ _1404_ _0630_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3775_ _1317_ _1319_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2726_ _0383_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__or2_1
X_2657_ _0316_ em0.mixed_sample\[2\] em0.mixed_sample\[1\] _0317_ vssd1 vssd1 vccd1
+ vccd1 _0319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2588_ _0269_ vssd1 vssd1 vccd1 vccd1 d13.nxt_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_4327_ clknet_leaf_6_clk _0050_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
X_4258_ clknet_leaf_5_clk _0021_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[5\] sky130_fd_sc_hd__dfrtp_2
X_3209_ _0767_ _0774_ _0766_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__a21oi_1
X_4189_ net119 _1705_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 d3.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3560_ _1121_ _1122_ _0762_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2511_ _0208_ _0209_ _0210_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3491_ d9.saw_temp\[3\] _0335_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2442_ net240 _0152_ _2023_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__o21ai_1
X_2373_ _1980_ _1982_ _1983_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ _1872_ d12.count\[5\] _0238_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__a21o_1
X_4043_ _1595_ em0.u1.R\[17\] _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3827_ _1386_ _1387_ _0683_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3758_ _1317_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2709_ _0328_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nand2_1
X_3689_ _0702_ _0806_ d8.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2991_ d10.saw_temp\[4\] d10.saw_temp\[3\] d10.saw_temp\[0\] _0573_ vssd1 vssd1 vccd1
+ vccd1 _0574_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3612_ _1169_ _1174_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_2
XFILLER_0_71_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3543_ _0801_ _0993_ _0991_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__o21a_1
X_3474_ _1033_ _1037_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2425_ _2023_ _2024_ _2025_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__and3_1
X_2356_ d7.count\[5\] d7.count\[4\] _1966_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__and3_1
X_2287_ _1872_ d6.count\[3\] d6.count\[4\] vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__o21a_1
X_4026_ _1553_ _1584_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ d4.count\[0\] d4.count\[1\] d4.count\[2\] vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__a21o_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _0755_ _0756_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__nand2_1
X_2141_ _1799_ _1800_ vssd1 vssd1 vccd1 vccd1 d2.nxt_count\[7\] sky130_fd_sc_hd__nor2_1
X_2072_ _1745_ _1746_ _1747_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2974_ _0551_ _0559_ _0564_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3526_ _0970_ _0972_ _0633_ _0968_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3457_ _0950_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__inv_2
X_3388_ _0951_ _0952_ _0646_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__mux2_1
X_2408_ _2010_ vssd1 vssd1 vccd1 vccd1 d8.nxt_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_2339_ _1956_ _1957_ _1958_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__o21a_2
X_4009_ _1514_ _1517_ _1515_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold50 d12.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 d2.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 p0.count\[1\] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 d6.saw_temp\[6\] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 d13.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2690_ _0347_ _0348_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ clknet_leaf_37_clk net46 net23 vssd1 vssd1 vccd1 vccd1 d9.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3311_ _0868_ _0869_ _0876_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__nand3_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ clknet_leaf_31_clk _0034_ net31 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _0805_ _0807_ _0634_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__mux2_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ d5.saw_temp\[4\] d5.saw_temp\[2\] d5.saw_temp\[1\] _0328_ vssd1 vssd1 vccd1
+ vccd1 _0740_ sky130_fd_sc_hd__o31a_1
X_2124_ d2.count\[1\] d2.count\[0\] d2.count\[2\] vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2055_ _1731_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__buf_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2957_ net133 _0547_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__xnor2_1
X_2888_ net139 _0501_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__xnor2_1
X_3509_ _1063_ _1064_ _1068_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__and4_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3860_ _1416_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2811_ d3.saw_temp\[2\] d3.saw_temp\[1\] _0446_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__and3_1
X_3791_ _1350_ _1351_ _0767_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2742_ d13.count\[4\] _1718_ _1722_ d13.count\[6\] vssd1 vssd1 vccd1 vccd1 _0397_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2673_ net12 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
X_4412_ clknet_leaf_0_clk d12.nxt_count\[3\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4343_ clknet_leaf_13_clk _0056_ net40 vssd1 vssd1 vccd1 vccd1 d7.saw_temp\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4274_ clknet_leaf_24_clk _0027_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[3\] sky130_fd_sc_hd__dfrtp_2
X_3225_ _0751_ _0790_ _0762_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__a21boi_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ _0683_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__buf_6
X_2107_ _1770_ _1771_ _1773_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__a21o_1
X_3087_ _0645_ _0653_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2038_ _1714_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__buf_6
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3989_ _1446_ _1441_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3010_ net252 _0585_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__and2_1
X_3912_ _0701_ _1360_ _0723_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3843_ _1402_ _1403_ _0640_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3774_ _1230_ _1249_ _1247_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2725_ _0363_ _0367_ _0382_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2656_ _0317_ em0.mixed_sample\[1\] vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2587_ _0266_ _0267_ _0268_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ clknet_leaf_6_clk _0049_ net35 vssd1 vssd1 vccd1 vccd1 d6.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
X_4257_ clknet_leaf_5_clk _0020_ net27 vssd1 vssd1 vccd1 vccd1 d2.saw_temp\[4\] sky130_fd_sc_hd__dfrtp_4
X_4188_ _1707_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
X_3208_ _0766_ _0767_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__and3_1
X_3139_ _0703_ _0704_ _0705_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold180 d11.saw_temp\[4\] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 d9.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3490_ _1052_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__and2_1
X_2510_ d11.count\[1\] d11.count\[0\] vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__nand2_1
X_2441_ d9.count\[6\] _0152_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2372_ _1735_ d8.count\[5\] d8.count\[4\] _1726_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__a22oi_1
X_4111_ d12.count\[8\] _1715_ _1718_ d12.count\[7\] _0231_ vssd1 vssd1 vccd1 vccd1
+ _1663_ sky130_fd_sc_hd__o221a_1
X_4042_ _1595_ em0.u1.R\[17\] _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3826_ d10.saw_temp\[6\] _0336_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ _1158_ _1209_ _1318_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2708_ _0365_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3688_ _1230_ _1249_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__xnor2_1
X_2639_ _0301_ _0302_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__nand2_1
X_4309_ clknet_leaf_19_clk _0042_ net39 vssd1 vssd1 vccd1 vccd1 d5.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2990_ d10.saw_temp\[6\] d10.saw_temp\[5\] d10.saw_temp\[2\] d10.saw_temp\[1\] vssd1
+ vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3611_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3542_ _0998_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__xnor2_2
X_3473_ _0750_ _1036_ _0722_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__a21o_1
X_2424_ d9.count\[0\] d9.count\[1\] vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2355_ _1969_ _1970_ vssd1 vssd1 vccd1 vccd1 d7.nxt_count\[4\] sky130_fd_sc_hd__nor2_1
X_2286_ _1777_ _1911_ _1913_ _1914_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__a211o_1
X_4025_ _1581_ _1583_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3809_ d6.saw_temp\[7\] _0726_ _0728_ d6.saw_temp\[5\] vssd1 vssd1 vccd1 vccd1 _1370_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ net186 _1797_ _1783_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__o21ai_1
X_2071_ d1.count\[0\] d1.count\[1\] vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2973_ _0563_ _0559_ _0551_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3525_ _1084_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__xnor2_2
X_3456_ _0945_ _0949_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__or2_1
X_3387_ d9.saw_temp\[7\] _0839_ _0688_ d9.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 _0952_
+ sky130_fd_sc_hd__o22a_1
X_2407_ _1990_ _2009_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and2_1
X_2338_ d7.count\[8\] _1805_ d7.count\[9\] vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__a21oi_1
X_2269_ _1900_ net195 vssd1 vssd1 vccd1 vccd1 d5.nxt_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4008_ _1523_ _1527_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold40 em0.u1.R\[20\] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 d10.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 em0.u1.count\[0\] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_1
Xhold62 em0.mixed_sample\[7\] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 d11.saw_temp\[1\] vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 d6.saw_temp\[3\] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _0749_ _0874_ _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__a21oi_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ clknet_leaf_31_clk _0033_ net31 vssd1 vssd1 vccd1 vccd1 d4.saw_temp\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _0702_ _0806_ d8.saw_temp\[0\] vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__mux2_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ d5.saw_temp\[7\] _0328_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__nand2_1
X_2123_ _1787_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2054_ _1712_ _1713_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2956_ _0549_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2887_ net206 _0497_ _0501_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3508_ _1069_ _1071_ _0306_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__o21ai_1
X_3439_ _0751_ _1002_ _0747_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__a21boi_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2810_ d3.saw_temp\[1\] _0446_ net224 vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__a21oi_1
X_3790_ d3.saw_temp\[6\] _0348_ _0738_ _0310_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__a31o_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2741_ d13.count\[1\] _1723_ _1718_ d13.count\[4\] vssd1 vssd1 vccd1 vccd1 _0396_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4411_ clknet_leaf_0_clk d12.nxt_count\[2\] net22 vssd1 vssd1 vccd1 vccd1 d12.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2672_ _0329_ _0330_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4342_ clknet_leaf_35_clk net47 net24 vssd1 vssd1 vccd1 vccd1 d8.count\[9\] sky130_fd_sc_hd__dfrtp_1
X_4273_ clknet_leaf_24_clk _0026_ net32 vssd1 vssd1 vccd1 vccd1 d3.saw_temp\[2\] sky130_fd_sc_hd__dfrtp_2
X_3224_ _0788_ _0789_ _0760_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__mux2_1
.ends

