module sync (
    input logic async_in, clk, nrst,
    output logic sync_sig
);
        

endmodule