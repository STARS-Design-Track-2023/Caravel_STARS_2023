* NGSPICE file created from sass_synth.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt sass_synth beat_led[0] beat_led[1] beat_led[2] beat_led[3] beat_led[4] beat_led[5]
+ beat_led[6] beat_led[7] cs hwclk mode_out[0] mode_out[1] multi[0] multi[1] multi[2]
+ multi[3] n_rst note1[0] note1[1] note1[2] note1[3] note2[0] note2[1] note2[2] note2[3]
+ note3[0] note3[1] note3[2] note3[3] note4[0] note4[1] note4[2] note4[3] piano_keys[0]
+ piano_keys[10] piano_keys[11] piano_keys[12] piano_keys[13] piano_keys[14] piano_keys[1]
+ piano_keys[2] piano_keys[3] piano_keys[4] piano_keys[5] piano_keys[6] piano_keys[7]
+ piano_keys[8] piano_keys[9] pwm_o seq_led_on seq_play seq_power tempo_select vccd1
+ vssd1
X_7963_ net130 _0126_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6914_ _3184_ _3186_ vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7894_ net114 inputcont.INTERNAL_SYNCED_I\[1\] net75 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6845_ sound2.divisor_m\[2\] _1469_ _2864_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3988_ pm.count\[1\] pm.count\[0\] pm.count\[2\] vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__and3_1
X_6776_ sound1.sdiv.Q\[3\] _2895_ sound1.sdiv.next_dived sound1.sdiv.Q\[2\] vssd1
+ vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5727_ sound4.sdiv.Q\[15\] _2182_ _2185_ sound4.sdiv.Q\[14\] _2194_ vssd1 vssd1 vccd1
+ vccd1 _0015_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5658_ sound4.sdiv.A\[12\] _2062_ _2069_ _2140_ _2067_ vssd1 vssd1 vccd1 vccd1 _2141_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4609_ _0983_ _0978_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5589_ sound4.divisor_m\[11\] _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7328_ _3486_ _3490_ _3497_ vssd1 vssd1 vccd1 vccd1 _3498_ sky130_fd_sc_hd__nand3_1
XFILLER_0_102_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7259_ _2843_ _1618_ _3436_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__o21ai_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4960_ _1470_ _1506_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4891_ sound2.count\[4\] _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__xor2_1
X_3911_ _0575_ net66 vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__nor2_8
X_6630_ sound1.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ _0478_ _0485_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6561_ _2927_ _2929_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5512_ _0550_ _2001_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[2\] sky130_fd_sc_hd__nor2_1
X_3773_ inputcont.INTERNAL_SYNCED_I\[5\] vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
X_8300_ net122 _0400_ net83 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6492_ sound1.divisor_m\[10\] _2875_ _2864_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8231_ net129 sound3.osc.next_count\[12\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_5443_ _1779_ _1936_ _1948_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8162_ net140 _0283_ net101 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[15\] sky130_fd_sc_hd__dfrtp_1
X_5374_ sound4.count\[6\] _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7113_ sound2.sdiv.A\[24\] _3168_ sound2.sdiv.next_dived _3364_ vssd1 vssd1 vccd1
+ vccd1 _0231_ sky130_fd_sc_hd__a22o_1
X_4325_ _0894_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nand2_1
Xfanout105 net106 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_8
Xfanout127 net134 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_4
Xfanout138 net145 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
XFILLER_0_10_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout116 net119 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_4
X_8093_ net117 _0235_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[1\] sky130_fd_sc_hd__dfrtp_1
X_7044_ _3302_ _3303_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__or2_1
X_4256_ _0838_ _0813_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__and3b_1
X_4187_ seq.tempo_select.state\[1\] seq.clk_div.count\[12\] _0779_ seq.clk_div.count\[6\]
+ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7946_ net128 _0109_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7877_ net111 seq.encode.inter_keys\[10\] net72 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_sync\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6828_ sound2.count_m\[13\] _2857_ _3128_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6759_ sound1.sdiv.C\[1\] sound1.sdiv.C\[0\] sound1.sdiv.C\[2\] vssd1 vssd1 vccd1
+ vccd1 _3105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5090_ _1584_ _1595_ _1602_ _1620_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__or4_1
X_4110_ seq.player_6.state\[0\] _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__and2_1
X_4041_ _0675_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__buf_12
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5992_ _2402_ _2427_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7800_ net113 oct.next_state\[1\] net74 vssd1 vssd1 vccd1 vccd1 oct.state\[1\] sky130_fd_sc_hd__dfstp_1
X_7731_ net120 _0016_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[16\] sky130_fd_sc_hd__dfrtp_1
X_4943_ _1004_ _1321_ _1338_ _1158_ _1493_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7662_ _3722_ _2156_ vssd1 vssd1 vccd1 vccd1 _3723_ sky130_fd_sc_hd__xor2_1
X_6613_ _2903_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__and2_1
X_4874_ _0683_ _1323_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__or2_1
X_3825_ _0485_ _0501_ _0492_ _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__a211o_1
X_7593_ _3675_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_1
X_6544_ _2909_ _2915_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__or2_1
X_6475_ sound1.divisor_m\[3\] _2005_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8214_ net145 _0335_ net106 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5426_ sound4.count\[0\] _1779_ _1936_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[0\]
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_112_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8145_ net117 _0266_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[26\] sky130_fd_sc_hd__dfrtp_1
X_5357_ sound4.count\[4\] _1866_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__or2_1
X_8076_ net116 _0218_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[11\] sky130_fd_sc_hd__dfrtp_1
X_4308_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__nor3b_1
X_5288_ _1773_ _1775_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__or2_1
X_4239_ seq.clk_div.count\[8\] _0824_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__nand2_1
X_7027_ _3277_ _3280_ _3288_ vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7929_ net129 _0092_ net90 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_123_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _0680_ _0958_ _1154_ _0950_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ sound1.sdiv.Q\[5\] _0579_ _2690_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5211_ sound3.count\[6\] _1732_ _1721_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__o21ai_1
X_6191_ sound2.sdiv.Q\[0\] sound2.sdiv.Q\[1\] sound2.sdiv.Q\[2\] _0578_ _2499_ vssd1
+ vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__o311a_1
X_5142_ _0948_ _1578_ _1617_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__o211a_2
XFILLER_0_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5073_ _1018_ _1556_ _1603_ _0971_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__a22o_1
X_4024_ _0581_ _0583_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5975_ _2409_ sound1.divisor_m\[4\] _2410_ sound1.divisor_m\[3\] vssd1 vssd1 vccd1
+ vccd1 _2411_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7714_ _3756_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4926_ _0993_ _1383_ _1471_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4857_ _0685_ _1323_ _1338_ _1165_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7645_ _2069_ _2140_ vssd1 vssd1 vccd1 vccd1 _3711_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3808_ _0473_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nand2_1
X_7576_ _3665_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6527_ _2897_ sound1.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__and2b_1
X_4788_ net39 _1316_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__nand2_8
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6458_ sound1.count_m\[16\] _2836_ _2854_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6389_ pm.current_waveform\[2\] _2812_ _2808_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5409_ net63 _1784_ _1781_ _1038_ _1769_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__o221a_1
X_8128_ net120 _0249_ net81 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8059_ net116 _0201_ net77 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5760_ _2207_ _2212_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4711_ sound1.count\[7\] _1272_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_1
X_5691_ _2169_ _2170_ _2171_ _2172_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7430_ _3586_ _3588_ vssd1 vssd1 vccd1 vccd1 _3589_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4642_ _0695_ _0977_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__or2_4
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7361_ _3448_ _3526_ vssd1 vssd1 vccd1 vccd1 _3527_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4573_ _1136_ _1137_ _1143_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7292_ sound3.divisor_m\[3\] sound3.divisor_m\[2\] sound3.divisor_m\[1\] sound3.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3465_ sky130_fd_sc_hd__or4_1
X_6312_ _2740_ _2742_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6243_ _2672_ _2675_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6174_ _2374_ _2574_ _2608_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__a21o_1
X_5125_ _1642_ _1649_ _1655_ sound3.count\[2\] vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5056_ _0677_ _1574_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__or2_1
X_4007_ wave.mode\[0\] inputcont.INTERNAL_MODE _0658_ vssd1 vssd1 vccd1 vccd1 _0659_
+ sky130_fd_sc_hd__and3_1
X_5958_ _2377_ _2380_ _2388_ _2393_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__and4bb_1
X_4909_ sound2.count\[16\] _1459_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5889_ sound4.count_m\[13\] _2142_ sound4.divisor_m\[13\] _2324_ vssd1 vssd1 vccd1
+ vccd1 _2325_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7628_ _2132_ _3697_ vssd1 vssd1 vccd1 vccd1 _3699_ sky130_fd_sc_hd__or2b_1
XFILLER_0_105_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7559_ _3655_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 inputcont.u1.ff_intermediate\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6930_ _1311_ _3201_ vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__nand2_1
X_6861_ sound2.divisor_m\[8\] _3147_ _3142_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5812_ _2256_ _2257_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6792_ sound1.sdiv.Q\[19\] _2893_ _0867_ sound1.sdiv.Q\[18\] _2849_ vssd1 vssd1 vccd1
+ vccd1 _0160_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5743_ sound4.count\[15\] _2201_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5674_ _2154_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__nor2_1
X_7413_ _3570_ _3572_ vssd1 vssd1 vccd1 vccd1 _3574_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4625_ _0959_ _1082_ _1192_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7344_ _3510_ _3511_ _3503_ _3507_ vssd1 vssd1 vccd1 vccd1 _3512_ sky130_fd_sc_hd__o211ai_1
X_4556_ _1025_ _1038_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nor2_4
XFILLER_0_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7275_ sound3.divisor_m\[2\] _3449_ vssd1 vssd1 vccd1 vccd1 _3450_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4487_ _0685_ _0977_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6226_ sound1.sdiv.Q\[5\] _2293_ _2658_ _2292_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__o2bb2a_1
X_6157_ sound2.sdiv.Q\[2\] _0578_ _2591_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__and3_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _1189_ _1565_ _1637_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__o211a_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ sound3.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__inv_2
X_5039_ _1569_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 mode_out[1] sky130_fd_sc_hd__buf_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 note2[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5390_ _0973_ _1777_ _1800_ _1016_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4341_ seq.player_5.state\[0\] _0890_ _0892_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4272_ _0850_ _0813_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__and3b_1
X_7060_ sound2.divisor_m\[17\] _3308_ _3177_ vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6011_ sound2.count_m\[15\] _2446_ sound2.count_m\[14\] _2440_ vssd1 vssd1 vccd1
+ vccd1 _2447_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7962_ net130 _0125_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6913_ sound2.divisor_m\[3\] _3185_ vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7893_ net114 inputcont.INTERNAL_SYNCED_I\[0\] net75 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6844_ _3137_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3987_ pm.count\[1\] pm.count\[0\] vssd1 vssd1 vccd1 vccd1 pm.next_count\[1\] sky130_fd_sc_hd__xor2_1
X_6775_ _2435_ _0866_ _2588_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5726_ sound4.count\[7\] _2186_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5657_ _2073_ _2138_ _2139_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__a21o_1
X_4608_ _0943_ _1028_ _1175_ _0976_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5588_ sound4.divisor_m\[10\] _2030_ _2036_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7327_ _3495_ _3496_ vssd1 vssd1 vccd1 vccd1 _3497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4539_ _0944_ _1012_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7258_ _2543_ _2005_ vssd1 vssd1 vccd1 vccd1 _3436_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6209_ _2640_ _2642_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__xor2_1
X_7189_ sound3.count_m\[8\] _3132_ _3395_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__a21o_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3910_ _0577_ vssd1 vssd1 vccd1 vccd1 sound3.sdiv.next_start sky130_fd_sc_hd__inv_2
X_4890_ _1139_ _1327_ _1435_ _1440_ _1317_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3841_ _0500_ _0491_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__nor2_2
XFILLER_0_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6560_ _2927_ _2929_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__or2_1
X_3772_ inputcont.INTERNAL_SYNCED_I\[9\] inputcont.INTERNAL_SYNCED_I\[10\] _0454_
+ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5511_ rate_clk.count\[1\] rate_clk.count\[0\] rate_clk.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _2001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6491_ _1157_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8230_ net129 sound3.osc.next_count\[11\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_5442_ sound4.count\[4\] _1944_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8161_ net132 _0282_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[14\] sky130_fd_sc_hd__dfrtp_1
X_5373_ _1880_ _1883_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7112_ _3360_ _3363_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__xor2_1
X_8092_ net117 _0234_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[0\] sky130_fd_sc_hd__dfrtp_1
X_4324_ seq.player_6.state\[0\] seq.player_6.state\[1\] seq.player_6.state\[2\] seq.player_6.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__or4_1
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout106 net3 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_8
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_4
X_7043_ _3299_ _3301_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__and2_1
Xfanout117 net119 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_4
Xfanout139 net145 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_4
XFILLER_0_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4255_ seq.clk_div.count\[12\] _0835_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4186_ seq.clk_div.count\[10\] vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__inv_2
X_7945_ net128 _0108_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7876_ net113 inputcont.u1.ff_intermediate\[7\] net74 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_6827_ sound2.count\[13\] _2855_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6758_ _2890_ _3103_ _3104_ _2894_ sound1.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 _0136_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6689_ sound1.divisor_m\[17\] _3036_ _2903_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__o21a_1
X_5709_ _0576_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__buf_6
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8359_ net136 sound4.osc.next_count\[17\] net97 vssd1 vssd1 vccd1 vccd1 sound4.count\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _0676_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__nor2_8
XFILLER_0_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5991_ _2400_ _2401_ _2397_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4942_ _1129_ _1347_ _1343_ _1014_ _1427_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__o221a_1
X_7730_ net120 _0015_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7661_ _2053_ _3720_ vssd1 vssd1 vccd1 vccd1 _3722_ sky130_fd_sc_hd__and2b_1
X_6612_ sound1.divisor_m\[9\] sound1.divisor_m\[8\] sound1.divisor_m\[7\] _2948_ vssd1
+ vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__or4_1
X_4873_ sound2.count\[14\] _1422_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3824_ _0481_ _0482_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nand2_2
X_7592_ sound4.divisor_m\[14\] _3674_ _2186_ vssd1 vssd1 vccd1 vccd1 _3675_ sky130_fd_sc_hd__mux2_1
X_6543_ _2913_ _2914_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6474_ _2865_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8213_ net145 _0334_ net106 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5425_ _1935_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8144_ net117 _0265_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[25\] sky130_fd_sc_hd__dfrtp_1
X_5356_ sound4.count\[4\] _1866_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__nand2_1
X_4307_ _0876_ _0877_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__nand2_1
X_5287_ _1146_ _1777_ _1792_ _1134_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__o221a_1
X_8075_ net116 _0217_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[10\] sky130_fd_sc_hd__dfrtp_1
X_4238_ seq.clk_div.count\[8\] _0824_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__or2_1
X_7026_ _3286_ _3287_ vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4169_ seq.encode.keys_edge_det\[2\] inputcont.INTERNAL_SYNCED_I\[0\] vssd1 vssd1
+ vccd1 vccd1 _0769_ sky130_fd_sc_hd__and2b_1
X_7928_ net128 _0091_ net89 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7859_ net107 seq.clk_div.next_count\[16\] net68 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5210_ sound3.count\[6\] _1732_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6190_ sound2.sdiv.Q\[4\] _0578_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__nand2_1
X_5141_ _1001_ _1570_ _1668_ _1671_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__o211a_1
X_5072_ _1556_ _1557_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ _0588_ _0584_ _0585_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__or3b_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5974_ sound1.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__inv_2
X_7713_ wave_comb.u1.M\[2\] net34 _0645_ vssd1 vssd1 vccd1 vccd1 _3756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4925_ _1095_ _1343_ _1472_ _1473_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4856_ _1126_ _1347_ _1341_ _1166_ _1406_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__o221a_1
X_7644_ _2069_ _2140_ vssd1 vssd1 vccd1 vccd1 _3710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3807_ _0477_ _0478_ _0479_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__and4b_1
X_7575_ sound4.divisor_m\[7\] _3664_ _3419_ vssd1 vssd1 vccd1 vccd1 _3665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6526_ sound1.sdiv.A\[1\] _2895_ sound1.sdiv.next_dived _2899_ vssd1 vssd1 vccd1
+ vccd1 _0109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4787_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__buf_4
X_6457_ sound1.count\[16\] _2201_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6388_ _2439_ _2581_ _2805_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__mux2_1
X_5408_ _0954_ _1777_ _1792_ _0985_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8127_ net120 _0248_ net81 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[8\] sky130_fd_sc_hd__dfrtp_2
X_5339_ _1844_ _1845_ _1849_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__or3_2
X_8058_ net109 _0200_ net70 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[12\] sky130_fd_sc_hd__dfrtp_1
X_7009_ _3164_ _3271_ _3272_ _3174_ sound2.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _0219_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _1274_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_5690_ sound4.sdiv.A\[23\] _2038_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__and2_2
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4641_ _1210_ _0869_ _0965_ _1011_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7360_ sound3.divisor_m\[10\] _3515_ vssd1 vssd1 vccd1 vccd1 _3526_ sky130_fd_sc_hd__or2_1
X_4572_ _0981_ _1138_ _1139_ _0969_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7291_ sound3.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _3464_ sky130_fd_sc_hd__inv_2
X_6311_ _2703_ _2707_ _2741_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6242_ sound4.sdiv.Q\[5\] _2290_ _2674_ _2292_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6173_ _2507_ _2573_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__and2_1
X_5124_ _1005_ _1578_ _1550_ _1017_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__o221a_2
X_5055_ _1057_ _1567_ _1565_ _1056_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__o221a_1
X_4006_ inputcont.u3.next_in vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _2389_ _2390_ _2391_ _2392_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__and4b_1
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4908_ _1010_ _1456_ _1458_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7627_ _3697_ _2132_ vssd1 vssd1 vccd1 vccd1 _3698_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5888_ sound4.count_m\[12\] vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4839_ _0954_ _1347_ _1345_ _1182_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7558_ sound4.divisor_m\[0\] _1859_ _3419_ vssd1 vssd1 vccd1 vccd1 _3655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7489_ _3437_ _3637_ _3639_ _3440_ sound3.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _0332_
+ sky130_fd_sc_hd__a32o_1
X_6509_ sound1.divisor_m\[16\] _2886_ _2864_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 inputcont.u1.ff_intermediate\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6860_ _1412_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__inv_2
X_5811_ _2248_ _2252_ _2247_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__a21boi_1
X_6791_ sound1.sdiv.Q\[18\] _2893_ _0867_ sound1.sdiv.Q\[17\] _2848_ vssd1 vssd1 vccd1
+ vccd1 _0159_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5742_ sound4.sdiv.Q\[22\] _2182_ _2185_ sound4.sdiv.Q\[21\] _2202_ vssd1 vssd1 vccd1
+ vccd1 _0022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5673_ _2155_ _2049_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7412_ _3570_ _3572_ vssd1 vssd1 vccd1 vccd1 _3573_ sky130_fd_sc_hd__nor2_1
X_4624_ _1193_ _0967_ _0943_ _1158_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7343_ sound3.sdiv.A\[8\] _3509_ vssd1 vssd1 vccd1 vccd1 _3511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4555_ _0959_ net63 vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7274_ sound3.divisor_m\[1\] sound3.divisor_m\[0\] _3448_ vssd1 vssd1 vccd1 vccd1
+ _3449_ sky130_fd_sc_hd__o21a_1
X_4486_ _0695_ _0970_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6225_ _2620_ _2657_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6156_ sound2.sdiv.Q\[0\] sound2.sdiv.Q\[1\] _0578_ _2499_ vssd1 vssd1 vccd1 vccd1
+ _2591_ sky130_fd_sc_hd__o211a_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _1204_ _1553_ _1580_ _1199_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__o22a_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _2521_ sound3.divisor_m\[14\] sound3.divisor_m\[13\] _2522_ vssd1 vssd1 vccd1
+ vccd1 _2523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5038_ _1563_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6989_ _3164_ _3253_ _3254_ _3174_ sound2.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _0217_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 multi[0] sky130_fd_sc_hd__clkbuf_4
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 note3[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4340_ seq.player_6.state\[0\] _0894_ _0896_ _0910_ vssd1 vssd1 vccd1 vccd1 _0911_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4271_ seq.clk_div.count\[16\] _0847_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6010_ sound2.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7961_ net130 _0124_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[16\] sky130_fd_sc_hd__dfrtp_1
X_7892_ net113 seq.encode.keys_sync\[1\] net74 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6912_ sound2.divisor_m\[2\] sound2.divisor_m\[1\] sound2.divisor_m\[0\] _3177_ vssd1
+ vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6843_ sound2.divisor_m\[1\] _3136_ _2864_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3986_ pm.count\[0\] vssd1 vssd1 vccd1 vccd1 pm.next_count\[0\] sky130_fd_sc_hd__inv_2
X_6774_ sound1.sdiv.Q\[0\] sound1.sdiv.next_dived _2436_ vssd1 vssd1 vccd1 vccd1 _0142_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5725_ sound4.sdiv.Q\[14\] _2182_ _2185_ sound4.sdiv.Q\[13\] _2193_ vssd1 vssd1 vccd1
+ vccd1 _0014_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5656_ _2070_ _2072_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4607_ _0954_ _0994_ _0992_ _1129_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5587_ sound4.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7326_ _3491_ _3494_ vssd1 vssd1 vccd1 vccd1 _3496_ sky130_fd_sc_hd__nand2_1
X_4538_ _0677_ _1084_ _1090_ _0952_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o22a_1
X_7257_ _3435_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
X_4469_ _0674_ _0977_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__nor2_4
X_6208_ sound4.sdiv.Q\[2\] _2641_ _2582_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__a21o_1
X_7188_ sound3.count\[8\] _2863_ vssd1 vssd1 vccd1 vccd1 _3395_ sky130_fd_sc_hd__and2_1
X_6139_ _2374_ _2574_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3840_ inputcont.INTERNAL_SYNCED_I\[3\] _0502_ _0512_ _0513_ vssd1 vssd1 vccd1 vccd1
+ _0514_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3771_ inputcont.INTERNAL_SYNCED_I\[8\] _0443_ _0444_ vssd1 vssd1 vccd1 vccd1 _0454_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5510_ rate_clk.count\[1\] rate_clk.count\[0\] vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6490_ _2005_ _1196_ _2874_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ sound4.count\[4\] _1944_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__nand2_1
X_8160_ net132 _0281_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[13\] sky130_fd_sc_hd__dfrtp_1
X_5372_ _0679_ net63 _1784_ _1882_ _1778_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__o311a_1
XFILLER_0_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7111_ _3343_ _3361_ _3362_ _3352_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__o211a_1
X_8091_ net117 _0233_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4323_ select1.sequencer_on _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__and2_1
Xfanout129 net134 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_8
X_7042_ _3299_ _3301_ vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__nor2_1
Xfanout107 net115 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_4
X_4254_ seq.clk_div.count\[12\] _0835_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4185_ seq.clk_div.count\[18\] vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__inv_2
X_7944_ net125 _0107_ net86 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ net110 inputcont.u1.ff_intermediate\[6\] net71 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6826_ sound2.count_m\[12\] _2857_ _3127_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__a21o_1
X_6757_ sound1.sdiv.C\[1\] sound1.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3969_ net34 _0632_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__nor2_2
X_5708_ sound4.sdiv.Q\[7\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[6\] vssd1
+ vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6688_ sound1.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5639_ sound4.divisor_m\[1\] _2121_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8358_ net136 sound4.osc.next_count\[16\] net97 vssd1 vssd1 vccd1 vccd1 sound4.count\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7309_ _3468_ _3471_ _3479_ vssd1 vssd1 vccd1 vccd1 _3481_ sky130_fd_sc_hd__or3b_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8289_ net121 _0389_ net82 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5990_ _2382_ _2425_ _2389_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__a21o_1
X_4941_ _1020_ _1333_ _1345_ _1083_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__o221a_1
X_4872_ sound2.count\[14\] _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7660_ _3681_ _3720_ _3721_ _2184_ sound4.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 _0421_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6611_ _2962_ _2963_ _2975_ _2966_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3823_ _0479_ _0478_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7591_ _1817_ vssd1 vssd1 vccd1 vccd1 _3674_ sky130_fd_sc_hd__inv_2
X_6542_ _2910_ _2912_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6473_ sound1.divisor_m\[2\] _2862_ _2864_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8212_ net142 _0333_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5424_ _1861_ _1886_ _1934_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8143_ net117 _0264_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5355_ _0696_ _1792_ _1794_ _1140_ _1865_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4306_ seq.player_2.state\[0\] seq.player_2.state\[1\] seq.player_2.state\[2\] seq.player_2.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__or4_1
X_5286_ _1154_ _1794_ _1796_ _1042_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__o22a_1
X_8074_ net116 _0216_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[9\] sky130_fd_sc_hd__dfrtp_1
X_4237_ _0824_ _0825_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[7\] sky130_fd_sc_hd__nor2_1
X_7025_ _3282_ _3285_ vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__nand2_1
X_4168_ _0766_ _0765_ _0768_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_2.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4099_ seq.player_7.state\[1\] seq.player_7.state\[2\] seq.player_7.state\[3\] _0722_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__a311o_1
X_7927_ net129 _0090_ net90 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[1\] sky130_fd_sc_hd__dfrtp_4
X_7858_ net108 seq.clk_div.next_count\[15\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6809_ sound2.count\[4\] _2855_ vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__and2_1
X_7789_ net107 inputcont.u1.ff_intermediate\[11\] net68 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_61_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5140_ _0973_ _1553_ _1574_ _0979_ _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5071_ sound3.count\[4\] _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__xnor2_1
X_4022_ _0594_ _0669_ _0596_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5973_ sound1.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7712_ _3755_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4924_ _1041_ _1323_ _1327_ _1096_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4855_ _1159_ _1343_ _1333_ _0997_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7643_ _3681_ _3708_ _3709_ _2184_ sound4.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _0416_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4786_ net39 _1325_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__or2_1
X_3806_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__buf_2
X_7574_ _1897_ vssd1 vssd1 vccd1 vccd1 _3664_ sky130_fd_sc_hd__inv_2
X_6525_ _2891_ _2898_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6456_ sound1.count_m\[15\] _2836_ _2853_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6387_ _2811_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
X_5407_ _1912_ _1914_ _1917_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__or3b_1
X_8126_ net136 _0247_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[7\] sky130_fd_sc_hd__dfrtp_4
X_5338_ _1125_ _1796_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__o21ai_1
X_8057_ net116 _0199_ net77 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[11\] sky130_fd_sc_hd__dfrtp_2
X_7008_ _3259_ _3262_ _3270_ vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__o21bai_1
X_5269_ net47 _1770_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4640_ _0909_ _0937_ _1138_ _0974_ _0688_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__o32a_1
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6310_ _2698_ _2702_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__and2_1
X_4571_ _1000_ _1140_ _1141_ _0976_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__o22a_1
X_7290_ _3461_ _3462_ sound3.sdiv.A\[3\] _3463_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6241_ _2639_ _2673_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6172_ _2585_ _2606_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5123_ _1025_ _1028_ _1553_ _1650_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__o311a_1
X_5054_ _0959_ _1133_ _1553_ _1578_ _0983_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__o32a_1
X_4005_ pm.count\[7\] _0655_ pm.count\[8\] vssd1 vssd1 vccd1 vccd1 pm.next_count\[8\]
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ sound1.divisor_m\[9\] sound1.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5887_ _2322_ sound4.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__or2_1
X_4907_ _0688_ _1418_ _1317_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__o211a_1
X_4838_ _1129_ _1341_ _1336_ _1175_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7626_ _2133_ _2093_ vssd1 vssd1 vccd1 vccd1 _3697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7557_ sound4.count_m\[18\] _2843_ _2206_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__a21o_1
X_4769_ _0499_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7488_ _3622_ _3631_ _3638_ _3636_ vssd1 vssd1 vccd1 vccd1 _3639_ sky130_fd_sc_hd__a31o_1
X_6508_ _1219_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6439_ _1073_ _2843_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8109_ net110 sound2.osc.next_count\[10\] net71 vssd1 vssd1 vccd1 vccd1 sound2.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 inputcont.u1.ff_intermediate\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5810_ _2254_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__nand2_1
X_6790_ sound1.sdiv.Q\[17\] _2893_ _0867_ sound1.sdiv.Q\[16\] _2847_ vssd1 vssd1 vccd1
+ vccd1 _0158_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ sound4.count\[14\] _2201_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7411_ sound3.divisor_m\[16\] _3571_ vssd1 vssd1 vccd1 vccd1 _3572_ sky130_fd_sc_hd__xnor2_1
X_5672_ _2046_ _2048_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4623_ _0992_ _1028_ _1020_ _0990_ _1130_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7342_ sound3.sdiv.A\[8\] _3509_ vssd1 vssd1 vccd1 vccd1 _3510_ sky130_fd_sc_hd__and2_1
X_4554_ _1124_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7273_ sound3.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _3448_ sky130_fd_sc_hd__inv_4
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6224_ sound1.sdiv.Q\[3\] _2656_ _2621_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__a21oi_1
X_4485_ _0678_ _1055_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6155_ _2279_ _2586_ _2589_ _2289_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__a2bb2o_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ sound3.count_m\[12\] vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__inv_2
X_5106_ _1200_ _1567_ _1550_ _0686_ _1636_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__o221a_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ net46 _1555_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6988_ _3233_ _3237_ _3251_ _3241_ _3250_ vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__a311o_1
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5939_ sound1.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7609_ _2120_ _2125_ vssd1 vssd1 vccd1 vccd1 _3685_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 beat_led[0] sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 multi[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 note3[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4270_ seq.clk_div.count\[16\] _0847_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7960_ net130 _0123_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6911_ sound2.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__inv_2
X_7891_ net114 seq.encode.keys_sync\[0\] net75 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6842_ _1404_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6773_ _0866_ _3114_ _2277_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__o21ai_1
X_3985_ _0646_ vssd1 vssd1 vccd1 vccd1 wave_comb.u1.next_dived sky130_fd_sc_hd__buf_4
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5724_ sound4.count\[6\] _2186_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5655_ _2079_ _2137_ _2077_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4606_ _0950_ _0996_ _1176_ _0981_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7325_ _3491_ _3494_ vssd1 vssd1 vccd1 vccd1 _3495_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5586_ _2067_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__nor2_1
X_4537_ _0683_ _0981_ _0992_ _1052_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7256_ sound3.divisor_m\[17\] _1604_ _3419_ vssd1 vssd1 vccd1 vccd1 _3435_ sky130_fd_sc_hd__mux2_1
X_4468_ _1019_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__or2_4
X_7187_ sound3.count_m\[7\] _3132_ _3394_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__a21o_1
X_6207_ _0576_ _2370_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and2_1
X_6138_ _2507_ _2573_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__xor2_1
X_4399_ _0686_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__nand2_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _2439_ _2504_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__xnor2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3770_ _0441_ _0445_ _0447_ _0452_ _0453_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__o2111ai_4
XFILLER_0_104_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5440_ _1947_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5371_ _1057_ _1792_ _1794_ _1063_ _1881_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7110_ sound2.sdiv.A\[22\] sound2.sdiv.A\[21\] _3329_ vssd1 vssd1 vccd1 vccd1 _3362_
+ sky130_fd_sc_hd__o21ai_1
X_8090_ net118 _0232_ net79 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[25\] sky130_fd_sc_hd__dfrtp_1
X_4322_ seq.beat\[3\] seq.encode.play _0874_ inputcont.INTERNAL_SYNCED_I\[5\] vssd1
+ vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__a31o_1
Xfanout119 net2 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_4
X_7041_ sound2.divisor_m\[16\] _3300_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__xnor2_1
Xfanout108 net115 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_4
X_4253_ _0837_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
X_4184_ _0777_ _0778_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[1\] sky130_fd_sc_hd__nor2_1
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7943_ net125 _0106_ net86 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7874_ net108 inputcont.u1.ff_intermediate\[5\] net69 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6825_ sound2.count\[12\] _2855_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__and2_1
X_6756_ sound1.sdiv.C\[1\] sound1.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3968_ _0630_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__or2_4
X_5707_ sound4.sdiv.Q\[6\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[5\] vssd1
+ vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a22o_1
X_6687_ sound1.sdiv.A\[17\] _2895_ sound1.sdiv.next_dived _3044_ vssd1 vssd1 vccd1
+ vccd1 _0125_ sky130_fd_sc_hd__a22o_1
X_3899_ _0554_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nand2_8
XFILLER_0_72_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5638_ sound4.sdiv.A\[26\] sound4.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8357_ net121 sound4.osc.next_count\[15\] net82 vssd1 vssd1 vccd1 vccd1 sound4.count\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5569_ sound4.divisor_m\[16\] _2051_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7308_ _3468_ _3471_ _3479_ vssd1 vssd1 vccd1 vccd1 _3480_ sky130_fd_sc_hd__o21bai_2
X_8288_ net121 _0388_ net82 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[2\] sky130_fd_sc_hd__dfrtp_4
X_7239_ _3424_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4940_ _1028_ _1341_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4871_ _0695_ _1417_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6610_ _2969_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__inv_2
X_3822_ _0443_ _0444_ inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1 vccd1 vccd1 _0500_
+ sky130_fd_sc_hd__o21ai_4
X_7590_ _3673_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__clkbuf_1
X_6541_ _2910_ _2912_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6472_ _2863_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8211_ net142 _0332_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5423_ _1911_ _1918_ _1925_ _1933_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__or4b_1
X_5354_ _1138_ _1769_ _1778_ _1864_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8142_ net116 _0263_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4305_ select1.sequencer_on _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__and2_1
X_8073_ net116 _0215_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[8\] sky130_fd_sc_hd__dfrtp_1
X_5285_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__clkbuf_4
X_4236_ seq.clk_div.count\[7\] _0822_ _0813_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7024_ _3282_ _3285_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__or2_1
X_4167_ seq.player_2.state\[1\] seq.player_2.state\[2\] _0762_ seq.player_2.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4098_ seq.player_7.state\[0\] _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__and2_1
X_7926_ net128 _0089_ net89 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7857_ net108 seq.clk_div.next_count\[14\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6808_ sound2.count_m\[3\] _2857_ _3118_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7788_ net128 inputcont.u1.ff_intermediate\[10\] net89 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6739_ _0866_ _3089_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout90 net95 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_4
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _1135_ _1550_ _1570_ _1140_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__o221a_1
X_4021_ _0668_ _0602_ _0592_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5972_ _2407_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__inv_2
X_7711_ wave_comb.u1.M\[1\] net33 _0645_ vssd1 vssd1 vccd1 vccd1 _3755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4923_ _1347_ _1336_ _0960_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7642_ _2138_ _3707_ vssd1 vssd1 vccd1 vccd1 _3709_ sky130_fd_sc_hd__or2b_1
X_4854_ _0677_ _1336_ _1345_ _1077_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7573_ _3663_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3805_ _0480_ _0481_ _0482_ net67 vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and4_1
X_4785_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__buf_4
X_6524_ sound1.sdiv.A\[0\] _2897_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6455_ sound1.count\[15\] _2201_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__and2_1
X_6386_ pm.current_waveform\[1\] _2810_ _2808_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5406_ sound4.count\[17\] _1222_ _1913_ _1915_ _1916_ vssd1 vssd1 vccd1 vccd1 _1917_
+ sky130_fd_sc_hd__o311a_1
X_8125_ net136 _0246_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[6\] sky130_fd_sc_hd__dfrtp_2
X_5337_ _1199_ _1800_ _1846_ _1847_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5268_ _1778_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__buf_4
X_8056_ net109 _0198_ net70 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[10\] sky130_fd_sc_hd__dfrtp_2
X_7007_ _3259_ _3262_ _3270_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__or3b_1
X_4219_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__buf_4
X_5199_ _1727_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7909_ net128 _0072_ net89 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4570_ _1038_ _1034_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6240_ sound4.sdiv.Q\[3\] _2641_ _2642_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__a21o_1
X_6171_ _2600_ _2605_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5122_ _1011_ _1559_ _1572_ _1020_ _1652_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__o221a_1
X_5053_ sound3.count\[0\] _1583_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__xor2_1
X_4004_ _0657_ _0655_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[7\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5955_ sound1.count_m\[9\] sound1.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 _2391_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5886_ sound4.count_m\[16\] vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _1324_ _1333_ _1055_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7625_ _3695_ _3696_ sound4.sdiv.A\[6\] _2183_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4837_ sound2.count\[10\] _1387_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7556_ sound4.count_m\[17\] _2843_ _2205_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4768_ _0507_ _1312_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__nand2_1
X_7487_ _3630_ _3623_ _3627_ vssd1 vssd1 vccd1 vccd1 _3638_ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6507_ _2885_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
X_4699_ sound1.count\[4\] _1263_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__nand2_1
X_6438_ sound1.count_m\[6\] _2836_ _2844_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6369_ _2794_ _2796_ net53 vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__or3_1
X_8108_ net110 sound2.osc.next_count\[9\] net71 vssd1 vssd1 vccd1 vccd1 sound2.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_8039_ net109 _0181_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 inputcont.u1.ff_intermediate\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5740_ _0575_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7410_ sound3.divisor_m\[15\] _3561_ _3448_ vssd1 vssd1 vccd1 vccd1 _3571_ sky130_fd_sc_hd__o21a_1
X_5671_ _2053_ _2153_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4622_ _1107_ _1100_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__or2_2
XFILLER_0_130_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7341_ sound3.divisor_m\[9\] _3508_ vssd1 vssd1 vccd1 vccd1 _3509_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4553_ _0683_ _1034_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7272_ sound3.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _3447_ sky130_fd_sc_hd__inv_2
X_4484_ _0676_ _0695_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__or2_4
XFILLER_0_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6223_ _0579_ _2434_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6154_ _2587_ _2588_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ sound3.count_m\[13\] vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__inv_2
X_5105_ _0683_ _1107_ _1570_ _1562_ _1198_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__o32a_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6987_ _3250_ _3252_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__nand2_1
X_5938_ _2289_ _2372_ _2373_ _2290_ sound4.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2374_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5869_ _2291_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7608_ sound4.sdiv.A\[1\] _2183_ sound4.sdiv.next_dived _3684_ vssd1 vssd1 vccd1
+ vccd1 _0406_ sky130_fd_sc_hd__a22o_1
X_7539_ sound4.count_m\[0\] _3403_ _2187_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 multi[2] sky130_fd_sc_hd__buf_2
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 beat_led[1] sky130_fd_sc_hd__clkbuf_4
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 note3[2] sky130_fd_sc_hd__buf_2
XFILLER_0_101_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6910_ _3176_ _3179_ vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__or2_1
X_7890_ net114 seq.encode.next_play net75 vssd1 vssd1 vccd1 vccd1 seq.encode.play
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6841_ _3135_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6772_ _3098_ _3100_ _3113_ _3096_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3984_ _0645_ _0571_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5723_ sound4.sdiv.Q\[13\] _2182_ _2185_ sound4.sdiv.Q\[12\] _2192_ vssd1 vssd1 vccd1
+ vccd1 _0013_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5654_ _2083_ _2135_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_60_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4605_ _0996_ _1019_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7324_ sound3.divisor_m\[7\] _3493_ vssd1 vssd1 vccd1 vccd1 _3494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5585_ _2063_ _2065_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__and2_1
X_4536_ _0685_ _0684_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nor2_8
XFILLER_0_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7255_ _3434_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
X_4467_ _0676_ _0695_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__nor2_8
X_7186_ _1642_ _2843_ vssd1 vssd1 vccd1 vccd1 _3394_ sky130_fd_sc_hd__nor2_1
X_6206_ sound4.sdiv.Q\[3\] _0576_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__nand2_1
X_4398_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__buf_4
X_6137_ _2289_ _2571_ _2572_ _2301_ sound3.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2573_
+ sky130_fd_sc_hd__a32o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _2289_ _2502_ _2503_ _2295_ sound2.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2504_
+ sky130_fd_sc_hd__a32o_1
X_5019_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__buf_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5370_ _1056_ _1777_ _1800_ _1053_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ _0890_ _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nand2_1
Xfanout109 net110 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_4
X_7040_ sound2.divisor_m\[15\] sound2.divisor_m\[14\] _3283_ _3177_ vssd1 vssd1 vccd1
+ vccd1 _3300_ sky130_fd_sc_hd__o31a_1
X_4252_ _0835_ _0813_ _0836_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__and3b_1
X_4183_ seq.clk_div.count\[1\] seq.clk_div.count\[0\] _0719_ vssd1 vssd1 vccd1 vccd1
+ _0778_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7942_ net126 _0105_ net87 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[16\] sky130_fd_sc_hd__dfrtp_2
X_7873_ net107 inputcont.u1.ff_intermediate\[4\] net68 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6824_ sound2.count_m\[11\] _2857_ _3126_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__a21o_1
X_6755_ _3102_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3967_ _0607_ _0629_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__and2_1
X_5706_ sound4.sdiv.Q\[5\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[4\] vssd1
+ vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6686_ _3042_ _3043_ vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3898_ sound4.sdiv.dived _0557_ _0560_ sound2.sdiv.dived _0567_ vssd1 vssd1 vccd1
+ vccd1 _0568_ sky130_fd_sc_hd__a221o_2
XFILLER_0_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5637_ _2117_ _2119_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8356_ net120 sound4.osc.next_count\[14\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_5568_ _2036_ _2033_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__and2_1
X_7307_ _3477_ _3478_ vssd1 vssd1 vccd1 vccd1 _3479_ sky130_fd_sc_hd__nand2_1
X_4519_ _0967_ _1025_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__or2_1
X_8287_ net123 _0387_ net84 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7238_ sound3.divisor_m\[10\] _1690_ _3419_ vssd1 vssd1 vccd1 vccd1 _3424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5499_ _1779_ _1936_ _1992_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__and4_1
X_7169_ sound2.sdiv.Q\[25\] _3167_ _1311_ sound2.sdiv.Q\[24\] _3133_ vssd1 vssd1 vccd1
+ vccd1 _0265_ sky130_fd_sc_hd__a221o_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4870_ _1111_ _1325_ _1334_ _1058_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3821_ _0499_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkinv_4
XFILLER_0_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6540_ sound1.divisor_m\[3\] _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6471_ _0575_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__clkbuf_8
X_8210_ net144 _0331_ net105 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5422_ sound4.count\[1\] _1931_ _1909_ sound4.count\[11\] _1932_ vssd1 vssd1 vccd1
+ vccd1 _1933_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5353_ _1135_ _1784_ _1796_ _1141_ _1863_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__o221a_1
X_8141_ net109 _0262_ net70 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4304_ _0702_ seq.encode.play _0874_ inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1
+ vccd1 vccd1 _0875_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8072_ net116 _0214_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5284_ _1782_ _1771_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__or2_1
X_4235_ seq.clk_div.count\[6\] seq.clk_div.count\[7\] _0819_ vssd1 vssd1 vccd1 vccd1
+ _0824_ sky130_fd_sc_hd__and3_1
X_7023_ _2441_ _3284_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__xnor2_1
X_4166_ _0766_ _0765_ _0767_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_2.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4097_ seq.encode.keys_edge_det\[8\] inputcont.INTERNAL_SYNCED_I\[6\] vssd1 vssd1
+ vccd1 vccd1 _0721_ sky130_fd_sc_hd__and2b_1
X_7925_ net127 _0088_ net88 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7856_ net108 seq.clk_div.next_count\[13\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6807_ _1318_ _2843_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7787_ net113 inputcont.u1.ff_intermediate\[9\] net74 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_4999_ _1535_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_6738_ net55 _3087_ _3084_ _3085_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6669_ sound1.divisor_m\[15\] sound1.divisor_m\[14\] _3011_ vssd1 vssd1 vccd1 vccd1
+ _3028_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8339_ net138 _0439_ net99 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.M\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout91 net95 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_8
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout80 net3 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_8
XFILLER_0_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _0599_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5971_ sound1.count_m\[17\] _2405_ sound1.count_m\[16\] _2406_ vssd1 vssd1 vccd1
+ vccd1 _2407_ sky130_fd_sc_hd__o22a_1
X_7710_ _3754_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4922_ _1101_ _1333_ _1345_ _1097_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7641_ _3707_ _2138_ vssd1 vssd1 vccd1 vccd1 _3708_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4853_ _1398_ _1400_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7572_ sound4.divisor_m\[6\] _1884_ _3419_ vssd1 vssd1 vccd1 vccd1 _3663_ sky130_fd_sc_hd__mux2_1
X_3804_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[3\]
+ inputcont.INTERNAL_SYNCED_I\[2\] inputcont.INTERNAL_SYNCED_I\[4\] vssd1 vssd1 vccd1
+ vccd1 _0483_ sky130_fd_sc_hd__o41ai_1
X_4784_ _1330_ _1334_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__or2_1
X_6523_ sound1.divisor_m\[1\] _2896_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__xnor2_1
X_6454_ sound1.count_m\[14\] _2836_ _2852_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5405_ sound4.count\[18\] _1778_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6385_ _2294_ _2310_ _2805_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8124_ net136 _0245_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[5\] sky130_fd_sc_hd__dfrtp_2
X_5336_ _1198_ _1769_ _1777_ _1189_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__o22a_1
X_8055_ net109 _0197_ net70 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[9\] sky130_fd_sc_hd__dfrtp_2
X_5267_ _1772_ _1773_ _1777_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__nand3_4
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7006_ _3268_ _3269_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__nand2_1
X_4218_ _0719_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__and2_1
X_5198_ _1721_ _1725_ _1726_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4149_ seq.player_3.state\[0\] seq.player_3.state\[1\] _0753_ vssd1 vssd1 vccd1 vccd1
+ _0756_ sky130_fd_sc_hd__and3_1
X_7908_ net128 _0071_ net89 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7839_ net143 _0062_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6170_ sound3.sdiv.Q\[3\] _2301_ _2603_ _2604_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _0997_ _1562_ _1565_ _0973_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__o221a_1
X_5052_ _1554_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__nand2_1
X_4003_ pm.count\[7\] vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5954_ sound1.count_m\[8\] sound1.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5885_ _2313_ sound4.divisor_m\[4\] _2317_ _2319_ _2320_ vssd1 vssd1 vccd1 vccd1
+ _2321_ sky130_fd_sc_hd__a2111oi_1
X_4905_ _1450_ _1334_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7624_ _2099_ _2131_ _2185_ vssd1 vssd1 vccd1 vccd1 _3696_ sky130_fd_sc_hd__o21ai_1
X_4836_ _1107_ net63 _1322_ _1380_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__o311a_2
X_7555_ sound4.count_m\[16\] _2843_ _2204_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6506_ sound1.divisor_m\[15\] _2884_ _2864_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4767_ sound2.count\[3\] vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7486_ _3629_ _3630_ _3631_ _3636_ vssd1 vssd1 vccd1 vccd1 _3637_ sky130_fd_sc_hd__o211ai_1
X_4698_ _1265_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6437_ _1237_ _2843_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6368_ _2762_ _2791_ _2792_ _2793_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__nor4_1
X_8107_ net110 sound2.osc.next_count\[8\] net71 vssd1 vssd1 vccd1 vccd1 sound2.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_5319_ sound4.count\[8\] _1829_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__and2_1
X_6299_ _2728_ _2729_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__xnor2_2
X_8038_ net109 _0180_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 inputcont.u1.ff_intermediate\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5670_ _2050_ _2052_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4621_ _0939_ _1014_ _1188_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7340_ sound3.divisor_m\[8\] _3448_ _3501_ vssd1 vssd1 vccd1 vccd1 _3508_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4552_ _0679_ _0971_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7271_ _3442_ sound3.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _3446_ sky130_fd_sc_hd__or2b_1
X_4483_ _0679_ _0950_ _1040_ _1053_ _0992_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o32a_1
XFILLER_0_52_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6222_ wave_comb.u1.next_start _2654_ _2655_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__a21bo_1
X_6153_ sound1.sdiv.Q\[2\] _0579_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ sound3.divisor_m\[1\] _2517_ _2518_ _2519_ vssd1 vssd1 vccd1 vccd1 _2520_
+ sky130_fd_sc_hd__o211ai_1
X_5104_ _1181_ _1559_ _1578_ _1028_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__o221a_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _1560_ _1551_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__or2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6986_ _3233_ _3237_ _3251_ _3241_ vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5937_ sound4.sdiv.Q\[1\] _2181_ _2370_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5868_ _2303_ _2304_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__nor2_1
X_7607_ _2123_ _3682_ vssd1 vssd1 vccd1 vccd1 _3684_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5799_ wave_comb.u1.next_dived _2245_ _2246_ _0573_ wave_comb.u1.A\[7\] vssd1 vssd1
+ vccd1 vccd1 _0035_ sky130_fd_sc_hd__a32o_1
X_4819_ _1318_ _1352_ _1360_ sound2.count\[12\] _1369_ vssd1 vssd1 vccd1 vccd1 _1370_
+ sky130_fd_sc_hd__a221o_1
X_7538_ sound3.sdiv.Q\[27\] _3440_ _3437_ sound3.sdiv.Q\[26\] vssd1 vssd1 vccd1 vccd1
+ _0366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7469_ sound3.sdiv.A\[23\] _3595_ vssd1 vssd1 vccd1 vccd1 _3622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 beat_led[2] sky130_fd_sc_hd__clkbuf_4
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 note3[3] sky130_fd_sc_hd__buf_2
Xoutput35 net58 vssd1 vssd1 vccd1 vccd1 note1[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6840_ sound2.divisor_m\[0\] _1477_ _2864_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__mux2_1
X_6771_ sound1.divisor_m\[18\] sound1.divisor_m\[17\] sound1.sdiv.A\[26\] _3036_ vssd1
+ vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__or4_1
X_3983_ _0644_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__buf_4
X_5722_ sound4.count\[5\] _2186_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5653_ sound4.sdiv.A\[8\] _2082_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4604_ _1001_ _1028_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nor2_2
X_5584_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7323_ _3448_ _3492_ vssd1 vssd1 vccd1 vccd1 _3493_ sky130_fd_sc_hd__and2_1
X_4535_ sound1.count\[2\] _1032_ _1072_ sound1.count\[6\] _1105_ vssd1 vssd1 vccd1
+ vccd1 _1106_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7254_ sound3.divisor_m\[16\] _3433_ _3419_ vssd1 vssd1 vccd1 vccd1 _3434_ sky130_fd_sc_hd__mux2_1
X_4466_ _0992_ _1033_ _1035_ _0981_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__o221a_1
X_7185_ sound3.count_m\[6\] _3132_ _3393_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a21o_1
X_6205_ sound4.sdiv.Q\[4\] _0576_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4397_ _0918_ _0941_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__or2_1
X_6136_ _2570_ _2275_ sound3.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6067_ _2500_ _2276_ _2499_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__or3b_1
X_5018_ _0540_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__or2_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6969_ _3224_ _3228_ _3235_ vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4320_ seq.player_5.state\[0\] seq.player_5.state\[1\] seq.player_5.state\[2\] seq.player_5.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__or4_1
X_4251_ seq.clk_div.count\[11\] _0832_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4182_ seq.clk_div.count\[1\] seq.clk_div.count\[0\] vssd1 vssd1 vccd1 vccd1 _0777_
+ sky130_fd_sc_hd__and2_1
X_7941_ net126 _0104_ net87 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7872_ net111 inputcont.u1.ff_intermediate\[3\] net72 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6823_ sound2.count\[11\] _2855_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__and2_1
X_6754_ _0867_ _2893_ sound1.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3966_ _0607_ _0629_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__nor2_2
X_6685_ _3031_ _3035_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__nand2_1
X_5705_ sound4.sdiv.Q\[4\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[3\] vssd1
+ vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3897_ sound3.sdiv.dived _0563_ _0566_ sound1.sdiv.dived vssd1 vssd1 vccd1 vccd1
+ _0567_ sky130_fd_sc_hd__a22o_1
X_5636_ sound4.divisor_m\[2\] _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__xnor2_1
X_8355_ net120 sound4.osc.next_count\[13\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5567_ sound4.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__inv_2
X_7306_ _3474_ _3476_ vssd1 vssd1 vccd1 vccd1 _3478_ sky130_fd_sc_hd__nand2_1
X_4518_ _1075_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__nand2_1
X_5498_ sound4.count\[16\] _1988_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__or2_1
X_8286_ net121 _0386_ net82 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[0\] sky130_fd_sc_hd__dfrtp_4
X_7237_ _3423_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__clkbuf_1
X_4449_ _1018_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__or2_4
XFILLER_0_0_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7168_ sound2.sdiv.Q\[24\] _3167_ _1311_ sound2.sdiv.Q\[23\] _3131_ vssd1 vssd1 vccd1
+ vccd1 _0264_ sky130_fd_sc_hd__a221o_1
X_6119_ _2551_ sound3.count_m\[0\] _2552_ _2553_ _2554_ vssd1 vssd1 vccd1 vccd1 _2555_
+ sky130_fd_sc_hd__o2111a_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _3350_ _3351_ _3352_ vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__nand3_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3820_ _0472_ _0487_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__o21ba_4
XFILLER_0_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6470_ _1032_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5421_ sound4.count\[1\] _1931_ _1891_ sound4.count\[15\] vssd1 vssd1 vccd1 vccd1
+ _1932_ sky130_fd_sc_hd__o2bb2a_1
X_5352_ _1127_ _1777_ _1800_ _1126_ _1862_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8140_ net109 _0261_ net70 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8071_ net116 _0213_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[6\] sky130_fd_sc_hd__dfrtp_1
X_4303_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__nor3b_1
X_7022_ _3177_ _3283_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__nand2_1
X_5283_ _1793_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4234_ _0822_ _0823_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[6\] sky130_fd_sc_hd__nor2_1
X_4165_ seq.player_2.state\[2\] _0764_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4096_ _0717_ _0716_ _0720_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_8.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_7924_ net127 _0087_ net88 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[17\] sky130_fd_sc_hd__dfrtp_1
X_7855_ net108 seq.clk_div.next_count\[12\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6806_ sound2.count_m\[2\] _2857_ _3117_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4998_ _1533_ _1534_ _1504_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7786_ net113 inputcont.u1.ff_intermediate\[8\] net74 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6737_ _3084_ _3085_ net55 _3087_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3949_ _0459_ _0481_ inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1 vccd1 vccd1 _0613_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6668_ sound1.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6599_ sound1.sdiv.A\[8\] _2895_ _2964_ _2965_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__a22o_1
X_5619_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8338_ net139 _0438_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.M\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8269_ net123 _0369_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout92 net94 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_8
XFILLER_0_92_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout81 net3 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_8
XFILLER_0_64_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout70 net71 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_6
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ sound1.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _1341_ _1322_ _0948_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__a21o_1
X_7640_ _2139_ _2073_ vssd1 vssd1 vccd1 vccd1 _3707_ sky130_fd_sc_hd__or2b_1
X_4852_ _1005_ _1322_ _1339_ _0964_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_117_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7571_ _3662_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4783_ net42 _1313_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__nand2_1
X_6522_ sound1.sdiv.A\[26\] sound1.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6453_ sound1.count\[14\] _2201_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5404_ sound4.count\[18\] _1778_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6384_ _2809_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
X_8123_ net136 _0244_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[4\] sky130_fd_sc_hd__dfrtp_1
X_5335_ _1204_ _1786_ _1790_ _1014_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8054_ net116 _0196_ net77 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[8\] sky130_fd_sc_hd__dfrtp_2
X_5266_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__buf_6
X_4217_ _0786_ _0795_ _0801_ _0810_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__or4bb_1
X_7005_ _3265_ _3267_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__nand2_1
X_5197_ sound3.count\[0\] sound3.count\[1\] sound3.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1726_ sky130_fd_sc_hd__nand3_1
X_4148_ seq.player_3.state\[0\] _0753_ _0755_ vssd1 vssd1 vccd1 vccd1 seq.player_3.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_4079_ _0709_ vssd1 vssd1 vccd1 vccd1 seq_power_on sky130_fd_sc_hd__clkbuf_1
X_7907_ net128 _0070_ net89 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[0\] sky130_fd_sc_hd__dfrtp_1
X_7838_ net143 _0061_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7769_ net144 pm.next_count\[8\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5120_ _1016_ _1580_ _1570_ _1024_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__o22a_1
X_5051_ _0996_ _1025_ _1559_ _1577_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__o311a_1
X_4002_ _0655_ _0656_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ sound1.count_m\[15\] _2381_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5884_ sound4.count_m\[2\] sound4.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__and2b_1
X_4904_ sound2.count\[15\] _1454_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7623_ _2099_ _2131_ vssd1 vssd1 vccd1 vccd1 _3695_ sky130_fd_sc_hd__and2_1
X_4835_ _1317_ _1382_ _1385_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4766_ _1314_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__or2_4
X_7554_ sound4.count_m\[15\] _2843_ _2203_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__a21o_1
X_6505_ _1215_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7485_ _3634_ _3635_ vssd1 vssd1 vccd1 vccd1 _3636_ sky130_fd_sc_hd__nand2_1
X_4697_ _1263_ _1264_ _1256_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__and3b_1
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6436_ _0554_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6367_ _2783_ _2786_ _2795_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5318_ _1778_ _1824_ _1828_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8106_ net111 sound2.osc.next_count\[7\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6298_ _2695_ _2697_ _2694_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__a21oi_2
X_5249_ _1761_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
X_8037_ net109 _0179_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4620_ _0677_ _0958_ _1077_ _0981_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4551_ sound1.count\[13\] _1120_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__or2_1
X_7270_ _3437_ _3444_ _3445_ _3440_ sound3.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _0307_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4482_ net64 _1001_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__nor2_4
XFILLER_0_110_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6221_ wave_comb.u1.Q\[4\] _0573_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__nand2_1
X_6152_ sound1.sdiv.Q\[0\] sound1.sdiv.Q\[1\] _0579_ _2434_ vssd1 vssd1 vccd1 vccd1
+ _2587_ sky130_fd_sc_hd__o211a_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5103_ _1176_ _1562_ _1572_ _0954_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__o221a_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ sound3.divisor_m\[2\] sound3.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__or2b_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _1564_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__buf_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6985_ _3240_ vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _2181_ _2370_ _2371_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5867_ _2302_ _2300_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__and2b_1
X_7606_ _3681_ _3682_ _3683_ _2184_ sound4.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _0405_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5798_ _2238_ _2243_ _2244_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4818_ sound2.count\[12\] _1360_ _1368_ sound2.count\[7\] vssd1 vssd1 vccd1 vccd1
+ _1369_ sky130_fd_sc_hd__a2bb2o_1
X_7537_ sound3.sdiv.Q\[26\] _3654_ _3643_ sound3.sdiv.Q\[25\] _3406_ vssd1 vssd1 vccd1
+ vccd1 _0365_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4749_ _1256_ _1302_ _1303_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7468_ sound3.sdiv.A\[23\] _3595_ vssd1 vssd1 vccd1 vccd1 _3621_ sky130_fd_sc_hd__or2_1
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 beat_led[3] sky130_fd_sc_hd__clkbuf_4
X_6419_ seq.beat\[2\] _2832_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__nand2_1
X_7399_ sound3.divisor_m\[14\] _3552_ vssd1 vssd1 vccd1 vccd1 _3561_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 note4[0] sky130_fd_sc_hd__buf_2
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 note1[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6770_ _3112_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
X_3982_ _0554_ _0568_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ sound4.sdiv.Q\[12\] _2182_ _2185_ sound4.sdiv.Q\[11\] _2191_ vssd1 vssd1 vccd1
+ vccd1 _0012_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5652_ _2089_ _2134_ _2087_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8371_ net144 wave_comb.u1.next_dived net105 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.dived
+ sky130_fd_sc_hd__dfrtp_1
X_4603_ _0695_ net64 net63 vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__a21o_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5583_ _2063_ _2065_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7322_ sound3.divisor_m\[6\] _3483_ vssd1 vssd1 vccd1 vccd1 _3492_ sky130_fd_sc_hd__or2_1
X_4534_ _1073_ _1089_ _1104_ sound1.count\[0\] vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7253_ _1608_ vssd1 vssd1 vccd1 vccd1 _3433_ sky130_fd_sc_hd__inv_2
X_4465_ _0940_ _0944_ _1004_ _0974_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__a211o_1
X_7184_ sound3.count\[6\] _2863_ vssd1 vssd1 vccd1 vccd1 _3393_ sky130_fd_sc_hd__and2_1
X_6204_ _2631_ _2637_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__xnor2_1
X_4396_ _0966_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6135_ _2275_ _2570_ sound3.sdiv.Q\[1\] _0577_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__a2bb2o_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ sound2.sdiv.Q\[0\] _0578_ _2499_ _2501_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__a31o_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ net56 _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__or2_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6968_ _3224_ _3228_ _3235_ vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__nand3_1
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5919_ _2346_ sound4.count_m\[0\] _2347_ _2348_ _2354_ vssd1 vssd1 vccd1 vccd1 _2355_
+ sky130_fd_sc_hd__o2111a_1
X_6899_ _0578_ vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__buf_6
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4250_ seq.clk_div.count\[10\] seq.clk_div.count\[11\] _0829_ vssd1 vssd1 vccd1 vccd1
+ _0835_ sky130_fd_sc_hd__and3_1
X_4181_ _0700_ seq.clk_div.count\[0\] vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[0\]
+ sky130_fd_sc_hd__nor2_1
X_7940_ net126 _0103_ net87 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7871_ net108 inputcont.u1.ff_intermediate\[2\] net69 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6822_ sound2.count_m\[10\] _2857_ _3125_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__a21o_1
X_6753_ sound1.sdiv.A\[26\] _2895_ sound1.sdiv.next_dived _3101_ vssd1 vssd1 vccd1
+ vccd1 _0134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _0446_ _0628_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3896_ net65 vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__inv_2
X_6684_ _3040_ _3041_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__nand2_1
X_5704_ sound4.sdiv.Q\[3\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[2\] vssd1
+ vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5635_ sound4.divisor_m\[1\] sound4.divisor_m\[0\] _2036_ vssd1 vssd1 vccd1 vccd1
+ _2118_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8354_ net120 sound4.osc.next_count\[12\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_5566_ _2046_ _2048_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__nand2_1
X_7305_ _3474_ _3476_ vssd1 vssd1 vccd1 vccd1 _3477_ sky130_fd_sc_hd__or2_1
X_4517_ _0684_ _0939_ _1077_ _1081_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__o311a_1
X_5497_ sound4.count\[16\] _1988_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__nand2_1
X_8285_ net123 _0385_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[18\] sky130_fd_sc_hd__dfrtp_1
X_7236_ sound3.divisor_m\[9\] _3422_ _3419_ vssd1 vssd1 vccd1 vccd1 _3423_ sky130_fd_sc_hd__mux2_1
X_4448_ _0675_ _0945_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__nor2_4
XFILLER_0_95_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _0949_ _0909_ _0940_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nand3_4
X_7167_ sound2.sdiv.Q\[23\] _3167_ _3349_ sound2.sdiv.Q\[22\] _3130_ vssd1 vssd1 vccd1
+ vccd1 _0263_ sky130_fd_sc_hd__a221o_1
X_6118_ _2547_ sound3.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__or2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ sound2.sdiv.A\[20\] sound2.sdiv.A\[19\] _3329_ vssd1 vssd1 vccd1 vccd1 _3352_
+ sky130_fd_sc_hd__o21ai_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ sound2.count_m\[3\] _2484_ sound2.divisor_m\[1\] _2480_ vssd1 vssd1 vccd1
+ vccd1 _2485_ sky130_fd_sc_hd__a22o_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5420_ _0997_ _1781_ _1926_ _1930_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__o211a_2
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5351_ _1139_ _1786_ _1790_ _1134_ _1834_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__o221a_1
X_4302_ _0871_ _0872_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__nand2_1
X_8070_ net117 _0212_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[5\] sky130_fd_sc_hd__dfrtp_1
X_5282_ _1771_ _1775_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4233_ seq.clk_div.count\[6\] _0819_ _0813_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__o21ai_1
X_7021_ sound2.divisor_m\[13\] _3274_ vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__or2_1
X_4164_ seq.player_2.state\[2\] seq.player_2.state\[3\] vssd1 vssd1 vccd1 vccd1 _0766_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4095_ seq.player_8.state\[1\] seq.player_8.state\[2\] _0713_ seq.player_8.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a31o_1
X_7923_ net127 _0086_ net88 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7854_ net108 seq.clk_div.next_count\[11\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_7785_ net142 inputcont.u1.ff_intermediate\[14\] net103 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_MODE
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6805_ _1470_ _2843_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__nor2_1
X_6736_ sound1.sdiv.A\[22\] sound1.sdiv.A\[21\] sound1.sdiv.A\[20\] sound1.sdiv.A\[19\]
+ _3055_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__o41a_1
X_4997_ sound2.count\[12\] sound2.count\[13\] _1527_ sound2.count\[14\] vssd1 vssd1
+ vccd1 vccd1 _1534_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3948_ inputcont.INTERNAL_SYNCED_I\[4\] vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6667_ _2890_ _3025_ _3026_ _2894_ sound1.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _0123_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3879_ _0549_ _0534_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__nand2_4
X_6598_ _2962_ _2963_ _0866_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__a21oi_1
X_5618_ sound4.divisor_m\[5\] _2100_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8337_ net138 _0437_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[5\] sky130_fd_sc_hd__dfrtp_1
X_5549_ sound4.divisor_m\[12\] _2031_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8268_ net123 _0368_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[1\] sky130_fd_sc_hd__dfrtp_1
X_8199_ net142 _0320_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[14\] sky130_fd_sc_hd__dfrtp_1
X_7219_ _1641_ vssd1 vssd1 vccd1 vccd1 _3412_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout82 net3 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_8
Xfanout71 net76 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_6
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _0996_ _1025_ _1339_ _1393_ _0977_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__o32a_1
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4851_ _0869_ _1343_ _1345_ _1001_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3802_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1
+ vccd1 vccd1 _0481_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7570_ sound4.divisor_m\[5\] _1810_ _3419_ vssd1 vssd1 vccd1 vccd1 _3662_ sky130_fd_sc_hd__mux2_1
X_4782_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__clkbuf_8
X_6521_ _2893_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6452_ sound1.count_m\[13\] _2836_ _2851_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5403_ _1222_ _1913_ sound4.count\[17\] vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__o21a_1
X_6383_ pm.current_waveform\[0\] _2806_ _2808_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__mux2_1
X_8122_ net136 _0243_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5334_ _0686_ _1784_ _1781_ _1146_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__o22ai_1
X_8053_ net116 _0195_ net77 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[7\] sky130_fd_sc_hd__dfrtp_2
X_5265_ _1765_ _1775_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__or2_1
X_5196_ sound3.count\[0\] sound3.count\[1\] sound3.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1725_ sky130_fd_sc_hd__a21o_1
X_4216_ _0804_ _0805_ _0808_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__and4_1
X_7004_ _3265_ _3267_ vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4147_ seq.player_3.state\[1\] seq.player_3.state\[2\] seq.player_3.state\[3\] _0754_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__a311o_1
X_4078_ net1 net20 vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7906_ net115 _0069_ net76 vssd1 vssd1 vccd1 vccd1 seq.beat\[3\] sky130_fd_sc_hd__dfrtp_4
X_7837_ net143 _0060_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7768_ net144 pm.next_count\[7\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6719_ _3072_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7699_ _3747_ vssd1 vssd1 vccd1 vccd1 _3748_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5050_ _0993_ _1012_ _1578_ _1580_ _0948_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__o32a_1
X_4001_ pm.count\[6\] _0652_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__nor2_1
X_5952_ _2382_ _2384_ _2386_ _2387_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__and4_1
X_4903_ _0683_ _1316_ _1451_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__a211o_2
XFILLER_0_48_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5883_ _2318_ sound4.divisor_m\[6\] sound4.divisor_m\[5\] _2312_ vssd1 vssd1 vccd1
+ vccd1 _2319_ sky130_fd_sc_hd__a22o_1
X_7622_ _3681_ _3693_ _3694_ _2184_ sound4.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _0410_
+ sky130_fd_sc_hd__a32o_1
X_4834_ _1151_ _1323_ _1339_ _1095_ _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4765_ _1314_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nor2_4
X_7553_ sound4.count_m\[14\] _3403_ _2202_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6504_ _2883_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7484_ sound3.sdiv.A\[25\] _3595_ vssd1 vssd1 vccd1 vccd1 _3635_ sky130_fd_sc_hd__or2_1
X_4696_ sound1.count\[0\] sound1.count\[1\] sound1.count\[2\] sound1.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6435_ sound1.count_m\[5\] _2836_ _2842_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6366_ _2779_ _2782_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5317_ _1154_ _1784_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8105_ net111 sound2.osc.next_count\[6\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6297_ _2726_ _2727_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__nand2_1
X_8036_ net109 _0178_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[9\] sky130_fd_sc_hd__dfrtp_1
X_5248_ _1721_ _1759_ _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__and3_1
X_5179_ _0680_ _0959_ _1574_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4550_ sound1.count\[13\] _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4481_ _0944_ _0969_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__or2_1
X_6220_ wave_comb.u1.Q\[3\] _2653_ _0645_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__mux2_1
X_6151_ sound1.sdiv.Q\[3\] _0579_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _0996_ _1550_ _1630_ _1632_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__o211a_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ sound3.count_m\[1\] sound3.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__or2b_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _1547_ _1563_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__or2_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6984_ _3248_ _3249_ vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__nand2_1
X_5935_ sound4.sdiv.Q\[1\] _0576_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__nand2_1
X_5866_ _2300_ _2302_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7605_ sound4.divisor_m\[0\] sound4.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3683_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4817_ _1362_ _1364_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__and3_1
X_5797_ _2238_ _2243_ _2244_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7536_ sound3.sdiv.Q\[25\] _3654_ _3643_ sound3.sdiv.Q\[24\] _3405_ vssd1 vssd1 vccd1
+ vccd1 _0364_ sky130_fd_sc_hd__a221o_1
X_4748_ sound1.count\[16\] _1299_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__or2_1
X_7467_ sound3.sdiv.A\[23\] _3463_ sound3.sdiv.next_dived _3620_ vssd1 vssd1 vccd1
+ vccd1 _0329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4679_ sound1.count\[4\] _1145_ _1249_ sound1.count\[12\] vssd1 vssd1 vccd1 vccd1
+ _1250_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6418_ seq.beat\[2\] _2832_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__or2_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 note4[1] sky130_fd_sc_hd__clkbuf_4
X_7398_ sound3.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _3560_ sky130_fd_sc_hd__inv_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 beat_led[4] sky130_fd_sc_hd__buf_2
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 note1[2] sky130_fd_sc_hd__clkbuf_4
X_6349_ _2772_ _2778_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8019_ net126 _0161_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3981_ net34 _0643_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__nor2_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ sound4.count\[4\] _2186_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5651_ _2093_ _2132_ _2133_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ _1009_ _1051_ _1106_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8370_ net119 rate_clk.next_count\[7\] net80 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_5582_ sound4.divisor_m\[12\] _2064_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__xor2_1
X_7321_ sound3.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _3491_ sky130_fd_sc_hd__inv_2
X_4533_ _1094_ _1099_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__and3_2
XFILLER_0_53_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7252_ _3432_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6203_ _2292_ _2634_ _2635_ _2636_ _2279_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__o32a_1
X_4464_ _0952_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__nor2_4
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7183_ sound3.count_m\[5\] _3132_ _3392_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__a21o_1
X_4395_ _0918_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6134_ _2516_ _2556_ _2569_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__o21a_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _2500_ sound2.sdiv.next_start vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__nor2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _0546_ _1546_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6967_ _3233_ _3234_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5918_ _2350_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6898_ sound2.divisor_m\[0\] sound2.sdiv.Q\[27\] _3171_ vssd1 vssd1 vccd1 vccd1 _3173_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _2181_ _2284_ _2285_ _2286_ _0645_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7519_ sound3.sdiv.Q\[8\] _3654_ _3643_ sound3.sdiv.Q\[7\] _3387_ vssd1 vssd1 vccd1
+ vccd1 _0347_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4180_ _0774_ _0773_ _0776_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_1.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7870_ net111 inputcont.u1.ff_intermediate\[1\] net72 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6821_ sound2.count\[10\] _2855_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6752_ _3098_ _3100_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3964_ _0626_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3895_ sound1.sdiv.C\[4\] sound1.sdiv.C\[3\] sound1.sdiv.C\[2\] _0564_ sound1.sdiv.C\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__a311oi_4
X_6683_ sound1.sdiv.A\[16\] _3039_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__or2_1
X_5703_ sound4.sdiv.Q\[2\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[1\] vssd1
+ vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5634_ sound4.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8353_ net119 sound4.osc.next_count\[11\] net80 vssd1 vssd1 vccd1 vccd1 sound4.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_7304_ sound3.divisor_m\[5\] _3475_ vssd1 vssd1 vccd1 vccd1 _3476_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ sound4.divisor_m\[17\] _2047_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4516_ _1082_ _1084_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__and3_1
X_8284_ net123 _0384_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[17\] sky130_fd_sc_hd__dfrtp_1
X_5496_ _1991_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7235_ _1714_ vssd1 vssd1 vccd1 vccd1 _3422_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4447_ _0674_ _0964_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nor2_4
X_7166_ sound2.sdiv.Q\[22\] _3167_ _3349_ sound2.sdiv.Q\[21\] _3129_ vssd1 vssd1 vccd1
+ vccd1 _0262_ sky130_fd_sc_hd__a221o_1
X_6117_ _2509_ sound3.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__or2_1
X_4378_ _0926_ _0936_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__nor2_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ sound2.sdiv.A\[20\] _3329_ _3343_ vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__o21bai_1
X_6048_ sound2.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__inv_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ net140 _0141_ net101 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5350_ _1804_ _1822_ _1852_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4301_ seq.player_1.state\[0\] seq.player_1.state\[1\] seq.player_1.state\[2\] seq.player_1.state\[3\]
+ _0698_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__o41a_1
XFILLER_0_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5281_ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4232_ seq.clk_div.count\[6\] _0819_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__and2_1
X_7020_ sound2.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4163_ seq.player_2.state\[2\] seq.player_2.state\[3\] _0764_ _0765_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_2.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_4094_ _0717_ _0716_ _0718_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_8.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_7922_ net126 _0085_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7853_ net108 seq.clk_div.next_count\[10\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4996_ sound2.count\[13\] sound2.count\[14\] _1530_ vssd1 vssd1 vccd1 vccd1 _1533_
+ sky130_fd_sc_hd__and3_1
X_7784_ net118 inputcont.INTERNAL_OCTAVE_INPUT net79 vssd1 vssd1 vccd1 vccd1 inputcont.u2.next_in
+ sky130_fd_sc_hd__dfrtp_1
X_6804_ sound2.count_m\[1\] _2857_ _3116_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__a21o_1
X_6735_ _3069_ _3073_ _3078_ _3081_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3947_ inputcont.INTERNAL_SYNCED_I\[10\] _0610_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6666_ _3014_ _3018_ _3024_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__a21o_1
X_3878_ _0545_ _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__and3_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6597_ _2962_ _2963_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__or2_1
X_5617_ sound4.divisor_m\[4\] _2026_ _2036_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8336_ net137 _0436_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[4\] sky130_fd_sc_hd__dfrtp_1
X_5548_ sound4.divisor_m\[11\] sound4.divisor_m\[10\] _2030_ vssd1 vssd1 vccd1 vccd1
+ _2031_ sky130_fd_sc_hd__or3_1
X_8267_ net123 _0367_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[0\] sky130_fd_sc_hd__dfrtp_1
X_7218_ _3411_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__clkbuf_1
X_5479_ _1977_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__inv_2
X_8198_ net133 _0319_ net94 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[13\] sky130_fd_sc_hd__dfrtp_1
X_7149_ sound2.sdiv.Q\[5\] _3168_ _3164_ sound2.sdiv.Q\[4\] vssd1 vssd1 vccd1 vccd1
+ _0245_ sky130_fd_sc_hd__a22o_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout72 net76 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_8
Xfanout83 net85 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_8
XFILLER_0_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout94 net95 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _0978_ _0944_ _1333_ _1347_ _0997_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__o32a_1
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3801_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\]
+ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__o31ai_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6520_ _2890_ _2891_ _2892_ _2894_ sound1.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _0108_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4781_ _1319_ _1331_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6451_ sound1.count\[13\] _2201_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6382_ _2807_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5402_ _1772_ _1773_ _1777_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__and3_1
X_8121_ net136 _0242_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5333_ _1011_ _1015_ _1842_ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8052_ net117 _0194_ net78 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[6\] sky130_fd_sc_hd__dfrtp_2
X_5264_ _1766_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__or2_1
X_5195_ _1724_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_4215_ _0806_ seq.clk_div.count\[9\] seq.tempo_select.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0809_ sky130_fd_sc_hd__a21o_1
X_7003_ sound2.divisor_m\[12\] _3266_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__xnor2_1
X_4146_ seq.player_3.state\[0\] _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__and2_1
X_4077_ _0708_ vssd1 vssd1 vccd1 vccd1 seq_play_on sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7905_ net115 _0068_ net76 vssd1 vssd1 vccd1 vccd1 seq.beat\[2\] sky130_fd_sc_hd__dfrtp_4
X_7836_ net143 _0059_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7767_ net144 pm.next_count\[6\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4979_ sound2.count\[8\] _1520_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__and2_1
X_6718_ sound1.sdiv.A\[20\] _3055_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__xor2_1
X_7698_ sound4.sdiv.C\[2\] sound4.sdiv.C\[1\] sound4.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3747_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6649_ sound1.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8319_ net124 _0419_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4000_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5951_ _2385_ sound1.divisor_m\[12\] sound1.count_m\[10\] _2378_ vssd1 vssd1 vccd1
+ vccd1 _2387_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4902_ _0688_ _1334_ _1452_ _1317_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__o211ai_1
X_5882_ sound4.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7621_ _2129_ _3692_ vssd1 vssd1 vccd1 vccd1 _3694_ sky130_fd_sc_hd__or2b_1
X_4833_ _1134_ _1343_ _1333_ _1146_ _1383_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7552_ sound4.count_m\[13\] _3403_ _2200_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__a21o_1
X_4764_ _0698_ _0504_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__or2_2
X_7483_ sound3.sdiv.A\[25\] _3595_ vssd1 vssd1 vccd1 vccd1 _3634_ sky130_fd_sc_hd__nand2_1
X_6503_ sound1.divisor_m\[14\] _2882_ _2864_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6434_ sound1.count\[5\] _2201_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__and2_1
X_4695_ sound1.count\[0\] sound1.count\[1\] sound1.count\[2\] sound1.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6365_ _2762_ _2791_ _2792_ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6296_ _2725_ _2717_ _2721_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__or3_1
X_5316_ _1166_ _1800_ _1796_ _0677_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__o22a_1
X_8104_ net111 sound2.osc.next_count\[5\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5247_ sound3.count\[18\] _1756_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__nand2_1
X_8035_ net109 _0177_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[8\] sky130_fd_sc_hd__dfrtp_1
X_5178_ _1158_ _1578_ _1550_ _1004_ _1708_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__o221a_1
X_4129_ seq.player_5.state\[2\] _0740_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7819_ net114 seq.player_4.next_state\[1\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4480_ sound1.count\[2\] _1032_ _1050_ sound1.count\[11\] vssd1 vssd1 vccd1 vccd1
+ _1051_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6150_ _2289_ _2583_ _2584_ _2290_ sound4.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1 _2585_
+ sky130_fd_sc_hd__a32o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _1129_ _1580_ _1570_ _1182_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__o221a_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ sound3.count_m\[0\] vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__inv_2
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _0698_ _0540_ _1557_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__o21ai_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6983_ _3244_ _3247_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5934_ _2314_ _2321_ _2356_ _2369_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__a31o_1
X_5865_ _2275_ _2292_ _2301_ sound3.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__a2bb2o_1
X_7604_ sound4.divisor_m\[0\] sound4.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3682_ sky130_fd_sc_hd__nand2_1
X_4816_ _1085_ _1322_ _1339_ _1078_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5796_ wave_comb.u1.A\[6\] _2224_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7535_ sound3.sdiv.Q\[24\] _3654_ _3643_ sound3.sdiv.Q\[23\] _3404_ vssd1 vssd1 vccd1
+ vccd1 _0363_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4747_ sound1.count\[16\] _1299_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7466_ _3618_ _3619_ vssd1 vssd1 vccd1 vccd1 _3620_ sky130_fd_sc_hd__xnor2_1
X_4678_ _1239_ _1241_ _1244_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__and4_2
X_7397_ _3437_ _3558_ _3559_ _3440_ sound3.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _0320_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6417_ _2831_ _2832_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 note1[3] sky130_fd_sc_hd__clkbuf_4
X_6348_ sound4.sdiv.Q\[8\] _2290_ _2369_ _2773_ _2777_ vssd1 vssd1 vccd1 vccd1 _2778_
+ sky130_fd_sc_hd__a221oi_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 note4[2] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 beat_led[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6279_ _2708_ _2710_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__xnor2_1
X_8018_ net126 _0160_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _0630_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5650_ sound4.sdiv.A\[6\] _2092_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__nand2_1
X_4601_ _1121_ _1122_ _1145_ sound1.count\[4\] _1171_ vssd1 vssd1 vccd1 vccd1 _1172_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5581_ _2036_ _2031_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__nand2_1
X_7320_ _3437_ _3489_ _3490_ _3440_ sound3.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _0312_
+ sky130_fd_sc_hd__a32o_1
X_4532_ _0981_ _1041_ _1101_ _0990_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7251_ sound3.divisor_m\[15\] _3431_ _3419_ vssd1 vssd1 vccd1 vccd1 _3432_ sky130_fd_sc_hd__mux2_1
X_4463_ _0685_ _0677_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6202_ sound3.sdiv.Q\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7182_ sound3.count\[5\] _2863_ vssd1 vssd1 vccd1 vccd1 _3392_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4394_ _0909_ _0955_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6133_ _2544_ _2568_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ sound2.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__inv_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _0699_ net46 vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__and2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _3229_ _3232_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__nand2_1
X_5917_ _2346_ sound4.count_m\[0\] _2351_ _2352_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6897_ _3165_ _3171_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5848_ net30 net31 vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5779_ _2225_ _2222_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7518_ _0577_ vssd1 vssd1 vccd1 vccd1 _3654_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7449_ _3599_ _3602_ _3605_ vssd1 vssd1 vccd1 vccd1 _3606_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6820_ sound2.count_m\[9\] _2857_ _3124_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6751_ _3089_ _3092_ _3099_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ _0456_ _0625_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6682_ sound1.sdiv.A\[16\] _3039_ vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__nand2_1
X_3894_ sound1.sdiv.start vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__inv_2
X_5702_ sound4.sdiv.Q\[1\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[0\] vssd1
+ vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5633_ _2114_ _2115_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5564_ _2036_ _2034_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8352_ net119 sound4.osc.next_count\[10\] net80 vssd1 vssd1 vccd1 vccd1 sound4.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7303_ sound3.divisor_m\[4\] _3465_ _3448_ vssd1 vssd1 vccd1 vccd1 _3475_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4515_ _0952_ _1000_ _1003_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8283_ net123 _0383_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[16\] sky130_fd_sc_hd__dfrtp_1
X_5495_ _1779_ _1936_ _1989_ _1990_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7234_ _2843_ _1706_ _3421_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o21ai_1
X_4446_ _0683_ _0947_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__nor2_2
X_7165_ sound2.sdiv.Q\[21\] _3167_ _3349_ sound2.sdiv.Q\[20\] _3128_ vssd1 vssd1 vccd1
+ vccd1 _0261_ sky130_fd_sc_hd__a221o_1
X_4377_ _0944_ _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__or2_4
X_6116_ _2545_ sound3.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__or2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ sound2.sdiv.A\[21\] _3329_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__xnor2_1
X_6047_ sound2.divisor_m\[1\] _2480_ _2481_ _2482_ vssd1 vssd1 vccd1 vccd1 _2483_
+ sky130_fd_sc_hd__o211ai_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ net137 sound2.sdiv.next_dived net98 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.dived
+ sky130_fd_sc_hd__dfrtp_1
X_6949_ _3206_ _3209_ _3217_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4300_ _0702_ seq.encode.play _0870_ inputcont.INTERNAL_SYNCED_I\[0\] vssd1 vssd1
+ vccd1 vccd1 _0871_ sky130_fd_sc_hd__a31o_2
X_5280_ _1767_ _1773_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__or2_1
X_4231_ _0821_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4162_ seq.player_2.state\[1\] _0762_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__nor2_1
X_4093_ _0698_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__clkbuf_8
X_7921_ net126 _0084_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7852_ net108 seq.clk_div.next_count\[9\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_7783_ net142 inputcont.INTERNAL_MODE net103 vssd1 vssd1 vccd1 vccd1 inputcont.u3.next_in
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4995_ sound2.count\[13\] _1530_ _1532_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[13\]
+ sky130_fd_sc_hd__a21oi_1
X_6803_ sound2.count\[1\] _2855_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__and2_1
X_6734_ sound1.sdiv.A\[23\] _3055_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__nand2_1
X_3946_ _0608_ _0609_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6665_ _3014_ _3018_ _3024_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3877_ _0518_ _0527_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6596_ _2946_ _2953_ _2951_ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__o21a_1
X_5616_ _2097_ _2098_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8335_ net137 _0435_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5547_ sound4.divisor_m\[9\] _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__or2_1
X_8266_ net141 _0366_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[27\] sky130_fd_sc_hd__dfrtp_1
X_5478_ sound4.count\[12\] _1973_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7217_ sound3.divisor_m\[2\] _3410_ _3142_ vssd1 vssd1 vccd1 vccd1 _3411_ sky130_fd_sc_hd__mux2_1
X_4429_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__buf_4
X_8197_ net133 _0318_ net94 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[12\] sky130_fd_sc_hd__dfrtp_1
X_7148_ sound2.sdiv.Q\[4\] _3168_ _3164_ sound2.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1
+ _0244_ sky130_fd_sc_hd__a22o_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7079_ sound2.sdiv.A\[19\] _3329_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout73 net76 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_4
XFILLER_0_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout95 net3 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_8
Xfanout84 net85 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_8
XFILLER_0_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[6\] vssd1 vssd1 vccd1 vccd1 _0479_
+ sky130_fd_sc_hd__o21ai_4
X_4780_ _1315_ _1330_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6450_ sound1.count_m\[12\] _2836_ _2850_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6381_ wave_comb.u1.dived _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__and3_1
X_5401_ sound4.count\[7\] _1897_ _1903_ sound4.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1912_ sky130_fd_sc_hd__a2bb2o_1
X_8120_ net136 _0241_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5332_ _1200_ _1792_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8051_ net112 _0193_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[5\] sky130_fd_sc_hd__dfrtp_2
X_5263_ _0698_ _0673_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__nor2_1
X_5194_ _1721_ _1722_ _1723_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__and3_1
X_4214_ seq.tempo_select.state\[1\] _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__nand2_1
X_7002_ sound2.divisor_m\[11\] _3256_ _3177_ vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__o21a_1
X_4145_ seq.encode.keys_edge_det\[4\] inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1
+ vccd1 vccd1 _0753_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ net1 net19 vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7904_ net115 _0067_ net76 vssd1 vssd1 vccd1 vccd1 seq.beat\[1\] sky130_fd_sc_hd__dfrtp_4
X_7835_ net143 _0058_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7766_ net144 pm.next_count\[5\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_4978_ _1520_ _1521_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[7\] sky130_fd_sc_hd__nor2_1
XFILLER_0_128_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6717_ sound1.sdiv.A\[20\] _2895_ _3069_ _3071_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7697_ sound4.sdiv.C\[1\] sound4.sdiv.C\[0\] sound4.sdiv.C\[2\] vssd1 vssd1 vccd1
+ vccd1 _3746_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3929_ _0593_ net57 _0590_ _0521_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__o31a_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6648_ _2890_ _3008_ _3009_ _2894_ sound1.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _0121_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6579_ sound1.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8318_ net124 _0418_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8249_ net135 _0349_ net96 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5950_ _2383_ sound1.count_m\[12\] _2385_ sound1.divisor_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2386_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4901_ _1138_ _1324_ _1315_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7620_ _3692_ _2129_ vssd1 vssd1 vccd1 vccd1 _3693_ sky130_fd_sc_hd__or2b_1
X_5881_ _2315_ sound4.divisor_m\[8\] _2316_ sound4.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4832_ _1012_ _1338_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__or2_2
X_7551_ sound4.count_m\[12\] _3403_ _2199_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__a21o_1
X_7482_ sound3.sdiv.A\[25\] _3463_ sound3.sdiv.next_dived _3633_ vssd1 vssd1 vccd1
+ vccd1 _0331_ sky130_fd_sc_hd__a22o_1
X_6502_ _1235_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__inv_2
X_4694_ _1262_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6433_ sound1.count_m\[4\] _2836_ _2841_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6364_ _2772_ _2778_ vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6295_ _2717_ _2721_ _2725_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__o21ai_1
X_5315_ _0685_ _1769_ _1794_ _1077_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__o221a_1
X_8103_ net111 sound2.osc.next_count\[4\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_5246_ sound3.count\[18\] _1756_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8034_ net109 _0176_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[7\] sky130_fd_sc_hd__dfrtp_1
X_5177_ _1014_ _1567_ _1570_ _1083_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__o22a_1
X_4128_ seq.player_5.state\[2\] seq.player_5.state\[3\] vssd1 vssd1 vccd1 vccd1 _0742_
+ sky130_fd_sc_hd__nand2_1
X_4059_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__buf_12
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7818_ net114 seq.player_4.next_state\[0\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7749_ net143 _0034_ net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6080_ _2510_ _2512_ _2515_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__nand3b_1
X_5100_ _1026_ _1567_ _1574_ _1175_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__o22a_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6982_ _3244_ _3247_ vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__or2_1
X_5933_ sound4.count_m\[17\] _2349_ sound4.count_m\[18\] _2368_ vssd1 vssd1 vccd1
+ vccd1 _2369_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5864_ sound3.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7603_ _1764_ vssd1 vssd1 vccd1 vccd1 _3681_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4815_ _1083_ _1321_ _1341_ _1079_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7534_ sound3.sdiv.Q\[23\] _3654_ _3643_ sound3.sdiv.Q\[22\] _3402_ vssd1 vssd1 vccd1
+ vccd1 _0362_ sky130_fd_sc_hd__a221o_1
X_5795_ wave_comb.u1.next_dived _2242_ _2243_ _0573_ wave_comb.u1.A\[6\] vssd1 vssd1
+ vccd1 vccd1 _0034_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4746_ _1301_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7465_ sound3.sdiv.A\[21\] _3595_ _3616_ vssd1 vssd1 vccd1 vccd1 _3619_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4677_ _0992_ _1245_ _1246_ _1247_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__o211a_1
X_7396_ _3546_ _3549_ _3557_ vssd1 vssd1 vccd1 vccd1 _3559_ sky130_fd_sc_hd__a21o_1
X_6416_ seq.beat\[1\] seq.beat\[0\] _2830_ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__and3_1
X_6347_ _2292_ _2776_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__nor2_1
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 beat_led[6] sky130_fd_sc_hd__clkbuf_4
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 note2[0] sky130_fd_sc_hd__clkbuf_4
X_6278_ _2672_ _2675_ _2709_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__o21a_1
X_5229_ sound3.count\[12\] _1744_ _1721_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__o21ai_1
X_8017_ net126 _0159_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4600_ sound1.count\[10\] _1157_ _1170_ sound1.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _1171_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5580_ sound4.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__inv_2
X_4531_ _0977_ _0950_ _0996_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7250_ _1615_ vssd1 vssd1 vccd1 vccd1 _3431_ sky130_fd_sc_hd__inv_2
X_4462_ _0679_ _0971_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__or2_2
XFILLER_0_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6201_ sound3.sdiv.Q\[3\] _0577_ _2633_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7181_ sound3.count_m\[4\] _3132_ _3391_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__a21o_1
X_4393_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__buf_8
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6132_ _2552_ _2567_ _2546_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__a21oi_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _2459_ _2469_ _2487_ _2498_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__a31o_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _1545_ vssd1 vssd1 vccd1 vccd1 sound3.sdiv.next_dived sky130_fd_sc_hd__buf_4
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6965_ _3229_ _3232_ vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__or2_2
X_5916_ sound4.divisor_m\[2\] sound4.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6896_ sound2.sdiv.A\[0\] _3170_ vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5847_ _2181_ _2284_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5778_ _2227_ _2228_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7517_ sound3.sdiv.Q\[7\] _3440_ _3437_ sound3.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1
+ _0346_ sky130_fd_sc_hd__a22o_1
X_4729_ _1287_ _1288_ _1256_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7448_ sound3.sdiv.A\[18\] _3595_ _3600_ _3603_ _3604_ vssd1 vssd1 vccd1 vccd1 _3605_
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_114_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7379_ sound3.divisor_m\[12\] sound3.divisor_m\[11\] _3526_ vssd1 vssd1 vccd1 vccd1
+ _3543_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6750_ sound1.sdiv.A\[24\] sound1.sdiv.A\[23\] _3055_ vssd1 vssd1 vccd1 vccd1 _3099_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5701_ _2182_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ _0456_ _0625_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__or2_1
X_3893_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__inv_2
X_6681_ _3038_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5632_ _2111_ _2113_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8351_ net120 sound4.osc.next_count\[9\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_5563_ sound4.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7302_ sound3.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 _3474_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4514_ _0959_ _0952_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5494_ sound4.count\[15\] _1984_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__or2_1
X_8282_ net122 _0382_ net83 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[15\] sky130_fd_sc_hd__dfrtp_1
X_7233_ sound3.divisor_m\[8\] _2843_ vssd1 vssd1 vccd1 vccd1 _3421_ sky130_fd_sc_hd__nand2_1
X_4445_ _1015_ _0869_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__nand2_4
XFILLER_0_41_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4376_ _0675_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nor2_4
X_7164_ sound2.sdiv.Q\[20\] _3167_ _3349_ sound2.sdiv.Q\[19\] _3127_ vssd1 vssd1 vccd1
+ vccd1 _0260_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6115_ sound3.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__inv_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _1311_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__buf_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ sound2.divisor_m\[2\] sound2.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__or2b_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ net134 sound1.osc.next_count\[18\] net95 vssd1 vssd1 vccd1 vccd1 sound1.count\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_6948_ _3206_ _3209_ _3217_ vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__nand3_1
X_6879_ _3159_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4230_ _0819_ _0820_ _0813_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__and3b_1
X_4161_ seq.player_2.state\[0\] seq.player_2.state\[1\] _0761_ vssd1 vssd1 vccd1 vccd1
+ _0764_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ seq.player_8.state\[2\] _0715_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__xor2_1
X_7920_ net126 _0083_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[13\] sky130_fd_sc_hd__dfrtp_1
X_7851_ net108 seq.clk_div.next_count\[8\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6802_ sound2.count_m\[0\] _2857_ _3115_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7782_ net137 _0056_ net98 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4994_ sound2.count\[13\] _1530_ _1504_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__o21ai_1
X_6733_ sound1.sdiv.A\[23\] _3055_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__or2_1
X_3945_ inputcont.INTERNAL_SYNCED_I\[6\] inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1
+ vccd1 vccd1 _0609_ sky130_fd_sc_hd__nor2_1
X_6664_ _3022_ _3023_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5615_ sound4.sdiv.A\[5\] _2096_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__or2_1
X_3876_ _0520_ _0541_ net57 vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6595_ _2960_ _2961_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8334_ net138 _0434_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5546_ sound4.divisor_m\[8\] sound4.divisor_m\[7\] _2028_ vssd1 vssd1 vccd1 vccd1
+ _2029_ sky130_fd_sc_hd__or3_1
X_8265_ net141 _0365_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5477_ _1976_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
X_7216_ _1655_ vssd1 vssd1 vccd1 vccd1 _3410_ sky130_fd_sc_hd__inv_2
X_4428_ _0940_ _0974_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__or2_1
X_8196_ net133 _0317_ net94 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[11\] sky130_fd_sc_hd__dfrtp_1
X_7147_ sound2.sdiv.Q\[3\] _3168_ sound2.sdiv.next_dived sound2.sdiv.Q\[2\] vssd1
+ vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__a22o_1
X_4359_ _0928_ _0929_ _0892_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__o21a_1
X_7078_ sound2.sdiv.A\[19\] _3168_ sound2.sdiv.next_dived _3334_ vssd1 vssd1 vccd1
+ vccd1 _0226_ sky130_fd_sc_hd__a22o_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _2463_ sound2.divisor_m\[6\] sound2.divisor_m\[5\] _2464_ vssd1 vssd1 vccd1
+ vccd1 _2465_ sky130_fd_sc_hd__a22o_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout74 net75 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_6
XFILLER_0_107_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout96 net97 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_6
Xfanout85 net3 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_6
XFILLER_0_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6380_ _2280_ _2274_ _2805_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__mux2_1
X_5400_ sound4.count\[15\] _1891_ _1897_ sound4.count\[7\] _1910_ vssd1 vssd1 vccd1
+ vccd1 _1911_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5331_ _1771_ _1775_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__nor2_1
X_8050_ net112 _0192_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[4\] sky130_fd_sc_hd__dfrtp_4
X_7001_ sound2.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__inv_2
X_5262_ _0698_ _0587_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__or2_4
X_5193_ sound3.count\[0\] sound3.count\[1\] vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__nand2_1
X_4213_ seq.tempo_select.state\[0\] _0802_ seq.clk_div.count\[9\] _0806_ vssd1 vssd1
+ vccd1 vccd1 _0807_ sky130_fd_sc_hd__a211o_1
X_4144_ _0750_ _0749_ _0752_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_4.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4075_ _0706_ _0707_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__nor2_1
X_7903_ net115 _0066_ net76 vssd1 vssd1 vccd1 vccd1 seq.beat\[0\] sky130_fd_sc_hd__dfrtp_4
X_7834_ net144 _0057_ net105 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7765_ net144 pm.next_count\[4\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[4\] sky130_fd_sc_hd__dfrtp_1
X_6716_ _0866_ _3070_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__nor2_1
X_4977_ sound2.count\[7\] _1518_ _1504_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__o21ai_1
X_7696_ _3681_ _3744_ _3745_ _2184_ sound4.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 _0433_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3928_ _0545_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__inv_2
X_6647_ _2996_ _3000_ _3007_ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3859_ _0520_ _0524_ _0528_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a211o_1
X_6578_ _2942_ _2943_ _2940_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__o21a_1
X_5529_ _2012_ pm.current_waveform\[3\] vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__and2_1
X_8317_ net124 _0417_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[12\] sky130_fd_sc_hd__dfrtp_1
X_8248_ net135 _0348_ net96 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[9\] sky130_fd_sc_hd__dfrtp_1
X_8179_ net133 _0300_ net94 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4900_ net63 _1449_ _1450_ _0944_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__a22o_1
X_5880_ sound4.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4831_ _1053_ _1347_ _1341_ _0983_ _1381_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7550_ sound4.count_m\[11\] _3403_ _2198_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__a21o_1
X_4762_ _0698_ _0507_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nor2_1
X_7481_ _3629_ _3632_ vssd1 vssd1 vccd1 vccd1 _3633_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6501_ _2881_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
X_4693_ _1256_ _1260_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6432_ sound1.count\[4\] _2201_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6363_ _2766_ _2771_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8102_ net111 sound2.osc.next_count\[3\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6294_ _2289_ _2723_ _2724_ _2293_ sound1.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 _2725_
+ sky130_fd_sc_hd__a32o_1
X_5314_ _0997_ _1777_ _1792_ _1159_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__o22a_1
X_5245_ _1758_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_8033_ net109 _0175_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5176_ sound3.count\[8\] _1706_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__xnor2_1
X_4127_ seq.player_5.state\[2\] seq.player_5.state\[3\] _0740_ _0741_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_5.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4058_ _0698_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__inv_4
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7817_ net114 seq.player_5.next_state\[3\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_5.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7748_ net139 _0033_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7679_ _3733_ _3734_ sound4.sdiv.A\[22\] _2183_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_62_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _1547_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ sound2.divisor_m\[10\] _3246_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5932_ _2323_ _2367_ _2350_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5863_ _2281_ _2299_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5794_ _2240_ _2241_ _2239_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7602_ _3680_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _0680_ _1336_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__or2_1
X_7533_ sound3.sdiv.Q\[22\] _3654_ _3643_ sound3.sdiv.Q\[21\] _3401_ vssd1 vssd1 vccd1
+ vccd1 _0361_ sky130_fd_sc_hd__a221o_1
X_4745_ _1299_ _1300_ _1256_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7464_ sound3.sdiv.A\[22\] _3595_ vssd1 vssd1 vccd1 vccd1 _3618_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4676_ _0967_ _1004_ _1133_ _1110_ _0976_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7395_ _3546_ _3549_ _3557_ vssd1 vssd1 vccd1 vccd1 _3558_ sky130_fd_sc_hd__nand3_1
XFILLER_0_114_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6415_ seq.beat\[0\] _2830_ seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__a21oi_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 beat_led[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6346_ _2774_ _2775_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6277_ _2668_ _2671_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__or2_1
X_8016_ net126 _0158_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[17\] sky130_fd_sc_hd__dfrtp_1
X_5228_ sound3.count\[12\] _1744_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__and2_1
X_5159_ _1684_ _1689_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4530_ _1100_ _0959_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__or2_4
X_4461_ _0990_ _0973_ _0939_ _1010_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__o221a_2
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6200_ sound3.sdiv.Q\[3\] _0577_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__and3_1
X_7180_ sound3.count\[4\] _2863_ vssd1 vssd1 vccd1 vccd1 _3391_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6131_ _2560_ net60 _2554_ _2566_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__a31o_1
X_4392_ _0676_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__or2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _2472_ _2497_ _2477_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__a21o_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _0575_ _0563_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__nor2_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6964_ sound2.divisor_m\[8\] _3231_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5915_ sound4.count_m\[1\] sound4.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__and2b_1
X_6895_ sound2.divisor_m\[1\] _3169_ vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__xnor2_1
X_5846_ _2275_ _2282_ _2283_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5777_ wave_comb.u1.A\[3\] _2224_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7516_ sound3.sdiv.Q\[6\] _3440_ _3437_ sound3.sdiv.Q\[5\] vssd1 vssd1 vccd1 vccd1
+ _0345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4728_ sound1.count\[9\] sound1.count\[10\] _1278_ sound1.count\[11\] vssd1 vssd1
+ vccd1 vccd1 _1288_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7447_ sound3.sdiv.A\[18\] _3595_ _3589_ vssd1 vssd1 vccd1 vccd1 _3604_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4659_ _0680_ _0950_ _0939_ _0684_ _0992_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7378_ sound3.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _3542_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _2472_ _2497_ _2477_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ inputcont.INTERNAL_SYNCED_I\[9\] _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__xnor2_1
X_5700_ _0576_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3892_ sound3.sdiv.C\[4\] sound3.sdiv.C\[3\] sound3.sdiv.C\[2\] _0561_ sound3.sdiv.C\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__a311oi_4
X_6680_ sound1.divisor_m\[17\] _3037_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5631_ _2111_ _2113_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5562_ sound4.sdiv.A\[21\] _2038_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8350_ net120 sound4.osc.next_count\[8\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7301_ _3471_ _3473_ sound3.sdiv.A\[4\] _3463_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4513_ _0950_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8281_ net122 _0381_ net83 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7232_ _3420_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__clkbuf_1
X_5493_ _1988_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4444_ _0695_ _0964_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__nand2_8
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4375_ _0945_ net64 vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__nor2_8
X_7163_ sound2.sdiv.Q\[19\] _3167_ _3349_ sound2.sdiv.Q\[18\] _3126_ vssd1 vssd1 vccd1
+ vccd1 _0259_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6114_ _2544_ _2546_ _2548_ _2549_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _3164_ _3347_ _3348_ _3174_ sound2.sdiv.A\[21\] vssd1 vssd1 vccd1 vccd1 _0228_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ sound2.count_m\[1\] sound2.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ net125 sound1.osc.next_count\[17\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6947_ _3215_ _3216_ vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6878_ sound2.divisor_m\[14\] _1422_ _3142_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5829_ _2269_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4160_ seq.player_2.state\[0\] _0761_ _0763_ vssd1 vssd1 vccd1 vccd1 seq.player_2.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ seq.player_8.state\[2\] seq.player_8.state\[3\] vssd1 vssd1 vccd1 vccd1 _0717_
+ sky130_fd_sc_hd__nand2_1
X_7850_ net108 seq.clk_div.next_count\[7\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6801_ sound2.count\[0\] _2855_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__and2_1
X_7781_ net137 _0055_ net98 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[10\] sky130_fd_sc_hd__dfrtp_1
X_4993_ _1530_ _1531_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[12\] sky130_fd_sc_hd__nor2_1
X_6732_ sound1.sdiv.A\[23\] _2895_ sound1.sdiv.next_dived _3083_ vssd1 vssd1 vccd1
+ vccd1 _0131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3944_ inputcont.INTERNAL_SYNCED_I\[6\] inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1
+ vccd1 vccd1 _0608_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6663_ _3019_ _3021_ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3875_ _0546_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__inv_2
XFILLER_0_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5614_ sound4.sdiv.A\[5\] _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6594_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8333_ net138 _0433_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5545_ sound4.divisor_m\[6\] _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8264_ net140 _0364_ net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ _1779_ _1936_ _1974_ _1975_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8195_ net133 _0316_ net94 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[10\] sky130_fd_sc_hd__dfrtp_1
X_7215_ _3409_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__clkbuf_1
X_4427_ _0959_ _0992_ _0993_ _0994_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__o32a_1
X_7146_ sound2.sdiv.Q\[2\] _3168_ sound2.sdiv.next_dived sound2.sdiv.Q\[1\] vssd1
+ vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__a22o_1
X_4358_ select1.sequencer_on seq.player_6.state\[3\] _0893_ vssd1 vssd1 vccd1 vccd1
+ _0929_ sky130_fd_sc_hd__and3_1
X_7077_ _3332_ _3333_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__xnor2_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ seq.encode.keys_edge_det\[0\] seq.encode.keys_sync\[0\] vssd1 vssd1 vccd1
+ vccd1 _0863_ sky130_fd_sc_hd__or2b_1
X_6028_ sound2.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7979_ net125 sound1.osc.next_count\[0\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[0\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout97 net106 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_8
Xfanout86 net95 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_8
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout75 net76 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_8
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5330_ sound4.count\[9\] _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__xnor2_1
X_5261_ _1769_ _1770_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__and3_1
X_7000_ sound2.sdiv.A\[11\] _3168_ sound2.sdiv.next_dived _3264_ vssd1 vssd1 vccd1
+ vccd1 _0218_ sky130_fd_sc_hd__a22o_1
X_4212_ seq.clk_div.count\[8\] vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__inv_2
X_5192_ sound3.count\[0\] sound3.count\[1\] vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4143_ seq.player_4.state\[1\] seq.player_4.state\[2\] _0746_ seq.player_4.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__a31o_1
X_4074_ _0705_ _0707_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__nor2_1
X_7902_ net140 sound1.sdiv.next_dived net101 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.dived
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7833_ net113 seq.player_1.next_state\[3\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_1.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7764_ net144 pm.next_count\[3\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6715_ _3068_ _3063_ _3065_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4976_ sound2.count\[6\] sound2.count\[7\] _1515_ vssd1 vssd1 vccd1 vccd1 _1520_
+ sky130_fd_sc_hd__and3_1
X_7695_ sound4.sdiv.C\[1\] sound4.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3745_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3927_ _0590_ _0591_ _0523_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__o21a_1
X_6646_ _2996_ _3000_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3858_ _0529_ _0530_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__and3_1
X_3789_ net1 wave.mode\[0\] vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6577_ _2944_ _2945_ sound1.sdiv.A\[6\] _2895_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__a2bb2o_1
X_5528_ pm.count\[3\] vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8316_ net118 _0416_ net79 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8247_ net141 _0347_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[8\] sky130_fd_sc_hd__dfrtp_1
X_5459_ sound4.count\[7\] sound4.count\[8\] _1955_ vssd1 vssd1 vccd1 vccd1 _1962_
+ sky130_fd_sc_hd__and3_1
X_8178_ net133 _0299_ net94 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[12\] sky130_fd_sc_hd__dfrtp_2
X_7129_ _3349_ _3375_ _3376_ _3174_ sound2.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 _0235_
+ sky130_fd_sc_hd__a32o_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4830_ _1042_ _1336_ _1345_ _1154_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4761_ _0699_ net42 vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__and2_1
X_7480_ _3630_ _3631_ vssd1 vssd1 vccd1 vccd1 _3632_ sky130_fd_sc_hd__and2b_1
X_6500_ sound1.divisor_m\[13\] _1120_ _2864_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__mux2_1
X_4692_ sound1.count\[0\] sound1.count\[1\] sound1.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1261_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6431_ sound1.count_m\[3\] _2836_ _2840_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6362_ _2764_ _2765_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5313_ _1126_ _1781_ _1790_ _1165_ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8101_ net111 sound2.osc.next_count\[2\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6293_ sound1.sdiv.Q\[6\] _0579_ _2722_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__a21o_1
X_5244_ _1756_ _1757_ _1721_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8032_ net111 _0174_ net72 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[5\] sky130_fd_sc_hd__dfrtp_1
X_5175_ _1701_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__and2_1
X_4126_ seq.player_5.state\[1\] _0738_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4057_ select1.sequencer_on vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__buf_8
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7816_ net114 seq.player_5.next_state\[2\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_5.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7747_ net139 _0032_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4959_ _1470_ _1506_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7678_ _2045_ _2171_ _3732_ _1763_ vssd1 vssd1 vccd1 vccd1 _3734_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6629_ _2991_ _2992_ sound1.sdiv.A\[11\] _2895_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_6_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6980_ _3177_ _3245_ vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__and2_1
X_5931_ _2360_ net61 _2345_ _2366_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5862_ _2297_ _2298_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__nor2_1
X_5793_ _2239_ _2240_ _2241_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__nand3_1
X_7601_ sound4.divisor_m\[18\] _1913_ _2186_ vssd1 vssd1 vccd1 vccd1 _3680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4813_ _0960_ _1333_ _1345_ _0952_ _1363_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7532_ sound3.sdiv.Q\[21\] _3654_ _3643_ sound3.sdiv.Q\[20\] _3400_ vssd1 vssd1 vccd1
+ vccd1 _0360_ sky130_fd_sc_hd__a221o_1
X_4744_ sound1.count\[15\] _1296_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7463_ _3615_ _3617_ sound3.sdiv.A\[22\] _3463_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_114_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4675_ _0994_ _1025_ _1038_ _0954_ _0990_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__o32a_1
XFILLER_0_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7394_ _3555_ _3556_ vssd1 vssd1 vccd1 vccd1 _3557_ sky130_fd_sc_hd__nand2_1
X_6414_ seq.beat\[0\] _2830_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6345_ sound4.sdiv.Q\[6\] _2641_ _2736_ vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6276_ _2703_ _2707_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__xor2_1
X_5227_ _1746_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
X_8015_ net126 _0157_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[16\] sky130_fd_sc_hd__dfrtp_1
X_5158_ _1012_ _1578_ _1686_ _1688_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__o211a_1
X_5089_ _1605_ _1609_ _1616_ _1619_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__or4_1
X_4109_ _0456_ seq.encode.keys_edge_det\[7\] vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _0981_ _0997_ _1023_ _1030_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4391_ _0869_ _0939_ _0943_ _0948_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__o221a_1
X_6130_ _2565_ _2539_ sound3.divisor_m\[16\] _2538_ vssd1 vssd1 vccd1 vccd1 _2566_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _2491_ _2496_ _2479_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__a21o_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _1544_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6963_ sound2.sdiv.A\[26\] _3230_ vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__nor2_1
X_5914_ sound4.count_m\[17\] _2349_ _2322_ sound4.divisor_m\[17\] vssd1 vssd1 vccd1
+ vccd1 _2350_ sky130_fd_sc_hd__a2bb2o_1
X_6894_ sound2.sdiv.A\[26\] sound2.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5845_ _2275_ _2279_ _2282_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__nor3_1
XFILLER_0_75_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5776_ wave_comb.u1.A\[3\] _2224_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7515_ sound3.sdiv.Q\[5\] _3463_ _3437_ sound3.sdiv.Q\[4\] vssd1 vssd1 vccd1 vccd1
+ _0344_ sky130_fd_sc_hd__a22o_1
X_4727_ sound1.count\[10\] sound1.count\[11\] _1281_ vssd1 vssd1 vccd1 vccd1 _1287_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7446_ _3573_ _3581_ _3582_ vssd1 vssd1 vccd1 vccd1 _3603_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4658_ _0981_ _0994_ _0687_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7377_ _3437_ _3540_ _3541_ _3440_ sound3.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _0318_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4589_ _0685_ _0981_ _0939_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__o22a_1
X_6328_ _2756_ _2757_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__xor2_1
X_6259_ sound1.sdiv.Q\[5\] _2690_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3960_ _0622_ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3891_ sound3.sdiv.start vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5630_ sound4.divisor_m\[3\] _2112_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__xnor2_1
X_5561_ _2043_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7300_ _1545_ _3472_ vssd1 vssd1 vccd1 vccd1 _3473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5492_ sound4.count\[15\] _1984_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__and2_2
X_4512_ _0694_ _0996_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_4
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8280_ net122 _0380_ net83 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7231_ sound3.divisor_m\[7\] _1649_ _3419_ vssd1 vssd1 vccd1 vccd1 _3420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4443_ _1013_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4374_ _0686_ _0680_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nor2_4
X_7162_ sound2.sdiv.Q\[18\] _3167_ _3349_ sound2.sdiv.Q\[17\] _3125_ vssd1 vssd1 vccd1
+ vccd1 _0258_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6113_ _2514_ sound3.divisor_m\[6\] sound3.divisor_m\[5\] _2511_ vssd1 vssd1 vccd1
+ vccd1 _2549_ sky130_fd_sc_hd__a22o_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7093_ _3336_ _3343_ _3346_ vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__nand3_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ sound2.count_m\[0\] vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__inv_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7995_ net125 sound1.osc.next_count\[16\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6946_ _3211_ _3214_ vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6877_ _3158_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
X_5828_ _0569_ _2268_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5759_ _2207_ _2212_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7429_ sound3.divisor_m\[18\] _3587_ vssd1 vssd1 vccd1 vccd1 _3588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4090_ seq.player_8.state\[2\] seq.player_8.state\[3\] _0715_ _0716_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_8.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
XFILLER_0_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6800_ sound1.sdiv.Q\[27\] _2894_ _2890_ sound1.sdiv.Q\[26\] vssd1 vssd1 vccd1 vccd1
+ _0168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7780_ net139 _0054_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[9\] sky130_fd_sc_hd__dfrtp_1
X_4992_ sound2.count\[12\] _1527_ _1504_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__o21ai_1
X_6731_ _3081_ _3082_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3943_ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6662_ _3019_ _3021_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3874_ _0512_ _0544_ _0534_ _0545_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__o211a_2
XFILLER_0_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5613_ _2095_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6593_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__nor2_1
X_8332_ net138 _0432_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.C\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5544_ sound4.divisor_m\[5\] sound4.divisor_m\[4\] _2026_ vssd1 vssd1 vccd1 vccd1
+ _2027_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8263_ net140 _0363_ net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5475_ sound4.count\[9\] sound4.count\[10\] _1962_ sound4.count\[11\] vssd1 vssd1
+ vccd1 vccd1 _1975_ sky130_fd_sc_hd__a31o_1
X_8194_ net133 _0315_ net94 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7214_ sound3.divisor_m\[1\] _3408_ _3142_ vssd1 vssd1 vccd1 vccd1 _3409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4426_ net64 _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__nor2_8
X_7145_ sound2.sdiv.Q\[0\] sound2.sdiv.next_dived _2501_ vssd1 vssd1 vccd1 vccd1 _0241_
+ sky130_fd_sc_hd__a21o_1
X_4357_ select1.sequencer_on _0896_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7076_ _3322_ _3325_ _3321_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__a21bo_1
X_4288_ seq.clk_div.count\[21\] _0859_ _0862_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[21\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ sound2.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7978_ net131 sound1.sdiv.next_start net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.start
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6929_ _3187_ _3191_ _3199_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout87 net95 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_6
Xfanout98 net106 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_6
Xfanout76 net3 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__buf_6
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5260_ _0698_ _0605_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__or2_4
XFILLER_0_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4211_ _0789_ seq.clk_div.count\[14\] _0782_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__o21ai_1
X_5191_ sound3.count\[0\] _1721_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[0\]
+ sky130_fd_sc_hd__nand2_1
X_4142_ _0750_ _0749_ _0751_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_4.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_4073_ _0704_ _0707_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__nor2_1
X_7901_ net111 seq.encode.keys_sync\[10\] net72 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7832_ net113 seq.player_1.next_state\[2\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_7763_ net144 pm.next_count\[2\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4975_ _1518_ _1519_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6714_ _3063_ _3065_ _3068_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__a21o_1
X_3926_ _0515_ _0521_ _0519_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__o21ba_1
X_7694_ sound4.sdiv.C\[1\] sound4.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6645_ _3005_ _3006_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3857_ _0525_ _0526_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__nand2_1
X_6576_ _2942_ _2943_ _0866_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ _0468_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_4
X_5527_ _0651_ pm.current_waveform\[4\] vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__and2_1
X_8315_ net124 _0415_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8246_ net141 _0346_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _1961_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
X_8177_ net133 _0298_ net94 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[11\] sky130_fd_sc_hd__dfrtp_2
X_4409_ _0918_ _0909_ _0949_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__or3b_1
X_5389_ _1017_ _1784_ _1781_ _1020_ _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7128_ sound2.sdiv.C\[1\] sound2.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3376_ sky130_fd_sc_hd__or2_1
X_7059_ _3164_ _3316_ _3317_ _3174_ sound2.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 _0224_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4760_ _1311_ vssd1 vssd1 vccd1 vccd1 sound2.sdiv.next_dived sky130_fd_sc_hd__buf_4
XFILLER_0_28_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4691_ sound1.count\[0\] sound1.count\[1\] sound1.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1260_ sky130_fd_sc_hd__a21o_1
X_6430_ sound1.count\[3\] _2201_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6361_ wave_comb.u1.next_start _2789_ _2790_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5312_ _1004_ _1038_ _1786_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8100_ net111 sound2.osc.next_count\[1\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6292_ sound1.sdiv.Q\[6\] _2722_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5243_ sound3.count\[15\] sound3.count\[16\] _1750_ sound3.count\[17\] vssd1 vssd1
+ vccd1 vccd1 _1757_ sky130_fd_sc_hd__a31o_1
X_8031_ net111 _0173_ net72 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[4\] sky130_fd_sc_hd__dfrtp_1
X_5174_ _1591_ _1703_ _1587_ _1704_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__and4_1
X_4125_ seq.player_5.state\[0\] seq.player_5.state\[1\] _0737_ vssd1 vssd1 vccd1 vccd1
+ _0740_ sky130_fd_sc_hd__and3_1
X_4056_ _0682_ _0683_ _0694_ _0697_ vssd1 vssd1 vccd1 vccd1 oct.next_state\[2\] sky130_fd_sc_hd__a211o_1
XFILLER_0_66_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7815_ net114 seq.player_5.next_state\[1\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_5.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7746_ net139 _0031_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4958_ _1507_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3909_ _0575_ net147 vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nor2_8
X_7677_ _2171_ _3732_ _2045_ vssd1 vssd1 vccd1 vccd1 _3733_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4889_ _0696_ _1343_ _1436_ _1439_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6628_ _2989_ _2990_ _0866_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6559_ sound1.divisor_m\[5\] _2928_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8229_ net128 sound3.osc.next_count\[10\] net89 vssd1 vssd1 vccd1 vccd1 sound3.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5930_ sound4.count_m\[15\] _2341_ _2365_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__a21oi_1
X_5861_ _2294_ _2296_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7600_ _2005_ _1018_ _1779_ _3679_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5792_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4812_ _1039_ _1347_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__or2_1
X_7531_ sound3.sdiv.Q\[20\] _3654_ _3643_ sound3.sdiv.Q\[19\] _3399_ vssd1 vssd1 vccd1
+ vccd1 _0359_ sky130_fd_sc_hd__a221o_1
X_4743_ sound1.count\[15\] _1296_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7462_ _2863_ _0563_ _3616_ vssd1 vssd1 vccd1 vccd1 _3617_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4674_ _1018_ _0959_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__or2_2
X_6413_ _0811_ _2829_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__nor2_1
X_7393_ _3551_ _3554_ vssd1 vssd1 vccd1 vccd1 _3556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6344_ sound4.sdiv.Q\[7\] _0576_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__nand2_1
X_6275_ _2289_ _2705_ _2706_ _2290_ sound4.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 _2707_
+ sky130_fd_sc_hd__a32o_1
X_5226_ _1744_ _1745_ _1721_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__and3b_1
X_8014_ net127 _0156_ net88 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5157_ _1053_ _1572_ _1550_ _1125_ _1687_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__o221a_1
X_5088_ sound3.count\[18\] _1618_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__xnor2_1
X_4108_ _0726_ _0725_ _0728_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_7.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4039_ _0674_ _0678_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__nor2_8
XFILLER_0_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ net120 _0014_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4390_ _0950_ _0954_ _0958_ _0960_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _2493_ _2495_ _2459_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__o21ai_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5011_ _1504_ _1542_ _1543_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__and3_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6962_ sound2.divisor_m\[7\] _3221_ vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5913_ sound4.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__inv_2
X_6893_ _3164_ _3165_ _3166_ _3168_ sound2.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _0207_
+ sky130_fd_sc_hd__a32o_1
X_5844_ _2276_ _2277_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7514_ sound3.sdiv.Q\[4\] _3463_ _3437_ sound3.sdiv.Q\[3\] vssd1 vssd1 vccd1 vccd1
+ _0343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5775_ wave_comb.u1.A\[3\] _0573_ wave_comb.u1.next_dived _2226_ vssd1 vssd1 vccd1
+ vccd1 _0031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4726_ _1286_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7445_ _3564_ _3568_ _3575_ _3583_ _3601_ vssd1 vssd1 vccd1 vccd1 _3602_ sky130_fd_sc_hd__a2111o_1
X_4657_ _1220_ _1221_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7376_ _3529_ _3532_ _3539_ vssd1 vssd1 vccd1 vccd1 _3541_ sky130_fd_sc_hd__o21bai_1
X_6327_ sound2.sdiv.Q\[7\] _0578_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__nand2_1
X_4588_ _1100_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ sound1.sdiv.Q\[4\] _2656_ _2657_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__a21bo_1
X_6189_ _2279_ _2620_ _2622_ _2292_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__o22a_1
X_5209_ _1734_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3890_ _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5560_ sound4.sdiv.A\[22\] _2038_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__xor2_2
XFILLER_0_53_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4511_ _0680_ _0976_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5491_ _1987_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7230_ _2863_ vssd1 vssd1 vccd1 vccd1 _3419_ sky130_fd_sc_hd__buf_8
X_4442_ _0944_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7161_ sound2.sdiv.Q\[17\] _3167_ _3349_ sound2.sdiv.Q\[16\] _3124_ vssd1 vssd1 vccd1
+ vccd1 _0257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4373_ _0674_ _0677_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__nor2_8
XFILLER_0_111_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6112_ _2547_ sound3.divisor_m\[8\] _2513_ sound3.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2548_ sky130_fd_sc_hd__a22o_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _3336_ _3343_ _3346_ vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__a21o_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ sound2.count_m\[16\] _2471_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__and2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7994_ net125 sound1.osc.next_count\[15\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _3211_ _3214_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6876_ sound2.divisor_m\[13\] _3157_ _3142_ vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5827_ _0571_ _2267_ wave_comb.u1.C\[3\] vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5758_ wave_comb.u1.A\[0\] _2211_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__xnor2_1
X_4709_ _1272_ _1273_ _1256_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__and3b_1
XFILLER_0_17_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7428_ sound3.divisor_m\[17\] _3578_ _3448_ vssd1 vssd1 vccd1 vccd1 _3587_ sky130_fd_sc_hd__o21a_1
X_5689_ sound4.sdiv.A\[23\] _2038_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7359_ sound3.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _3525_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6730_ sound1.sdiv.A\[21\] _3055_ _3079_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4991_ sound2.count\[12\] _1527_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__and2_1
X_3942_ _0587_ _0606_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__nand2_8
XFILLER_0_46_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6661_ sound1.divisor_m\[15\] _3020_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__xnor2_1
X_3873_ _0520_ _0524_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__nand2_1
X_6592_ sound1.divisor_m\[8\] _2958_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__xnor2_1
X_5612_ sound4.divisor_m\[6\] _2094_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8331_ net124 _0431_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[26\] sky130_fd_sc_hd__dfrtp_4
X_5543_ sound4.divisor_m\[3\] sound4.divisor_m\[2\] sound4.divisor_m\[1\] sound4.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8262_ net140 _0362_ net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[23\] sky130_fd_sc_hd__dfrtp_1
X_5474_ _1973_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__inv_2
X_8193_ net133 _0314_ net94 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7213_ _1673_ vssd1 vssd1 vccd1 vccd1 _3408_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4425_ _0995_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__buf_8
X_7144_ sound2.sdiv.next_dived _3386_ _2276_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4356_ seq.player_7.state\[3\] _0897_ _0901_ seq.player_8.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _0927_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7075_ _3330_ _3331_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__or2b_1
X_4287_ seq.clk_div.count\[21\] _0859_ _0813_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__o21ai_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ sound2.count_m\[7\] _2460_ _2461_ sound2.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2462_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7977_ net131 _0140_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6928_ _3187_ _3191_ _3199_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6859_ _3146_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout88 net95 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_6
Xfanout99 net106 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_4
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout77 net80 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_8
XFILLER_0_36_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4210_ seq.clk_div.count\[10\] _0779_ _0777_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5190_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4141_ seq.player_4.state\[2\] _0748_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__xor2_1
X_4072_ _0701_ _0707_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__nor2_1
XFILLER_0_92_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7900_ net107 inputcont.INTERNAL_SYNCED_I\[7\] net68 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7831_ net113 seq.player_1.next_state\[1\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_7762_ net144 pm.next_count\[1\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4974_ sound2.count\[6\] _1515_ _1504_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__o21ai_1
X_6713_ _3066_ _3067_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7693_ _3743_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3925_ _0548_ _0543_ _0582_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nand3_2
XFILLER_0_46_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6644_ _3001_ _3004_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3856_ inputcont.INTERNAL_SYNCED_I\[3\] _0502_ _0512_ vssd1 vssd1 vccd1 vccd1 _0530_
+ sky130_fd_sc_hd__a21oi_1
X_6575_ _2942_ _2943_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3787_ _0462_ _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or2_1
X_5526_ _2009_ pm.current_waveform\[5\] vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and2_1
X_8314_ net124 _0414_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[9\] sky130_fd_sc_hd__dfrtp_1
X_8245_ net141 _0345_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[6\] sky130_fd_sc_hd__dfrtp_2
X_5457_ _1779_ _1936_ _1959_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4408_ _0978_ _0971_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__or2_4
X_8176_ net133 _0297_ net94 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5388_ _1025_ _1794_ _1796_ _1027_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__o221a_1
X_4339_ seq.player_7.state\[0\] _0898_ _0901_ seq.player_8.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _0910_ sky130_fd_sc_hd__a22o_1
X_7127_ sound2.sdiv.C\[1\] sound2.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3375_ sky130_fd_sc_hd__nand2_1
X_7058_ _3302_ _3306_ _3315_ vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6009_ sound2.count_m\[10\] _2443_ _2444_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4690_ _1259_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6360_ wave_comb.u1.Q\[8\] _0572_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5311_ _1811_ _1812_ _1818_ _1821_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__a211o_1
X_6291_ sound1.sdiv.Q\[5\] _2656_ _2690_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__a21o_1
X_8030_ net111 _0172_ net72 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[3\] sky130_fd_sc_hd__dfrtp_1
X_5242_ sound3.count\[16\] sound3.count\[17\] _1753_ vssd1 vssd1 vccd1 vccd1 _1756_
+ sky130_fd_sc_hd__and3_1
X_5173_ _1025_ _1046_ _1559_ _1578_ _1165_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__o32a_1
X_4124_ seq.player_5.state\[0\] _0737_ _0739_ vssd1 vssd1 vccd1 vccd1 seq.player_5.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
Xinput1 cs vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_8
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4055_ _0682_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7814_ net114 seq.player_5.next_state\[0\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_5.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7745_ net139 _0030_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[2\] sky130_fd_sc_hd__dfrtp_1
X_4957_ _1504_ _1505_ _1506_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3908_ _0576_ vssd1 vssd1 vccd1 vccd1 sound4.sdiv.next_start sky130_fd_sc_hd__inv_2
X_7676_ _2042_ _2168_ vssd1 vssd1 vccd1 vccd1 _3732_ sky130_fd_sc_hd__or2b_1
X_4888_ _1123_ _1339_ _1336_ _1141_ _1438_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6627_ _2989_ _2990_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3839_ _0480_ _0481_ _0482_ net67 vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6558_ sound1.divisor_m\[4\] _2919_ _2903_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6489_ sound1.divisor_m\[9\] _2005_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__nor2_1
X_5509_ rate_clk.count\[0\] vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8228_ net128 sound3.osc.next_count\[9\] net89 vssd1 vssd1 vccd1 vccd1 sound3.count\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8159_ net132 _0280_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5860_ _2294_ _2296_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _1015_ _1323_ _1327_ _0946_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__o221a_1
X_5791_ wave_comb.u1.A\[4\] wave_comb.u1.A\[3\] _2224_ vssd1 vssd1 vccd1 vccd1 _2240_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7530_ sound3.sdiv.Q\[19\] _3654_ _3643_ sound3.sdiv.Q\[18\] _3398_ vssd1 vssd1 vccd1
+ vccd1 _0358_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4742_ _1298_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_7461_ _3613_ _3614_ _3612_ vssd1 vssd1 vccd1 vccd1 _3616_ sky130_fd_sc_hd__a21oi_1
X_4673_ _0985_ _0939_ _1242_ _0950_ _1243_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6412_ _0719_ seq.encode.play vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__nand2_1
X_7392_ _3551_ _3554_ vssd1 vssd1 vccd1 vccd1 _3555_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6343_ net31 net30 vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__and2b_1
X_6274_ sound4.sdiv.Q\[5\] _2704_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5225_ sound3.count\[9\] sound3.count\[10\] _1738_ sound3.count\[11\] vssd1 vssd1
+ vccd1 vccd1 _1745_ sky130_fd_sc_hd__a31o_1
X_8013_ net127 _0155_ net88 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5156_ _0983_ _1580_ _1565_ _1146_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ _0695_ _1617_ _1591_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__o21a_1
X_4107_ seq.player_7.state\[1\] seq.player_7.state\[2\] _0722_ seq.player_7.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4038_ inputcont.u2.next_in inputcont.INTERNAL_OCTAVE_INPUT vssd1 vssd1 vccd1 vccd1
+ _0682_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5989_ _2384_ _2424_ _2377_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__a21o_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7728_ net120 _0013_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7659_ _3719_ _2154_ vssd1 vssd1 vccd1 vccd1 _3721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap63 _1040_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_8
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ sound2.count\[18\] _1539_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__nand2_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6961_ sound2.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5912_ sound4.divisor_m\[3\] sound4.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__or2b_1
X_6892_ _3167_ vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5843_ sound2.sdiv.Q\[0\] _0578_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7513_ sound3.sdiv.Q\[3\] _3463_ sound3.sdiv.next_dived sound3.sdiv.Q\[2\] vssd1
+ vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5774_ _2222_ _2225_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4725_ _1256_ _1284_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__and3_1
X_7444_ _3600_ vssd1 vssd1 vccd1 vccd1 _3601_ sky130_fd_sc_hd__inv_2
X_4656_ sound1.count\[11\] _1050_ _1224_ _1226_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__o211a_1
X_7375_ _3529_ _3532_ _3539_ vssd1 vssd1 vccd1 vccd1 _3540_ sky130_fd_sc_hd__or3b_1
X_4587_ _0685_ _0982_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__nor2_4
XFILLER_0_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6326_ sound2.sdiv.Q\[6\] _2660_ _2718_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__a21oi_1
X_6257_ _2687_ _2688_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__nand2_1
X_6188_ _2586_ _2621_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__xor2_1
X_5208_ _1732_ _1733_ _1721_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__and3b_1
X_5139_ _0869_ _1567_ _1550_ _0954_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4510_ _0990_ _0960_ _0994_ _1039_ _1080_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5490_ _1779_ _1936_ _1985_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4441_ _0675_ _0970_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__nor2_4
XFILLER_0_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7160_ sound2.sdiv.Q\[16\] _3167_ _3349_ sound2.sdiv.Q\[15\] _3123_ vssd1 vssd1 vccd1
+ vccd1 _0256_ sky130_fd_sc_hd__a221o_1
X_6111_ sound3.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__inv_2
X_4372_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__buf_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _3345_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ sound2.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__inv_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7993_ net125 sound1.osc.next_count\[14\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6944_ sound2.divisor_m\[6\] _3213_ vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875_ _1434_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5826_ _0646_ _2266_ _2267_ _0573_ wave_comb.u1.C\[2\] vssd1 vssd1 vccd1 vccd1 _0041_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5757_ wave_comb.u1.M\[1\] _2210_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4708_ sound1.count\[6\] _1269_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7427_ sound3.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 _3586_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5688_ sound4.sdiv.A\[20\] sound4.sdiv.A\[19\] _2038_ vssd1 vssd1 vccd1 vccd1 _2171_
+ sky130_fd_sc_hd__o21ai_4
X_4639_ _0949_ _0988_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7358_ _3437_ _3523_ _3524_ _3440_ sound3.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _0316_
+ sky130_fd_sc_hd__a32o_1
X_7289_ _0577_ vssd1 vssd1 vccd1 vccd1 _3463_ sky130_fd_sc_hd__clkbuf_8
X_6309_ _2735_ _2739_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4990_ _1529_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3941_ _0588_ _0589_ _0598_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__o31a_2
X_6660_ sound1.divisor_m\[14\] _3011_ _2903_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3872_ inputcont.INTERNAL_SYNCED_I\[3\] _0502_ _0543_ vssd1 vssd1 vccd1 vccd1 _0544_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6591_ sound1.sdiv.A\[26\] _2957_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__nor2_1
X_5611_ _2036_ _2027_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5542_ pm.current_waveform\[8\] _2024_ _2025_ vssd1 vssd1 vccd1 vccd1 pm.next_pwm_o
+ sky130_fd_sc_hd__o21a_1
X_8330_ net124 _0430_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8261_ net140 _0361_ net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[22\] sky130_fd_sc_hd__dfrtp_1
X_5473_ sound4.count\[10\] sound4.count\[11\] _1966_ vssd1 vssd1 vccd1 vccd1 _1973_
+ sky130_fd_sc_hd__and3_1
X_8192_ net142 _0313_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7212_ _3407_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4424_ _0686_ _0674_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nor2_1
X_4355_ net37 _0925_ _0698_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__mux2_2
X_7143_ _3373_ _3385_ vssd1 vssd1 vccd1 vccd1 _3386_ sky130_fd_sc_hd__nand2_1
X_7074_ sound2.sdiv.A\[18\] _3329_ vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__nand2_1
X_4286_ _0861_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[20\] sky130_fd_sc_hd__clkbuf_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ sound2.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7976_ net131 _0139_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6927_ _3197_ _3198_ vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6858_ sound2.divisor_m\[7\] _3145_ _3142_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout89 net90 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__buf_6
X_5809_ wave_comb.u1.A\[8\] _2224_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout78 net80 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_8
X_6789_ sound1.sdiv.Q\[16\] _2893_ _0867_ sound1.sdiv.Q\[15\] _2846_ vssd1 vssd1 vccd1
+ vccd1 _0157_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4140_ seq.player_4.state\[2\] seq.player_4.state\[3\] vssd1 vssd1 vccd1 vccd1 _0750_
+ sky130_fd_sc_hd__nand2_1
X_4071_ seq.beat\[3\] net52 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nand2_8
XFILLER_0_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7830_ net113 seq.player_1.next_state\[0\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7761_ net144 pm.next_count\[0\] net105 vssd1 vssd1 vccd1 vccd1 pm.count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4973_ sound2.count\[6\] _1515_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6712_ sound1.sdiv.A\[19\] _3055_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7692_ _1764_ _2182_ sound4.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3924_ _0584_ _0585_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6643_ _3001_ _3004_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3855_ _0513_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6574_ _2932_ _2933_ _2930_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3786_ inputcont.INTERNAL_SYNCED_I\[8\] _0448_ _0455_ _0466_ vssd1 vssd1 vccd1 vccd1
+ _0467_ sky130_fd_sc_hd__a211o_1
X_5525_ pm.count\[5\] vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8313_ net122 _0413_ net83 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[8\] sky130_fd_sc_hd__dfrtp_1
X_8244_ net141 _0344_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ sound4.count\[7\] _1955_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4407_ _0685_ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__nor2_4
X_8175_ net133 _0296_ net94 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5387_ _1024_ _1028_ _1786_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__or3_1
X_4338_ net36 _0908_ _0698_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__mux2_4
X_7126_ _3374_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_7057_ _3302_ _3306_ _3315_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__o21ai_1
X_4269_ _0849_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
X_6008_ sound2.divisor_m\[10\] sound2.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2444_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ net130 _0122_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6290_ _2289_ _2719_ _2720_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5310_ sound4.count\[16\] _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5241_ sound3.count\[16\] _1753_ _1755_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[16\]
+ sky130_fd_sc_hd__a21oi_1
X_5172_ _1159_ _1567_ _1565_ _0997_ _1702_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__o221a_1
X_4123_ seq.player_5.state\[1\] seq.player_5.state\[2\] seq.player_5.state\[3\] _0738_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a311o_1
X_4054_ _0695_ _0687_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__nand2_4
Xinput2 hwclk vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7813_ net107 seq.player_6.next_state\[3\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_6.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_7744_ net137 _0029_ net98 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ sound2.count\[0\] sound2.count\[1\] vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3907_ _0575_ _0556_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__nor2_4
X_7675_ sound4.sdiv.A\[21\] _2184_ _3681_ _3731_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__a22o_1
X_4887_ _1138_ _1323_ _1341_ _1126_ _1437_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6626_ _2970_ _2980_ _2976_ _2979_ _2974_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__o32a_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3838_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6557_ sound1.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5508_ _2000_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3769_ inputcont.INTERNAL_SYNCED_I\[5\] _0443_ inputcont.INTERNAL_SYNCED_I\[4\] inputcont.INTERNAL_SYNCED_I\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__or4b_2
X_6488_ _2873_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8227_ net129 sound3.osc.next_count\[8\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_5439_ _1779_ _1936_ _1945_ _1946_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__and4_1
X_8158_ net132 _0279_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[11\] sky130_fd_sc_hd__dfrtp_1
X_7109_ _3346_ _3350_ _3355_ vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__or3b_1
X_8089_ net118 _0231_ net79 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4810_ _0684_ _1077_ _1343_ _1338_ _0971_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__o32a_1
X_5790_ _2237_ _2238_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4741_ _1296_ _1297_ _1256_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__and3b_1
X_7460_ _3612_ _3613_ _3614_ vssd1 vssd1 vccd1 vccd1 _3615_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4672_ _0958_ _0944_ _1004_ _1025_ _0981_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__o32a_1
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6411_ _2828_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7391_ sound3.divisor_m\[14\] _3553_ vssd1 vssd1 vccd1 vccd1 _3554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6342_ _2766_ _2771_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6273_ sound4.sdiv.Q\[5\] _0576_ _2704_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__a21o_1
X_5224_ sound3.count\[10\] sound3.count\[11\] _1741_ vssd1 vssd1 vccd1 vccd1 _1744_
+ sky130_fd_sc_hd__and3_1
X_8012_ net127 _0154_ net88 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[13\] sky130_fd_sc_hd__dfrtp_1
X_5155_ _1134_ _1567_ _1570_ _1154_ _1685_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5086_ net64 _1603_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__nand2_1
X_4106_ _0726_ _0725_ _0727_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_7.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_4037_ _0676_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nor2_4
XFILLER_0_94_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _2387_ _2423_ _2386_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__a21bo_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7727_ net121 _0012_ net82 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4939_ _1189_ _1327_ _1365_ _0959_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7658_ _3719_ _2154_ vssd1 vssd1 vccd1 vccd1 _3720_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6609_ _0866_ _2972_ _2973_ sound1.sdiv.next_start _2974_ vssd1 vssd1 vccd1 vccd1
+ _0117_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7589_ sound4.divisor_m\[13\] _1875_ _2186_ vssd1 vssd1 vccd1 vccd1 _3673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap53 net54 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xmax_cap64 _0684_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_6
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6960_ _3164_ _3227_ _3228_ _3174_ sound2.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 _0214_
+ sky130_fd_sc_hd__a32o_1
X_5911_ _2316_ sound4.divisor_m\[7\] _2318_ sound4.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2347_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6891_ _0578_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__buf_6
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5842_ _2279_ _2277_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5773_ wave_comb.u1.A\[2\] _2224_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7512_ sound3.sdiv.Q\[2\] _3463_ sound3.sdiv.next_dived sound3.sdiv.Q\[1\] vssd1
+ vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ sound1.count\[10\] _1281_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7443_ _3591_ _3596_ vssd1 vssd1 vccd1 vccd1 _3600_ sky130_fd_sc_hd__nor2_1
X_4655_ sound1.count\[17\] _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__xnor2_1
X_7374_ _3537_ _3538_ vssd1 vssd1 vccd1 vccd1 _3539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4586_ _1150_ _1153_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__and3_2
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6325_ _2292_ _2751_ _2754_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6256_ sound2.sdiv.Q\[5\] _2686_ _2292_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__a21oi_1
X_6187_ sound1.sdiv.Q\[0\] sound1.sdiv.Q\[1\] sound1.sdiv.Q\[2\] _0579_ _2434_ vssd1
+ vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__o311a_1
X_5207_ sound3.count\[4\] _1728_ sound3.count\[5\] vssd1 vssd1 vccd1 vccd1 _1733_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5138_ _0959_ _0993_ _1580_ _1562_ _0985_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__o32a_1
X_5069_ _1126_ _1580_ _1598_ _1599_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ _0695_ _0678_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__or2_4
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6110_ sound3.count_m\[17\] _2543_ _2545_ sound3.divisor_m\[17\] vssd1 vssd1 vccd1
+ vccd1 _2546_ sky130_fd_sc_hd__a2bb2o_1
X_4371_ _0940_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ sound2.sdiv.A\[20\] _3329_ vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__xor2_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ sound2.count_m\[17\] _2470_ sound2.count_m\[18\] vssd1 vssd1 vccd1 vccd1 _2477_
+ sky130_fd_sc_hd__a21o_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7992_ net125 sound1.osc.next_count\[13\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6943_ _3177_ _3212_ vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6874_ _3156_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5825_ wave_comb.u1.C\[2\] wave_comb.u1.C\[0\] wave_comb.u1.C\[1\] vssd1 vssd1 vccd1
+ vccd1 _2267_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5756_ wave_comb.u1.M\[0\] _2209_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4707_ sound1.count\[6\] _1269_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__and2_1
X_5687_ sound4.sdiv.A\[22\] sound4.sdiv.A\[21\] _2038_ vssd1 vssd1 vccd1 vccd1 _2170_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7426_ sound3.sdiv.A\[17\] _3463_ sound3.sdiv.next_dived _3585_ vssd1 vssd1 vccd1
+ vccd1 _0323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4638_ sound1.count\[3\] _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__xnor2_1
X_7357_ _3503_ _3507_ _3521_ _3511_ _3520_ vssd1 vssd1 vccd1 vccd1 _3524_ sky130_fd_sc_hd__a311o_1
XFILLER_0_102_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4569_ _0945_ _1038_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__nor2_4
X_7288_ _3454_ _3452_ _3460_ _0563_ _2005_ vssd1 vssd1 vccd1 vccd1 _3462_ sky130_fd_sc_hd__a311o_1
X_6308_ _2289_ _2737_ _2738_ _2290_ sound4.sdiv.Q\[7\] vssd1 vssd1 vccd1 vccd1 _2739_
+ sky130_fd_sc_hd__a32o_1
X_6239_ _2668_ _2671_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3940_ _0603_ _0595_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__or3b_2
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3871_ _0513_ _0531_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6590_ sound1.divisor_m\[7\] _2948_ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__nor2_1
X_5610_ sound4.sdiv.A\[6\] _2092_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5541_ pm.current_waveform\[8\] _2024_ pm.count\[8\] vssd1 vssd1 vccd1 vccd1 _2025_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8260_ net132 _0360_ net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7211_ sound3.divisor_m\[0\] _1583_ _3142_ vssd1 vssd1 vccd1 vccd1 _3407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5472_ _1972_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
X_8191_ net142 _0312_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4423_ _0949_ _0909_ _0918_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nand3_4
X_4354_ seq.player_1.state\[2\] _0871_ _0873_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_
+ sky130_fd_sc_hd__a22o_1
X_7142_ sound2.sdiv.A\[25\] _3327_ _3177_ vssd1 vssd1 vccd1 vccd1 _3385_ sky130_fd_sc_hd__o21ai_1
X_7073_ sound2.sdiv.A\[18\] _3329_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__nor2_1
X_4285_ _0859_ _0813_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__and3b_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ sound2.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__inv_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7975_ net131 _0138_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _3193_ _3196_ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6857_ _1368_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5808_ wave_comb.u1.A\[8\] _2224_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6788_ sound1.sdiv.Q\[15\] _2893_ _0867_ sound1.sdiv.Q\[14\] _2845_ vssd1 vssd1 vccd1
+ vccd1 _0156_ sky130_fd_sc_hd__a221o_1
Xfanout68 net76 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_8
Xfanout79 net80 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_8
XFILLER_0_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5739_ sound4.sdiv.Q\[21\] _2182_ _2185_ sound4.sdiv.Q\[20\] _2200_ vssd1 vssd1 vccd1
+ vccd1 _0021_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7409_ sound3.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _3570_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4070_ _0703_ _0706_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__nor2_2
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7760_ net143 wave_comb.u1.next_start net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.start
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4972_ _1517_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6711_ sound1.sdiv.A\[19\] _3055_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7691_ _3681_ _2179_ _3742_ _2184_ sound4.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _0431_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3923_ _0581_ _0583_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6642_ sound1.divisor_m\[13\] _3003_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3854_ _0515_ _0518_ _0521_ _0523_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__o41a_1
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6573_ _2940_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__nand2_1
X_8312_ net123 _0412_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3785_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
X_5524_ _2007_ pm.current_waveform\[6\] vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8243_ net141 _0343_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[4\] sky130_fd_sc_hd__dfrtp_1
X_5455_ sound4.count\[7\] _1955_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__nand2_1
X_8174_ net132 _0295_ net93 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4406_ _0678_ _0964_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__nand2_8
X_7125_ _1311_ _3167_ sound2.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3374_ sky130_fd_sc_hd__mux2_1
X_5386_ _1892_ _1893_ _1896_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__and3_2
X_4337_ seq.player_1.state\[1\] _0871_ _0873_ _0907_ vssd1 vssd1 vccd1 vccd1 _0908_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7056_ _3313_ _3314_ vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__nor2_1
X_4268_ _0847_ _0813_ _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__and3b_1
X_6007_ sound2.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__inv_2
X_4199_ seq.tempo_select.state\[1\] _0791_ _0792_ seq.clk_div.count\[12\] vssd1 vssd1
+ vccd1 vccd1 _0793_ sky130_fd_sc_hd__o22a_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ net130 _0121_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7889_ net113 seq.encode.next_sequencer_on net74 vssd1 vssd1 vccd1 vccd1 select1.sequencer_on
+ sky130_fd_sc_hd__dfrtp_4
X_6909_ _3164_ _3181_ _3182_ _3174_ sound2.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _0209_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_92_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5240_ sound3.count\[16\] _1753_ _1721_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5171_ _1004_ _1038_ _1553_ _1580_ _1166_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__o32a_1
X_4122_ seq.player_5.state\[0\] _0737_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__and2_1
X_4053_ _0674_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__buf_12
Xinput3 n_rst vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_6
XFILLER_0_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7812_ net107 seq.player_6.next_state\[2\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_6.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_7743_ net137 _0028_ net98 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[0\] sky130_fd_sc_hd__dfrtp_1
X_4955_ sound2.count\[0\] sound2.count\[1\] vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3906_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7674_ _2040_ _3730_ vssd1 vssd1 vccd1 vccd1 _3731_ sky130_fd_sc_hd__xor2_1
X_4886_ _1129_ _1347_ _1345_ _1140_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6625_ _2987_ _2988_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3837_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__and3_1
X_6556_ sound1.sdiv.A\[4\] _2895_ sound1.sdiv.next_dived _2926_ vssd1 vssd1 vccd1
+ vccd1 _0112_ sky130_fd_sc_hd__a22o_1
X_3768_ inputcont.INTERNAL_SYNCED_I\[8\] _0448_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_
+ sky130_fd_sc_hd__a21oi_1
X_5507_ _1779_ _1998_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6487_ sound1.divisor_m\[8\] _2872_ _2864_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__mux2_1
X_8226_ net128 sound3.osc.next_count\[7\] net89 vssd1 vssd1 vccd1 vccd1 sound3.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5438_ sound4.count\[3\] _1940_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__or2_1
X_8157_ net132 _0278_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5369_ _1064_ _1781_ _1878_ _1879_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7108_ _3358_ _3359_ vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__nand2_1
X_8088_ net118 _0230_ net79 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[23\] sky130_fd_sc_hd__dfrtp_1
X_7039_ sound2.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ sound1.count\[12\] sound1.count\[13\] _1287_ sound1.count\[14\] vssd1 vssd1
+ vccd1 vccd1 _1297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4671_ _1012_ _1028_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__nor2_1
X_7390_ _3448_ _3552_ vssd1 vssd1 vccd1 vccd1 _3553_ sky130_fd_sc_hd__and2_1
X_6410_ pm.current_waveform\[8\] _2827_ _2808_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6341_ _2289_ _2769_ _2770_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6272_ sound4.sdiv.Q\[4\] _2641_ _2673_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5223_ sound3.count\[10\] _1741_ _1743_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[10\]
+ sky130_fd_sc_hd__a21oi_1
X_8011_ net127 _0153_ net88 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[12\] sky130_fd_sc_hd__dfrtp_1
X_5154_ _1151_ _1562_ _1574_ _1042_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__o22a_1
X_4105_ seq.player_7.state\[2\] _0724_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__xor2_1
X_5085_ sound3.count\[15\] _1615_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4036_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__inv_8
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ sound1.count_m\[10\] _2378_ _2390_ _2391_ _2379_ vssd1 vssd1 vccd1 vccd1 _2423_
+ sky130_fd_sc_hd__a221o_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7726_ net121 _0011_ net82 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[11\] sky130_fd_sc_hd__dfrtp_1
X_4938_ _1077_ _1323_ _1339_ _1193_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4869_ _0964_ _1418_ _1419_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__or3b_1
X_7657_ _2145_ _2150_ _3715_ _2147_ vssd1 vssd1 vccd1 vccd1 _3719_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6608_ sound1.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7588_ _3672_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6539_ sound1.divisor_m\[2\] sound1.divisor_m\[1\] sound1.divisor_m\[0\] _2903_ vssd1
+ vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8209_ net144 _0330_ net105 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[24\] sky130_fd_sc_hd__dfrtp_1
Xmax_cap65 _0565_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ sound4.divisor_m\[1\] vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__inv_2
X_6890_ sound2.divisor_m\[0\] sound2.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5841_ _2278_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5772_ _2223_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__buf_4
X_7511_ sound3.sdiv.Q\[1\] _3463_ sound3.sdiv.next_dived sound3.sdiv.Q\[0\] vssd1
+ vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__a22o_1
X_4723_ sound1.count\[10\] _1281_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7442_ sound3.sdiv.A\[19\] _3595_ vssd1 vssd1 vccd1 vccd1 _3599_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4654_ _0988_ _0955_ _0971_ _1069_ _1018_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7373_ _3534_ _3536_ vssd1 vssd1 vccd1 vccd1 _3538_ sky130_fd_sc_hd__nand2_1
X_4585_ _0967_ _1095_ _1042_ _0976_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6324_ sound1.sdiv.Q\[8\] _2293_ _2752_ _2753_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__o2bb2a_1
X_6255_ sound2.sdiv.Q\[5\] _0578_ _2686_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__a21o_1
X_5206_ sound3.count\[4\] sound3.count\[5\] _1728_ vssd1 vssd1 vccd1 vccd1 _1732_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_110_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6186_ sound1.sdiv.Q\[4\] _0579_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__nand2_1
X_5137_ _0978_ _0944_ _1565_ _1572_ _0997_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__o32a_1
XFILLER_0_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5068_ _1123_ _1559_ _1565_ _1127_ _1591_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__o221a_1
X_4019_ _0587_ _0597_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7709_ wave_comb.u1.M\[0\] net32 _0645_ vssd1 vssd1 vccd1 vccd1 _3754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _0937_ _0909_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _2474_ sound2.divisor_m\[4\] _2475_ sound2.divisor_m\[3\] vssd1 vssd1 vccd1
+ vccd1 _2476_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7991_ net125 sound1.osc.next_count\[12\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ sound2.divisor_m\[5\] sound2.divisor_m\[4\] _3194_ vssd1 vssd1 vccd1 vccd1
+ _3212_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6873_ sound2.divisor_m\[12\] _3155_ _3142_ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5824_ wave_comb.u1.C\[0\] wave_comb.u1.C\[1\] wave_comb.u1.C\[2\] vssd1 vssd1 vccd1
+ vccd1 _2266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5755_ wave_comb.u1.A\[10\] vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4706_ _1271_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
X_5686_ _2042_ _2044_ _2045_ _2168_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__or4b_2
X_7425_ _3583_ _3584_ vssd1 vssd1 vccd1 vccd1 _3585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4637_ _0981_ _1198_ _0992_ _1199_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__o221a_2
XFILLER_0_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7356_ _3520_ _3522_ vssd1 vssd1 vccd1 vccd1 _3523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4568_ _0959_ _1028_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nor2_4
X_7287_ _3454_ _3452_ _3460_ vssd1 vssd1 vccd1 vccd1 _3461_ sky130_fd_sc_hd__a21oi_1
X_6307_ sound4.sdiv.Q\[6\] _2736_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__nand2_1
X_4499_ _0988_ _0955_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__a21o_4
XFILLER_0_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6238_ sound3.sdiv.Q\[5\] _2301_ _2670_ _2292_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__o2bb2a_1
X_6169_ sound3.sdiv.Q\[2\] _2602_ _2292_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__a21o_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3870_ _0542_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__inv_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5540_ _0657_ pm.current_waveform\[7\] _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5471_ _1779_ _1936_ _1970_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7210_ sound3.count_m\[18\] _3403_ _3406_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4422_ _0674_ _0680_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nor2_4
X_8190_ net142 _0311_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4353_ seq.player_2.state\[2\] _0876_ _0878_ _0923_ vssd1 vssd1 vccd1 vccd1 _0924_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7141_ _3384_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
X_4284_ _0791_ _0858_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nand2_1
X_7072_ _3328_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__buf_4
X_6023_ _2442_ _2445_ _2453_ _2458_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__and4bb_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7974_ net131 _0137_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[2\] sky130_fd_sc_hd__dfrtp_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6925_ _3193_ _3196_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6856_ _3144_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
X_3999_ pm.count\[6\] _0652_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__and2_1
X_5807_ wave_comb.u1.A\[8\] _0573_ wave_comb.u1.next_dived _2253_ vssd1 vssd1 vccd1
+ vccd1 _0036_ sky130_fd_sc_hd__a22o_1
X_6787_ sound1.sdiv.Q\[14\] _2893_ _0867_ sound1.sdiv.Q\[13\] _2844_ vssd1 vssd1 vccd1
+ vccd1 _0155_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout69 net76 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_8
XFILLER_0_17_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5738_ sound4.count\[13\] _2186_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5669_ _2057_ _2061_ _2141_ _2148_ _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__a41o_1
X_7408_ _3564_ _3568_ vssd1 vssd1 vccd1 vccd1 _3569_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7339_ _3437_ _3506_ _3507_ _3440_ sound3.sdiv.A\[8\] vssd1 vssd1 vccd1 vccd1 _0314_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4971_ _1515_ _1516_ _1504_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__and3b_1
X_6710_ _3022_ _3026_ _3033_ _3042_ _3064_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_74_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7690_ _2178_ _2175_ _2176_ vssd1 vssd1 vccd1 vccd1 _3742_ sky130_fd_sc_hd__nand3_1
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3922_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6641_ _2903_ _3002_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3853_ _0514_ _0525_ _0526_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6572_ _2936_ _2939_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3784_ inputcont.INTERNAL_SYNCED_I\[6\] _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__or4b_1
X_8311_ net123 _0411_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[6\] sky130_fd_sc_hd__dfrtp_1
X_5523_ pm.count\[6\] vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8242_ net143 _0342_ net104 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[3\] sky130_fd_sc_hd__dfrtp_2
X_5454_ _1958_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_8173_ net132 _0294_ net93 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[7\] sky130_fd_sc_hd__dfrtp_4
X_4405_ _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5385_ _0960_ _1777_ _1894_ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4336_ seq.player_2.state\[1\] _0876_ _0878_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7124_ _3349_ _3371_ _3373_ _3174_ sound2.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _0233_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7055_ sound2.sdiv.A\[16\] _3311_ vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__nor2_1
X_4267_ seq.clk_div.count\[15\] _0844_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__or2_1
X_4198_ seq.tempo_select.state\[1\] seq.clk_div.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0792_ sky130_fd_sc_hd__nand2_1
X_6006_ sound2.count_m\[14\] _2440_ sound2.count_m\[13\] _2441_ vssd1 vssd1 vccd1
+ vccd1 _2442_ sky130_fd_sc_hd__a22o_1
X_7957_ net130 _0120_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7888_ net111 tempo_select_on net72 vssd1 vssd1 vccd1 vccd1 seq.encode.inter_keys\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6908_ _3175_ _3172_ _3180_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__nand3_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6839_ sound2.count_m\[18\] _3132_ _3134_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5170_ _0685_ _1562_ _1572_ _1126_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__o221a_1
X_4121_ _0612_ seq.encode.keys_edge_det\[6\] vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__nor2_1
X_4052_ _0676_ _0675_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__nor2_2
Xinput4 piano_keys[0] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_7811_ net107 seq.player_6.next_state\[1\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_6.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_7742_ net137 _0027_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[27\] sky130_fd_sc_hd__dfrtp_1
X_4954_ sound2.count\[0\] _1504_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[0\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3905_ rate_clk.count\[6\] rate_clk.count\[7\] _0552_ vssd1 vssd1 vccd1 vccd1 _0574_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7673_ sound4.sdiv.A\[19\] _2038_ _3728_ vssd1 vssd1 vccd1 vccd1 _3730_ sky130_fd_sc_hd__a21oi_1
X_4885_ _1135_ _1321_ _1333_ _1127_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6624_ _2983_ _2986_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__and2_1
X_3836_ _0471_ _0487_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__nand2_1
X_6555_ _2924_ _2925_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3767_ _0449_ inputcont.INTERNAL_SYNCED_I\[2\] inputcont.INTERNAL_SYNCED_I\[4\] _0450_
+ inputcont.INTERNAL_SYNCED_I\[0\] vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__a221o_1
X_5506_ sound4.count\[16\] sound4.count\[17\] sound4.count\[18\] _1988_ vssd1 vssd1
+ vccd1 vccd1 _1999_ sky130_fd_sc_hd__nand4_1
XFILLER_0_30_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8225_ net129 sound3.osc.next_count\[6\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_6486_ _1170_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5437_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8156_ net132 _0277_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5368_ _0677_ _1038_ _1796_ _1769_ _1059_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__o32a_1
X_5299_ _0954_ _1781_ _1805_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__o211ai_4
X_8087_ net117 _0229_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[22\] sky130_fd_sc_hd__dfrtp_1
X_7107_ sound2.sdiv.A\[23\] _3329_ vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__nand2_1
X_4319_ select1.sequencer_on _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__and2_1
X_7038_ _3164_ _3297_ _3298_ _3174_ sound2.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _0222_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4670_ _0969_ _1101_ _1240_ _0943_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6340_ _2569_ _2753_ sound3.sdiv.Q\[8\] _2301_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _2698_ _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5222_ sound3.count\[10\] _1741_ _1721_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o21ai_1
X_8010_ net128 _0152_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[11\] sky130_fd_sc_hd__dfrtp_1
X_5153_ _1095_ _1559_ _1553_ _1127_ _1591_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__o221a_1
X_4104_ seq.player_7.state\[2\] seq.player_7.state\[3\] vssd1 vssd1 vccd1 vccd1 _0726_
+ sky130_fd_sc_hd__nand2_1
X_5084_ _1610_ _1612_ _1614_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__and3_1
X_4035_ _0675_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _2408_ _2411_ _2412_ _2421_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__nor4_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7725_ net121 _0010_ net82 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[10\] sky130_fd_sc_hd__dfrtp_1
X_4937_ _1001_ _1480_ _1482_ _1487_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__o211a_2
XFILLER_0_74_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4868_ _0695_ _0499_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__or2_1
X_7656_ sound4.sdiv.A\[15\] _2183_ sound4.sdiv.next_dived _3718_ vssd1 vssd1 vccd1
+ vccd1 _0420_ sky130_fd_sc_hd__a22o_1
X_6607_ _2966_ _2964_ _2971_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3819_ _0492_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7587_ sound4.divisor_m\[12\] _1924_ _2186_ vssd1 vssd1 vccd1 vccd1 _3672_ sky130_fd_sc_hd__mux2_1
X_4799_ _1014_ _1338_ _1339_ _0688_ _1349_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__o221a_1
X_6538_ sound1.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6469_ _2861_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
X_8208_ net144 _0329_ net105 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[23\] sky130_fd_sc_hd__dfrtp_1
X_8139_ net109 _0260_ net70 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap66 _0559_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5840_ wave.mode\[0\] net1 wave.mode\[1\] vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__or3b_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ wave_comb.u1.M\[0\] wave_comb.u1.M\[1\] wave_comb.u1.M\[2\] _2209_ vssd1 vssd1
+ vccd1 vccd1 _2223_ sky130_fd_sc_hd__o31a_1
XFILLER_0_29_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7510_ _2275_ _3653_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__nand2_1
X_4722_ _1283_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7441_ sound3.sdiv.A\[19\] _3463_ sound3.sdiv.next_dived _3598_ vssd1 vssd1 vccd1
+ vccd1 _0325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4653_ sound1.count\[18\] _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__xnor2_1
X_7372_ _3534_ _3536_ vssd1 vssd1 vccd1 vccd1 _3537_ sky130_fd_sc_hd__or2_1
X_4584_ _0950_ _1125_ _1154_ _1000_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6323_ net1 wave.mode\[1\] wave.mode\[0\] vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__or3b_2
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6254_ sound2.sdiv.Q\[4\] _2660_ _2661_ vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5205_ sound3.count\[4\] _1728_ _1731_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
X_6185_ _2617_ _2599_ _2618_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5136_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5067_ _1134_ _1578_ _1553_ _1139_ _1597_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__o221a_1
X_4018_ _0662_ _0666_ vssd1 vssd1 vccd1 vccd1 seq.tempo_select.next_state\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5969_ sound1.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__inv_2
X_7708_ _3753_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7639_ _1763_ _3705_ _3706_ sound4.sdiv.next_start _2070_ vssd1 vssd1 vccd1 vccd1
+ _0415_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7990_ net125 sound1.osc.next_count\[11\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_6941_ sound2.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6872_ _1360_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5823_ _0646_ _2264_ _2265_ _0573_ wave_comb.u1.C\[1\] vssd1 vssd1 vccd1 vccd1 _0040_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ wave_comb.u1.next_dived _2207_ _2208_ _0573_ wave_comb.u1.A\[0\] vssd1 vssd1
+ vccd1 vccd1 _0028_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4705_ _1269_ _1270_ _1256_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__and3b_1
XFILLER_0_72_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5685_ sound4.sdiv.A\[18\] _2038_ _2158_ _2166_ _2167_ vssd1 vssd1 vccd1 vccd1 _2168_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7424_ _3569_ _3575_ _3573_ vssd1 vssd1 vccd1 vccd1 _3584_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4636_ _0958_ _1027_ _1203_ _1206_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__o211a_1
X_7355_ _3503_ _3507_ _3521_ _3511_ vssd1 vssd1 vccd1 vccd1 _3522_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6306_ sound4.sdiv.Q\[6\] _0576_ _2736_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__a21o_1
X_4567_ _0685_ _0678_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__nand2_8
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7286_ _3458_ _3459_ vssd1 vssd1 vccd1 vccd1 _3460_ sky130_fd_sc_hd__or2_1
X_4498_ _0949_ _0937_ _0974_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6237_ _2636_ _2669_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__xor2_1
X_6168_ sound3.sdiv.Q\[2\] _0577_ _2602_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__a21oi_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _1010_ _1567_ _1574_ _1027_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__o22a_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ sound3.divisor_m\[11\] sound3.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2535_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5470_ sound4.count\[10\] _1966_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4421_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7140_ sound2.sdiv.C\[5\] _0554_ vssd1 vssd1 vccd1 vccd1 _3384_ sky130_fd_sc_hd__and2_1
X_4352_ seq.player_3.state\[2\] _0881_ _0883_ _0922_ vssd1 vssd1 vccd1 vccd1 _0923_
+ sky130_fd_sc_hd__a22o_1
X_4283_ _0791_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__nor2_1
X_7071_ sound2.sdiv.A\[26\] _3327_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__nor2_1
X_6022_ _2454_ _2455_ _2456_ _2457_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__and4b_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7973_ net131 _0136_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6924_ _2484_ _3195_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6855_ sound2.divisor_m\[6\] _1378_ _3142_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__mux2_1
X_3998_ _0652_ _0653_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[5\] sky130_fd_sc_hd__nor2_1
X_5806_ _2249_ _2252_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6786_ sound1.sdiv.Q\[13\] _2893_ _2890_ sound1.sdiv.Q\[12\] _2842_ vssd1 vssd1 vccd1
+ vccd1 _0154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5737_ sound4.sdiv.Q\[20\] _2182_ _2185_ sound4.sdiv.Q\[19\] _2199_ vssd1 vssd1 vccd1
+ vccd1 _0020_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7407_ _3437_ _3567_ _3568_ _3440_ sound3.sdiv.A\[15\] vssd1 vssd1 vccd1 vccd1 _0321_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5668_ _2145_ _2150_ _2147_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4619_ _0950_ _1004_ _1189_ _0969_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5599_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__inv_2
X_7338_ _3495_ _3499_ _3505_ vssd1 vssd1 vccd1 vccd1 _3507_ sky130_fd_sc_hd__a21o_1
X_7269_ sound3.divisor_m\[0\] sound3.sdiv.Q\[27\] _3443_ vssd1 vssd1 vccd1 vccd1 _3445_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4970_ sound2.count\[3\] sound2.count\[4\] _1508_ sound2.count\[5\] vssd1 vssd1 vccd1
+ vccd1 _1516_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3921_ _0581_ _0583_ _0584_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__and4b_1
X_6640_ sound1.divisor_m\[12\] sound1.divisor_m\[11\] _2984_ vssd1 vssd1 vccd1 vccd1
+ _3002_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3852_ _0478_ _0485_ _0479_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6571_ _2936_ _2939_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8310_ net123 _0410_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5522_ _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[7\] sky130_fd_sc_hd__nor2_1
X_3783_ inputcont.INTERNAL_SYNCED_I\[3\] _0460_ _0462_ _0464_ vssd1 vssd1 vccd1 vccd1
+ net37 sky130_fd_sc_hd__a211o_1
XFILLER_0_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8241_ net143 _0341_ net104 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[2\] sky130_fd_sc_hd__dfrtp_2
X_5453_ _1779_ _1936_ _1956_ _1957_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8172_ net135 _0293_ net96 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[6\] sky130_fd_sc_hd__dfrtp_4
X_4404_ _0918_ _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5384_ _1015_ _1769_ _1784_ _1083_ _1833_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7123_ _3359_ _3367_ _3372_ _3370_ vssd1 vssd1 vccd1 vccd1 _3373_ sky130_fd_sc_hd__a31o_1
X_4335_ seq.player_3.state\[1\] _0881_ _0883_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_
+ sky130_fd_sc_hd__a22o_1
X_7054_ _3312_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__inv_2
X_4266_ seq.clk_div.count\[14\] seq.clk_div.count\[15\] _0841_ vssd1 vssd1 vccd1 vccd1
+ _0847_ sky130_fd_sc_hd__and3_1
X_4197_ seq.clk_div.count\[20\] vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__inv_2
X_6005_ sound2.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7956_ net130 _0119_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7887_ net144 net16 net105 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6907_ _3175_ _3172_ _3180_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__a21o_1
X_6838_ sound2.count\[18\] _2855_ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6769_ sound1.sdiv.C\[5\] _2843_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4120_ _0734_ _0733_ _0736_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_6.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4051_ _0693_ vssd1 vssd1 vccd1 vccd1 oct.next_state\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 piano_keys[10] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_1
X_7810_ net107 seq.player_6.next_state\[0\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_6.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7741_ net137 _0026_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4953_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__buf_4
X_3904_ _0573_ vssd1 vssd1 vccd1 vccd1 wave_comb.u1.next_start sky130_fd_sc_hd__inv_2
XFILLER_0_74_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7672_ sound4.sdiv.A\[20\] _2183_ _3681_ _3729_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__a22o_1
X_6623_ _2983_ _2986_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4884_ _1134_ _1338_ _1322_ _1041_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__o22a_1
X_3835_ _0509_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_4
XFILLER_0_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6554_ _2909_ _2915_ _2913_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__o21ai_1
X_3766_ _0443_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
X_6485_ _2871_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
X_5505_ sound4.count\[16\] sound4.count\[17\] _1988_ sound4.count\[18\] vssd1 vssd1
+ vccd1 vccd1 _1998_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8224_ net129 sound3.osc.next_count\[5\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5436_ sound4.count\[3\] _1940_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8155_ net131 _0276_ net92 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[8\] sky130_fd_sc_hd__dfrtp_1
X_5367_ _0959_ _1133_ _1786_ _1790_ _0983_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__o32a_1
XFILLER_0_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5298_ _0996_ _1784_ _1806_ _1808_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__o211a_1
X_8086_ net119 _0228_ net80 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[21\] sky130_fd_sc_hd__dfrtp_1
X_7106_ sound2.sdiv.A\[23\] _3329_ vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__or2_1
X_4318_ seq.beat\[3\] seq.encode.play _0870_ inputcont.INTERNAL_SYNCED_I\[4\] vssd1
+ vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__a31o_1
X_7037_ _3286_ _3290_ _3296_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__a21o_1
X_4249_ _0834_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ net125 _0102_ net86 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[13\] sky130_fd_sc_hd__dfrtp_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6270_ _2289_ _2700_ _2701_ _2301_ sound3.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 _2702_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5221_ _1741_ _1742_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[9\] sky130_fd_sc_hd__nor2_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5152_ sound3.count\[12\] _1681_ _1655_ sound3.count\[2\] _1682_ vssd1 vssd1 vccd1
+ vccd1 _1683_ sky130_fd_sc_hd__o221a_1
X_4103_ seq.player_7.state\[2\] seq.player_7.state\[3\] _0724_ _0725_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_7.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_5083_ _1011_ _1559_ _1613_ _1590_ _1591_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4034_ _0676_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__nand2_8
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5985_ sound1.count_m\[2\] _2413_ _2414_ _2418_ _2420_ vssd1 vssd1 vccd1 vccd1 _2421_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7724_ net120 _0009_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[9\] sky130_fd_sc_hd__dfrtp_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4936_ _1004_ _1483_ _1484_ _1486_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__o211a_1
XANTENNA_10 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4867_ _1314_ _1315_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7655_ _3717_ _2148_ vssd1 vssd1 vccd1 vccd1 _3718_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6606_ _2966_ _2964_ _2971_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7586_ _3671_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3818_ _0474_ _0491_ _0494_ _0495_ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__a221o_1
X_6537_ _2901_ _2906_ _2908_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4798_ _1199_ _1341_ _1343_ _1200_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6468_ sound1.divisor_m\[1\] _1008_ _2005_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__mux2_1
X_8207_ net142 _0328_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[22\] sky130_fd_sc_hd__dfrtp_1
X_6399_ _2819_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5419_ _0973_ _1786_ _1928_ _1929_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__o211a_1
X_8138_ net109 _0259_ net70 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[19\] sky130_fd_sc_hd__dfrtp_1
X_8069_ net117 _0211_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap67 _0483_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap56 _0542_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_2
XFILLER_0_78_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5770_ _2216_ _2218_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _1281_ _1282_ _1256_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7440_ _3596_ _3597_ vssd1 vssd1 vccd1 vccd1 _3598_ sky130_fd_sc_hd__xnor2_1
X_4652_ _1222_ _1216_ _1070_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7371_ sound3.divisor_m\[12\] _3535_ vssd1 vssd1 vccd1 vccd1 _3536_ sky130_fd_sc_hd__xnor2_1
X_4583_ _1018_ _0978_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__or2_4
XFILLER_0_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6322_ _2407_ _2432_ _2412_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6253_ sound2.sdiv.Q\[6\] _2295_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5204_ sound3.count\[4\] _1728_ _1721_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__o21ai_1
X_6184_ _2590_ _2595_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__nand2_1
X_5135_ _1591_ _1660_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5066_ _1129_ _1572_ _1574_ _1141_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4017_ _0664_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__nand2_1
X_5968_ _2397_ _2400_ _2401_ _2403_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7707_ sound4.sdiv.C\[5\] _0554_ vssd1 vssd1 vccd1 vccd1 _3753_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4919_ sound2.count\[2\] vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5899_ _2333_ sound4.divisor_m\[10\] sound4.divisor_m\[9\] _2334_ vssd1 vssd1 vccd1
+ vccd1 _2335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7638_ _2079_ _2137_ vssd1 vssd1 vccd1 vccd1 _3706_ sky130_fd_sc_hd__and2_1
X_7569_ _3661_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6940_ _3164_ _3209_ _3210_ _3174_ sound2.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _0212_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6871_ _3154_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5822_ wave_comb.u1.C\[0\] wave_comb.u1.C\[1\] vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5753_ wave_comb.u1.M\[0\] wave_comb.u1.Q\[11\] vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4704_ sound1.count\[4\] _1263_ sound1.count\[5\] vssd1 vssd1 vccd1 vccd1 _1270_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5684_ sound4.sdiv.A\[18\] _2038_ _2162_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7423_ _3581_ _3582_ vssd1 vssd1 vccd1 vccd1 _3583_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4635_ _0688_ _0967_ _0969_ _1204_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7354_ _3510_ vssd1 vssd1 vccd1 vccd1 _3521_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4566_ _0696_ _0939_ _1003_ _1041_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6305_ sound4.sdiv.Q\[5\] _2641_ _2704_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7285_ _3455_ _3457_ vssd1 vssd1 vccd1 vccd1 _3459_ sky130_fd_sc_hd__and2_1
X_4497_ _0677_ _0976_ _1038_ _1054_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__o311a_1
X_6236_ sound3.sdiv.Q\[3\] _2632_ _2633_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__a21o_1
X_6167_ _2570_ _2601_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__nor2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _1643_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ sound3.divisor_m\[10\] sound3.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2534_
+ sky130_fd_sc_hd__and2b_1
X_5049_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4420_ _0988_ _0937_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4351_ seq.player_4.state\[2\] _0886_ _0888_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4282_ seq.clk_div.count\[19\] _0855_ _0858_ _0813_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[19\]
+ sky130_fd_sc_hd__o211a_1
X_7070_ _3308_ _2471_ _2470_ vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__and3b_1
X_6021_ sound2.divisor_m\[9\] sound2.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__or2b_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7972_ net131 _0135_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.C\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6923_ _3177_ _3194_ vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__nand2_1
X_6854_ _3143_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
X_3997_ pm.count\[4\] _0649_ pm.count\[5\] vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__a21oi_1
X_5805_ _2250_ _2251_ _2240_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__or3b_1
XFILLER_0_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6785_ sound1.sdiv.Q\[12\] _2893_ _2890_ sound1.sdiv.Q\[11\] _2841_ vssd1 vssd1 vccd1
+ vccd1 _0153_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5736_ sound4.count\[12\] _2186_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5667_ _2149_ _2056_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7406_ _3555_ _3559_ _3566_ vssd1 vssd1 vccd1 vccd1 _3568_ sky130_fd_sc_hd__a21o_1
X_4618_ _1001_ net63 vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nor2_4
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5598_ sound4.divisor_m\[9\] _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__xnor2_1
X_7337_ _3495_ _3499_ _3505_ vssd1 vssd1 vccd1 vccd1 _3506_ sky130_fd_sc_hd__nand3_1
X_4549_ _1107_ _1108_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7268_ _3438_ _3443_ vssd1 vssd1 vccd1 vccd1 _3444_ sky130_fd_sc_hd__or2b_1
X_6219_ _2650_ _2652_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__xnor2_1
X_7199_ sound3.count_m\[13\] _3132_ _3400_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _0529_ _0549_ _0582_ _0525_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3851_ _0478_ _0485_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__or2_2
XFILLER_0_128_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6570_ sound1.divisor_m\[6\] _2938_ vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__xnor2_1
X_3782_ inputcont.INTERNAL_SYNCED_I\[6\] _0463_ _0450_ vssd1 vssd1 vccd1 vccd1 _0464_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5521_ rate_clk.count\[7\] _0553_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8240_ net143 _0340_ net104 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5452_ sound4.count\[6\] _1951_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__or2_1
X_8171_ net135 _0292_ net96 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[5\] sky130_fd_sc_hd__dfrtp_2
X_4403_ _0909_ _0936_ _0926_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__or3b_4
X_5383_ _1079_ _1800_ _1794_ _0952_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7122_ _3360_ _3363_ _3366_ vssd1 vssd1 vccd1 vccd1 _3372_ sky130_fd_sc_hd__or3_1
X_4334_ seq.player_4.state\[1\] _0886_ _0888_ _0904_ vssd1 vssd1 vccd1 vccd1 _0905_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7053_ sound2.sdiv.A\[16\] _3311_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__nand2_1
X_6004_ sound2.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__inv_2
X_4265_ _0846_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4196_ _0789_ seq.clk_div.count\[14\] seq.tempo_select.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0790_ sky130_fd_sc_hd__a21oi_1
X_7955_ net130 _0118_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7886_ net110 net15 net71 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6906_ _3176_ _3179_ vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6837_ sound2.count_m\[17\] _3132_ _3133_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6768_ _3111_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6699_ _3054_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5719_ sound4.sdiv.Q\[11\] _2182_ _2185_ sound4.sdiv.Q\[10\] _2190_ vssd1 vssd1 vccd1
+ vccd1 _0011_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8369_ net119 rate_clk.next_count\[6\] net80 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4050_ _0679_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__or2_1
Xinput6 piano_keys[11] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7740_ net137 _0025_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[25\] sky130_fd_sc_hd__dfrtp_1
X_4952_ _1317_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3903_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7671_ _3727_ _3728_ vssd1 vssd1 vccd1 vccd1 _3729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4883_ _1317_ _1426_ _1431_ _1433_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__and4_2
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6622_ sound1.divisor_m\[11\] _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__xnor2_1
X_3834_ net1 wave.mode\[1\] vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6553_ _2922_ _2923_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3765_ inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
X_6484_ sound1.divisor_m\[7\] _1089_ _2864_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__mux2_1
X_5504_ _1997_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_8223_ net129 sound3.osc.next_count\[4\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_5435_ _1943_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8154_ net132 _0275_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[7\] sky130_fd_sc_hd__dfrtp_1
X_5366_ sound4.count\[13\] _1875_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__or2_1
X_5297_ _1182_ _1794_ _1796_ _1175_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__o221a_1
X_8085_ net118 _0227_ net79 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[20\] sky130_fd_sc_hd__dfrtp_1
X_7105_ sound2.sdiv.A\[23\] _3168_ sound2.sdiv.next_dived _3357_ vssd1 vssd1 vccd1
+ vccd1 _0230_ sky130_fd_sc_hd__a22o_1
X_4317_ _0886_ _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__nand2_1
X_7036_ _3286_ _3290_ _3296_ vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__nand3_1
X_4248_ _0832_ _0813_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4179_ seq.player_1.state\[1\] seq.player_1.state\[2\] _0770_ seq.player_1.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__a31o_1
X_7938_ net127 _0101_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[12\] sky130_fd_sc_hd__dfrtp_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7869_ net113 inputcont.u1.ff_intermediate\[0\] net74 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5220_ sound3.count\[9\] _1738_ _1721_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5151_ sound3.count\[1\] _1673_ _1666_ sound3.count\[13\] vssd1 vssd1 vccd1 vccd1
+ _1682_ sky130_fd_sc_hd__o2bb2a_1
X_5082_ _1138_ _1551_ _1568_ _0688_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__o22a_1
X_4102_ seq.player_7.state\[1\] _0722_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4033_ oct.state\[0\] vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__buf_12
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ sound1.count_m\[3\] _2419_ sound1.divisor_m\[1\] _2415_ vssd1 vssd1 vccd1
+ vccd1 _2420_ sky130_fd_sc_hd__a22o_1
X_7723_ net136 _0008_ net97 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4935_ _0947_ _1325_ _1485_ _1033_ _1341_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__o32a_1
XANTENNA_11 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7654_ _2150_ _3715_ vssd1 vssd1 vccd1 vccd1 _3717_ sky130_fd_sc_hd__nand2_1
X_4866_ _0680_ _1321_ _1415_ _1416_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__o211a_1
X_6605_ _2969_ _2970_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7585_ sound4.divisor_m\[11\] _3670_ _2186_ vssd1 vssd1 vccd1 vccd1 _3671_ sky130_fd_sc_hd__mux2_1
X_3817_ inputcont.INTERNAL_SYNCED_I\[2\] _0459_ _0481_ vssd1 vssd1 vccd1 vccd1 _0496_
+ sky130_fd_sc_hd__and3_1
X_4797_ _0683_ _1107_ _1345_ _1347_ _1146_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__o32a_1
X_6536_ _2902_ _2905_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6467_ _2860_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
X_8206_ net144 _0327_ net105 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6398_ _2659_ _2682_ _2805_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5418_ _0959_ _0993_ _1800_ _1792_ _0869_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__o32a_1
X_5349_ sound4.count\[0\] _1859_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8137_ net109 _0258_ net70 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8068_ net117 _0210_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[3\] sky130_fd_sc_hd__dfrtp_1
X_7019_ _3164_ _3280_ _3281_ _3174_ sound2.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _0220_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ sound1.count\[9\] _1278_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4651_ _0685_ _0684_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 seq_power vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7370_ sound3.divisor_m\[11\] _3526_ _3448_ vssd1 vssd1 vccd1 vccd1 _3535_ sky130_fd_sc_hd__o21a_1
X_4582_ _0939_ _1134_ _1151_ _0981_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6321_ _2749_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6252_ _2678_ _2679_ _2683_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6183_ _2590_ _2595_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__nor2_1
X_5203_ _1730_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5134_ _0952_ _1025_ _1559_ _1661_ _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _1138_ _1562_ _1567_ _0696_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4016_ seq.tempo_select.state\[1\] seq.tempo_select.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _0665_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5967_ sound1.divisor_m\[5\] _2399_ _2402_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7706_ _3752_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__clkbuf_1
X_4918_ _1466_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5898_ sound4.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__inv_2
X_7637_ _2079_ _2137_ vssd1 vssd1 vccd1 vccd1 _3705_ sky130_fd_sc_hd__nor2_1
X_4849_ _0985_ _1323_ _1338_ _0948_ _1399_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__o221a_1
X_7568_ sound4.divisor_m\[4\] _1866_ _3419_ vssd1 vssd1 vccd1 vccd1 _3661_ sky130_fd_sc_hd__mux2_1
X_7499_ _3643_ _3644_ _3646_ _3440_ sound3.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 _0335_
+ sky130_fd_sc_hd__a32o_1
X_6519_ _2893_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6870_ sound2.divisor_m\[11\] _3153_ _3142_ vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__mux2_1
X_5821_ wave_comb.u1.C\[0\] wave_comb.u1.C\[1\] vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5752_ wave_comb.u1.M\[0\] wave_comb.u1.Q\[11\] vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4703_ sound1.count\[4\] sound1.count\[5\] _1263_ vssd1 vssd1 vccd1 vccd1 _1269_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5683_ _2164_ _2165_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__nor2_1
X_7422_ _3577_ _3580_ vssd1 vssd1 vccd1 vccd1 _3582_ sky130_fd_sc_hd__nand2_1
X_4634_ _0683_ _1107_ _1000_ _0943_ _1014_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7353_ _3518_ _3519_ vssd1 vssd1 vccd1 vccd1 _3520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4565_ _0943_ _1134_ _1135_ _0950_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6304_ _2730_ _2734_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__xor2_1
X_7284_ _3455_ _3457_ vssd1 vssd1 vccd1 vccd1 _3458_ sky130_fd_sc_hd__nor2_1
X_4496_ _0990_ _1056_ _1061_ _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__o211a_1
X_6235_ _2666_ _2667_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6166_ sound3.sdiv.Q\[0\] sound3.sdiv.Q\[1\] _0577_ vssd1 vssd1 vccd1 vccd1 _2601_
+ sky130_fd_sc_hd__o21ai_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _2531_ sound3.divisor_m\[10\] sound3.divisor_m\[9\] _2532_ vssd1 vssd1 vccd1
+ vccd1 _2533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5117_ _0971_ _1578_ _1645_ _1647_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__o211a_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5048_ _1551_ _1563_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6999_ _3262_ _3263_ vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4350_ seq.player_5.state\[2\] _0890_ _0892_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4281_ seq.clk_div.count\[18\] seq.clk_div.count\[19\] _0853_ vssd1 vssd1 vccd1 vccd1
+ _0858_ sky130_fd_sc_hd__nand3_1
X_6020_ sound2.count_m\[9\] sound2.divisor_m\[10\] vssd1 vssd1 vccd1 vccd1 _2456_
+ sky130_fd_sc_hd__or2b_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7971_ net130 _0134_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6922_ sound2.divisor_m\[3\] sound2.divisor_m\[2\] sound2.divisor_m\[1\] sound2.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__or4_1
X_6853_ sound2.divisor_m\[5\] _3141_ _3142_ vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__mux2_1
X_5804_ wave_comb.u1.A\[6\] wave_comb.u1.A\[5\] _2224_ vssd1 vssd1 vccd1 vccd1 _2251_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3996_ pm.count\[5\] pm.count\[4\] _0649_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__and3_1
X_6784_ sound1.sdiv.Q\[11\] _2893_ _2890_ sound1.sdiv.Q\[10\] _2840_ vssd1 vssd1 vccd1
+ vccd1 _0152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5735_ sound4.sdiv.Q\[19\] _2182_ _2185_ sound4.sdiv.Q\[18\] _2198_ vssd1 vssd1 vccd1
+ vccd1 _0019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5666_ sound4.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__inv_2
X_7405_ _3555_ _3559_ _3566_ vssd1 vssd1 vccd1 vccd1 _3567_ sky130_fd_sc_hd__nand3_1
XFILLER_0_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4617_ _0676_ _1003_ _1083_ _1000_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5597_ _2036_ _2029_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7336_ _3503_ _3504_ vssd1 vssd1 vccd1 vccd1 _3505_ sky130_fd_sc_hd__nand2_1
X_4548_ _0676_ _1003_ _1034_ _1109_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o311a_1
XFILLER_0_111_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7267_ sound3.sdiv.A\[0\] _3442_ vssd1 vssd1 vccd1 vccd1 _3443_ sky130_fd_sc_hd__xnor2_1
X_4479_ _1037_ _1045_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__and3_2
XFILLER_0_110_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6218_ _2610_ _2612_ _2651_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__a21bo_1
X_7198_ _1658_ _2843_ vssd1 vssd1 vccd1 vccd1 _3400_ sky130_fd_sc_hd__nor2_1
X_6149_ sound4.sdiv.Q\[2\] _0576_ _2582_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__a21o_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3850_ _0473_ _0486_ _0521_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__nor4_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ inputcont.INTERNAL_SYNCED_I\[5\] inputcont.INTERNAL_SYNCED_I\[4\] vssd1 vssd1
+ vccd1 vccd1 _0463_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5520_ _0575_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5451_ _1955_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__inv_2
X_8170_ net135 _0291_ net96 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[4\] sky130_fd_sc_hd__dfrtp_4
X_4402_ _0971_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__or2_4
X_5382_ _0684_ _1077_ _1792_ _1781_ _1039_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__o32a_1
XFILLER_0_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7121_ _3365_ _3366_ _3367_ _3370_ vssd1 vssd1 vccd1 vccd1 _3371_ sky130_fd_sc_hd__o211ai_1
X_4333_ seq.player_5.state\[1\] _0890_ _0892_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_
+ sky130_fd_sc_hd__a22o_1
X_7052_ _3310_ vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__inv_2
X_4264_ _0844_ _0813_ _0845_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__and3b_1
X_6003_ _2289_ _2437_ _2438_ _2293_ sound1.sdiv.Q\[2\] vssd1 vssd1 vccd1 vccd1 _2439_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ seq.clk_div.count\[2\] vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__inv_2
X_7954_ net130 _0117_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6905_ sound2.divisor_m\[2\] _3178_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__xnor2_1
X_7885_ net108 net14 net69 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6836_ sound2.count\[17\] _2855_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6767_ _2843_ _3110_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__and2_1
X_5718_ sound4.count\[3\] _2186_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3979_ _0640_ _0641_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6698_ sound1.divisor_m\[18\] sound1.divisor_m\[17\] _3036_ _2903_ vssd1 vssd1 vccd1
+ vccd1 _3054_ sky130_fd_sc_hd__o31a_1
XFILLER_0_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5649_ _2099_ _2131_ _2097_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8368_ net119 rate_clk.next_count\[5\] net80 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7319_ _3477_ _3480_ _3488_ vssd1 vssd1 vccd1 vccd1 _3490_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8299_ net122 _0399_ net83 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 piano_keys[12] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4951_ _1370_ _1414_ _1443_ _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__or4_1
X_3902_ _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7670_ _2041_ _2168_ vssd1 vssd1 vccd1 vccd1 _3728_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4882_ _0952_ _1025_ _1339_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__o31a_1
XFILLER_0_129_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6621_ _2903_ _2984_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__and2_1
X_3833_ _0508_ _0477_ _0505_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__a21o_2
XFILLER_0_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6552_ _2918_ _2921_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3764_ _0443_ _0444_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6483_ _2870_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5503_ _1779_ _1936_ _1995_ _1996_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__and4_1
XFILLER_0_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8222_ net128 sound3.osc.next_count\[3\] net89 vssd1 vssd1 vccd1 vccd1 sound3.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5434_ _1779_ _1936_ _1941_ _1942_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8153_ net132 _0274_ net93 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7104_ _3355_ _3356_ vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__xnor2_1
X_5365_ sound4.count\[13\] _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__nand2_1
X_5296_ _1129_ _1800_ _1792_ _1026_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__o22a_1
X_8084_ net118 _0226_ net79 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[19\] sky130_fd_sc_hd__dfrtp_1
X_4316_ seq.player_4.state\[0\] seq.player_4.state\[1\] seq.player_4.state\[2\] seq.player_4.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__or4_1
X_7035_ _3294_ _3295_ vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__nand2_1
X_4247_ seq.clk_div.count\[10\] _0829_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__or2_1
X_4178_ _0774_ _0773_ _0775_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_1.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7937_ net126 _0100_ net87 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[11\] sky130_fd_sc_hd__dfrtp_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7868_ net113 seq.encode.inter_keys\[1\] net74 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_sync\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6819_ sound2.count\[9\] _2855_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7799_ net113 oct.next_state\[0\] net74 vssd1 vssd1 vccd1 vccd1 oct.state\[0\] sky130_fd_sc_hd__dfstp_4
XFILLER_0_18_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5150_ _1675_ _1677_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__and3_2
X_5081_ _1611_ _1565_ _1213_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__a21o_1
X_4101_ seq.player_7.state\[0\] seq.player_7.state\[1\] _0721_ vssd1 vssd1 vccd1 vccd1
+ _0724_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4032_ oct.state\[1\] vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__buf_12
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5983_ sound1.divisor_m\[4\] vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7722_ net137 _0007_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[7\] sky130_fd_sc_hd__dfrtp_1
X_4934_ _0977_ _1419_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_12 net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7653_ _3681_ _3715_ _3716_ _2184_ sound4.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _0419_
+ sky130_fd_sc_hd__a32o_1
X_4865_ _1347_ _1323_ _0687_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6604_ sound1.sdiv.A\[8\] _2968_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4796_ _1346_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__buf_4
X_3816_ _0480_ _0481_ _0482_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__and3_1
X_7584_ _1909_ vssd1 vssd1 vccd1 vccd1 _3670_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6535_ sound1.sdiv.A\[2\] _2895_ sound1.sdiv.next_dived _2907_ vssd1 vssd1 vccd1
+ vccd1 _0110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8205_ net142 _0326_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[20\] sky130_fd_sc_hd__dfrtp_2
X_6466_ sound1.divisor_m\[0\] _2859_ _2005_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6397_ _2818_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5417_ _0985_ _1769_ _1796_ _0979_ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8136_ net110 _0257_ net71 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[17\] sky130_fd_sc_hd__dfrtp_1
X_5348_ _1041_ _1769_ _1777_ _1101_ _1858_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__o221ai_4
X_8067_ net117 _0209_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[2\] sky130_fd_sc_hd__dfrtp_1
X_7018_ _3268_ _3272_ _3279_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__nand3_1
X_5279_ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap58 net35 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_4
XFILLER_0_93_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4650_ sound1.count\[15\] _1215_ _1219_ sound1.count\[16\] vssd1 vssd1 vccd1 vccd1
+ _1221_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput21 tempo_select vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 piano_keys[1] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_6320_ sound1.sdiv.Q\[7\] _0579_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__nand2_1
X_4581_ _1107_ _1003_ _1040_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6251_ _2676_ _2677_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__or2b_1
XFILLER_0_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6182_ wave_comb.u1.next_start _2615_ _2616_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__a21o_1
X_5202_ _1728_ _1729_ _1721_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5133_ _1016_ _1553_ _1567_ _0997_ _1663_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ sound3.count\[6\] _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4015_ seq.tempo_select.state\[1\] seq.tempo_select.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _0664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5966_ sound1.divisor_m\[8\] sound1.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7705_ _2843_ _3751_ vssd1 vssd1 vccd1 vccd1 _3752_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4917_ _1014_ _1322_ _1467_ _0499_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__o22a_1
X_5897_ sound4.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4848_ _0954_ _1321_ _1327_ _0973_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__o22a_1
X_7636_ _3681_ _3703_ _3704_ _2184_ sound4.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 _0414_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7567_ _3660_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__clkbuf_1
X_4779_ _0698_ _0499_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7498_ _3645_ vssd1 vssd1 vccd1 vccd1 _3646_ sky130_fd_sc_hd__inv_2
X_6518_ _0579_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6449_ sound1.count\[12\] _2201_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8119_ net136 _0240_ net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _2263_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__clkbuf_1
X_5751_ sound4.sdiv.Q\[27\] _2183_ sound4.sdiv.next_dived sound4.sdiv.Q\[26\] vssd1
+ vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4702_ _1268_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7421_ _3577_ _3580_ vssd1 vssd1 vccd1 vccd1 _3581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5682_ sound4.sdiv.A\[18\] _2037_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _0978_ _0996_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__or2_2
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7352_ _3514_ _3517_ vssd1 vssd1 vccd1 vccd1 _3519_ sky130_fd_sc_hd__nand2_1
X_4564_ _1107_ net63 vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7283_ sound3.divisor_m\[3\] _3456_ vssd1 vssd1 vccd1 vccd1 _3457_ sky130_fd_sc_hd__xnor2_1
X_6303_ sound3.sdiv.Q\[7\] _2301_ _2732_ _2733_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6234_ _2619_ _2629_ _2628_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__a21o_1
X_4495_ _1000_ _1063_ _1064_ _0994_ _1065_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6165_ _2596_ _2599_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ sound3.count_m\[8\] vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__inv_2
X_5116_ _1083_ _1550_ _1565_ _0960_ _1646_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__o221a_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _0540_ _1552_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nand2_8
XFILLER_0_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6998_ _3248_ _3254_ _3261_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__and3_1
X_5949_ sound1.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7619_ _2130_ _2103_ vssd1 vssd1 vccd1 vccd1 _3692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4280_ _0857_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7970_ net131 _0133_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6921_ sound2.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__inv_2
X_6852_ _2863_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__buf_8
XFILLER_0_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5803_ _2239_ _2241_ _2244_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__nor3_1
XFILLER_0_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3995_ _0651_ _0649_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[4\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6783_ sound1.sdiv.Q\[10\] _2894_ _2890_ sound1.sdiv.Q\[9\] _2839_ vssd1 vssd1 vccd1
+ vccd1 _0151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5734_ sound4.count\[11\] _2186_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5665_ _2146_ _2147_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7404_ _3564_ _3565_ vssd1 vssd1 vccd1 vccd1 _3566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4616_ sound1.count\[5\] _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7335_ _3500_ _3502_ vssd1 vssd1 vccd1 vccd1 _3504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5596_ _2077_ _2078_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__nand2_1
X_4547_ _0958_ _1110_ _1115_ _1117_ _1070_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_20_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7266_ sound3.divisor_m\[1\] _3441_ vssd1 vssd1 vccd1 vccd1 _3442_ sky130_fd_sc_hd__xnor2_1
X_4478_ _1001_ _1047_ _1048_ _0947_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__o22a_1
X_7197_ sound3.count_m\[12\] _3132_ _3399_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21o_1
X_6217_ _2607_ _2609_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6148_ sound4.sdiv.Q\[2\] _2582_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__nand2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _2513_ sound3.divisor_m\[7\] _2514_ sound3.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2515_ sky130_fd_sc_hd__o22a_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3780_ _0447_ _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5450_ sound4.count\[6\] _1951_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4401_ _0675_ _0687_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5381_ _0946_ _1786_ _1790_ _0971_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7120_ sound2.sdiv.A\[25\] _3329_ vssd1 vssd1 vccd1 vccd1 _3370_ sky130_fd_sc_hd__xnor2_1
X_4332_ seq.player_6.state\[1\] _0894_ _0896_ _0902_ vssd1 vssd1 vccd1 vccd1 _0903_
+ sky130_fd_sc_hd__a22o_1
X_7051_ sound2.divisor_m\[17\] _3309_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__xnor2_1
X_4263_ seq.clk_div.count\[14\] _0841_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__or2_1
X_6002_ _2435_ _2277_ _2434_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4194_ seq.clk_div.count\[6\] seq.clk_div.count\[12\] seq.clk_div.count\[16\] _0779_
+ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__or4_1
X_7953_ net130 _0116_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6904_ sound2.divisor_m\[1\] sound2.divisor_m\[0\] _3177_ vssd1 vssd1 vccd1 vccd1
+ _3178_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7884_ net109 net13 net70 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6835_ _0554_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__buf_6
X_6766_ sound1.sdiv.C\[3\] _0565_ _3106_ sound1.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1
+ _3110_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3978_ _0446_ _0628_ _0626_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o21a_1
X_5717_ sound4.sdiv.Q\[10\] _2182_ _2185_ sound4.sdiv.Q\[9\] _2189_ vssd1 vssd1 vccd1
+ vccd1 _0010_ sky130_fd_sc_hd__a221o_1
X_6697_ _2890_ _3052_ _3053_ _2894_ sound1.sdiv.A\[18\] vssd1 vssd1 vccd1 vccd1 _0126_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5648_ _2103_ _2129_ _2130_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8367_ net119 rate_clk.next_count\[4\] net80 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5579_ _2060_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7318_ _3477_ _3480_ _3488_ vssd1 vssd1 vccd1 vccd1 _3489_ sky130_fd_sc_hd__nand3_1
X_8298_ net118 _0398_ net79 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[12\] sky130_fd_sc_hd__dfrtp_2
X_7249_ _3430_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput8 piano_keys[13] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _1444_ _1461_ _1479_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__or4_1
X_3901_ wave_comb.u1.C\[3\] wave_comb.u1.C\[2\] _0570_ wave_comb.u1.C\[5\] wave_comb.u1.C\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4881_ _0687_ _1001_ _1338_ _1336_ _1112_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__o32a_1
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6620_ sound1.divisor_m\[10\] _2977_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3832_ _0479_ _0478_ _0485_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__and3_1
X_6551_ _2918_ _2921_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5502_ sound4.count\[15\] sound4.count\[16\] _1984_ sound4.count\[17\] vssd1 vssd1
+ vccd1 vccd1 _1996_ sky130_fd_sc_hd__a31o_1
X_3763_ _0446_ inputcont.INTERNAL_SYNCED_I\[11\] inputcont.INTERNAL_SYNCED_I\[10\]
+ _0445_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or4_2
X_6482_ sound1.divisor_m\[6\] _1071_ _2864_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8221_ net128 sound3.osc.next_count\[2\] net89 vssd1 vssd1 vccd1 vccd1 sound3.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_5433_ sound4.count\[0\] sound4.count\[1\] sound4.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1942_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8152_ net131 _0273_ net92 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[5\] sky130_fd_sc_hd__dfrtp_1
X_5364_ _1778_ _1874_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__nand2_2
X_7103_ sound2.sdiv.A\[21\] _3329_ _3354_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__a21boi_1
X_4315_ select1.sequencer_on _0885_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__and2_1
X_5295_ _1176_ _1769_ _1777_ _1174_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o22a_1
X_8083_ net119 _0225_ net80 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[18\] sky130_fd_sc_hd__dfrtp_1
X_7034_ _3291_ _3293_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__nand2_1
X_4246_ seq.clk_div.count\[8\] seq.clk_div.count\[9\] seq.clk_div.count\[10\] _0824_
+ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__and4_1
X_4177_ seq.player_1.state\[2\] _0772_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7936_ net127 _0099_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7867_ net114 seq.encode.inter_keys\[0\] net75 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_sync\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6818_ sound2.count_m\[8\] _2857_ _3123_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__a21o_1
X_7798_ net142 net9 net103 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6749_ _3096_ _3097_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5080_ net56 _1551_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__or2_1
X_4100_ seq.player_7.state\[0\] _0721_ _0723_ vssd1 vssd1 vccd1 vccd1 seq.player_7.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_4031_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__inv_4
XFILLER_0_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5982_ sound1.divisor_m\[1\] _2415_ _2416_ _2417_ vssd1 vssd1 vccd1 vccd1 _2418_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7721_ net136 _0006_ net97 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4933_ _1041_ _1343_ _1333_ _1129_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__o22a_1
X_7652_ _2061_ _2141_ _2057_ vssd1 vssd1 vccd1 vccd1 _3716_ sky130_fd_sc_hd__a21o_1
X_4864_ _0684_ _1343_ _1333_ _0686_ _1341_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6603_ sound1.sdiv.A\[8\] _2968_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4795_ net39 _1315_ _1319_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__or3_1
X_3815_ _0483_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__nand2_1
X_7583_ _3669_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6534_ _2901_ _2906_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__xor2_1
X_6465_ _1104_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8204_ net142 _0325_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5416_ _0978_ _0944_ _1777_ _1794_ _1001_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__o32a_1
X_6396_ pm.current_waveform\[4\] _2817_ _2808_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8135_ net110 _0256_ net71 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[16\] sky130_fd_sc_hd__dfrtp_1
X_5347_ _0948_ _1800_ _1853_ _1857_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8066_ net117 _0208_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[1\] sky130_fd_sc_hd__dfrtp_1
X_5278_ net47 _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__or2_1
X_4229_ seq.clk_div.count\[4\] _0815_ seq.clk_div.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0820_ sky130_fd_sc_hd__a21o_1
X_7017_ _3268_ _3272_ _3279_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__a21o_1
Xmax_cap59 net60 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7919_ net126 _0082_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4580_ _0696_ _1055_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nand2_2
Xinput11 piano_keys[2] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6250_ wave_comb.u1.next_start _2681_ _2682_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6181_ wave_comb.u1.Q\[3\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__and3_1
X_5201_ sound3.count\[0\] sound3.count\[1\] sound3.count\[2\] sound3.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__a31o_1
X_5132_ _1113_ _1570_ _1574_ _1112_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__o221a_1
X_5063_ _1586_ _1593_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__nand2_1
X_4014_ _0662_ _0663_ vssd1 vssd1 vccd1 vccd1 seq.tempo_select.next_state\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _2396_ sound1.divisor_m\[7\] _2398_ sound1.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2401_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7704_ sound4.sdiv.C\[3\] _0556_ _3747_ sound4.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1
+ _3751_ sky130_fd_sc_hd__a31o_1
X_4916_ _1025_ _1028_ _1325_ _1418_ _1011_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__o32a_1
X_5896_ sound4.count_m\[14\] _2331_ sound4.count_m\[13\] _2142_ vssd1 vssd1 vccd1
+ vccd1 _2332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4847_ _0959_ _0993_ _1341_ _1336_ _0979_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__o32a_1
X_7635_ _2135_ _3702_ vssd1 vssd1 vccd1 vccd1 _3704_ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7566_ sound4.divisor_m\[3\] _1850_ _3419_ vssd1 vssd1 vccd1 vccd1 _3660_ sky130_fd_sc_hd__mux2_1
X_4778_ _0686_ _1321_ _1322_ _1134_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__o221a_1
X_7497_ sound3.sdiv.C\[2\] sound3.sdiv.C\[1\] sound3.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3645_ sky130_fd_sc_hd__and3_1
X_6517_ sound1.divisor_m\[0\] sound1.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6448_ sound1.count_m\[11\] _2836_ _2849_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6379_ net34 _2804_ _0700_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__o21a_4
X_8118_ net140 sound3.sdiv.next_dived net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.dived
+ sky130_fd_sc_hd__dfrtp_1
X_8049_ net112 _0191_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5750_ sound4.sdiv.Q\[26\] _2182_ _2185_ sound4.sdiv.Q\[25\] _2206_ vssd1 vssd1 vccd1
+ vccd1 _0026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4701_ _1256_ _1266_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__and3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5681_ _2162_ _2163_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__or2b_1
X_7420_ sound3.divisor_m\[17\] _3579_ vssd1 vssd1 vccd1 vccd1 _3580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4632_ _1003_ _1134_ _1125_ _0976_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7351_ _3514_ _3517_ vssd1 vssd1 vccd1 vccd1 _3518_ sky130_fd_sc_hd__or2_1
X_4563_ _1107_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__nor2_4
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7282_ sound3.divisor_m\[2\] sound3.divisor_m\[1\] sound3.divisor_m\[0\] _3448_ vssd1
+ vssd1 vccd1 vccd1 _3456_ sky130_fd_sc_hd__o31a_1
X_6302_ sound3.sdiv.Q\[6\] _2731_ _2292_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4494_ _0979_ _1003_ _0943_ _0983_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6233_ _2664_ _2665_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6164_ _2597_ _2506_ _2598_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__a21oi_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ sound3.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5115_ _1078_ _1559_ _1572_ _1039_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__o22a_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5046_ _1041_ _1562_ _1565_ _1101_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6997_ _3248_ _3254_ _3261_ vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5948_ sound1.count_m\[13\] _2376_ _2383_ sound1.count_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2384_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ sound4.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7618_ _3681_ _3690_ _3691_ _2184_ sound4.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 _0409_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7549_ sound4.count_m\[10\] _3403_ _2197_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6920_ sound2.sdiv.A\[3\] _3168_ sound2.sdiv.next_dived _3192_ vssd1 vssd1 vccd1
+ vccd1 _0210_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6851_ _1396_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5802_ _2247_ _2248_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__nand2_1
X_3994_ pm.count\[4\] vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__inv_2
X_6782_ sound1.sdiv.Q\[9\] _2894_ _2890_ sound1.sdiv.Q\[8\] _2838_ vssd1 vssd1 vccd1
+ vccd1 _0150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5733_ sound4.sdiv.Q\[18\] _2182_ _2185_ sound4.sdiv.Q\[17\] _2197_ vssd1 vssd1 vccd1
+ vccd1 _0018_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5664_ sound4.sdiv.A\[14\] _2144_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7403_ _3560_ _3563_ vssd1 vssd1 vccd1 vccd1 _3565_ sky130_fd_sc_hd__nand2_1
X_4615_ _1026_ _0939_ _1174_ _0990_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_60_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5595_ sound4.sdiv.A\[9\] _2076_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__or2_1
X_7334_ _3500_ _3502_ vssd1 vssd1 vccd1 vccd1 _3503_ sky130_fd_sc_hd__or2_2
XFILLER_0_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4546_ _0990_ _1064_ _1116_ _0994_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7265_ sound3.sdiv.A\[26\] sound3.divisor_m\[0\] vssd1 vssd1 vccd1 vccd1 _3441_ sky130_fd_sc_hd__and2b_1
X_4477_ _0990_ _0996_ _1040_ _0969_ _0943_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__o221a_1
X_6216_ _2648_ _2649_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__or2b_1
X_7196_ sound3.count\[12\] _2863_ vssd1 vssd1 vccd1 vccd1 _3399_ sky130_fd_sc_hd__and2_1
X_6147_ sound4.sdiv.Q\[0\] sound4.sdiv.Q\[1\] _0576_ _2370_ vssd1 vssd1 vccd1 vccd1
+ _2582_ sky130_fd_sc_hd__o211a_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ sound3.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__inv_2
X_5029_ _0698_ _0540_ net44 vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__or3_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4400_ _0674_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__nor2_8
XFILLER_0_124_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5380_ _1778_ _1887_ _1890_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__and3_2
XFILLER_0_1_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4331_ seq.player_7.state\[1\] _0898_ _0901_ seq.player_8.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _0902_ sky130_fd_sc_hd__a22o_1
X_7050_ _3177_ _3308_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__and2_1
X_4262_ seq.clk_div.count\[13\] seq.clk_div.count\[14\] _0838_ vssd1 vssd1 vccd1 vccd1
+ _0844_ sky130_fd_sc_hd__and3_1
X_6001_ sound1.sdiv.Q\[0\] _0579_ _2434_ _2436_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4193_ seq.tempo_select.state\[0\] seq.clk_div.count\[4\] vssd1 vssd1 vccd1 vccd1
+ _0787_ sky130_fd_sc_hd__nand2_1
X_7952_ net130 _0115_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6903_ sound2.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_106_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7883_ net110 net12 net71 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6834_ sound2.count_m\[16\] _2857_ _3131_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6765_ _2005_ _3108_ _3109_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3977_ _0638_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5716_ sound4.count\[2\] _2186_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6696_ _3050_ _3051_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5647_ sound4.sdiv.A\[4\] _2102_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8366_ net119 rate_clk.next_count\[3\] net80 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5578_ _2058_ _2060_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7317_ _3486_ _3487_ vssd1 vssd1 vccd1 vccd1 _3488_ sky130_fd_sc_hd__nand2_1
X_4529_ _0674_ _0687_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8297_ net118 _0397_ net79 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7248_ sound3.divisor_m\[14\] _1628_ _3419_ vssd1 vssd1 vccd1 vccd1 _3430_ sky130_fd_sc_hd__mux2_1
X_7179_ sound3.count_m\[3\] _3132_ _3390_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a21o_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 piano_keys[14] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ wave_comb.u1.start vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4880_ _1034_ _1427_ _1428_ _1430_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__o211a_1
X_3831_ _0507_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__inv_2
XFILLER_0_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6550_ _2419_ _2920_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__xnor2_1
X_3762_ inputcont.INTERNAL_SYNCED_I\[12\] vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5501_ sound4.count\[16\] sound4.count\[17\] _1988_ vssd1 vssd1 vccd1 vccd1 _1995_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6481_ _2869_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8220_ net135 sound3.osc.next_count\[1\] net96 vssd1 vssd1 vccd1 vccd1 sound3.count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_5432_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8151_ net131 _0272_ net92 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[4\] sky130_fd_sc_hd__dfrtp_1
X_5363_ _1107_ _1869_ _1872_ _1873_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7102_ sound2.sdiv.A\[22\] _3329_ vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__xor2_1
X_4314_ _0702_ seq.encode.play _0884_ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1
+ vccd1 vccd1 _0885_ sky130_fd_sc_hd__a31o_1
X_5294_ _1180_ _1786_ _1790_ _1028_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8082_ net119 _0224_ net80 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[17\] sky130_fd_sc_hd__dfrtp_1
X_7033_ _3291_ _3293_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__or2_1
X_4245_ _0831_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_4176_ seq.player_1.state\[2\] seq.player_1.state\[3\] vssd1 vssd1 vccd1 vccd1 _0774_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7935_ net125 _0098_ net86 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[9\] sky130_fd_sc_hd__dfrtp_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7866_ net110 seq.tempo_select.next_state\[1\] net71 vssd1 vssd1 vccd1 vccd1 seq.tempo_select.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6817_ sound2.count\[8\] _2855_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7797_ net118 net8 net79 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_6748_ sound1.sdiv.A\[25\] _3055_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6679_ _2903_ _3036_ vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8349_ net120 sound4.osc.next_count\[7\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4030_ oct.state\[2\] vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__buf_12
XFILLER_0_78_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5981_ sound1.divisor_m\[2\] sound1.count_m\[1\] vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__or2b_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7720_ net137 _0005_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4932_ _0944_ _1336_ _1345_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7651_ _2057_ _2061_ _2141_ vssd1 vssd1 vccd1 vccd1 _3715_ sky130_fd_sc_hd__nand3_1
X_6602_ sound1.divisor_m\[9\] _2967_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__xnor2_1
X_4863_ _1379_ _1388_ _1397_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3814_ _0479_ _0478_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__or2b_1
X_4794_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__buf_4
X_7582_ sound4.divisor_m\[10\] _1803_ _3419_ vssd1 vssd1 vccd1 vccd1 _3669_ sky130_fd_sc_hd__mux2_1
X_6533_ _2902_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6464_ sound1.count_m\[18\] _2857_ _2858_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__a21o_1
X_8203_ net142 _0324_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5415_ _0954_ _1784_ _1790_ _0948_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6395_ _2816_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8134_ net109 _0255_ net70 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[15\] sky130_fd_sc_hd__dfrtp_1
X_5346_ _1095_ _1792_ _1855_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8065_ net117 _0207_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[0\] sky130_fd_sc_hd__dfrtp_1
X_5277_ _0673_ _1773_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__or2_1
X_7016_ _3277_ _3278_ vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__nand2_1
X_4228_ seq.clk_div.count\[4\] seq.clk_div.count\[5\] _0815_ vssd1 vssd1 vccd1 vccd1
+ _0819_ sky130_fd_sc_hd__and3_1
X_4159_ seq.player_2.state\[1\] seq.player_2.state\[2\] seq.player_2.state\[3\] _0762_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__a311o_1
X_7918_ net126 _0081_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7849_ net108 seq.clk_div.next_count\[6\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 piano_keys[3] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6180_ _2613_ _2614_ wave_comb.u1.Q\[2\] _0569_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__a2bb2o_1
X_5200_ sound3.count\[0\] sound3.count\[1\] sound3.count\[2\] sound3.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__and4_1
X_5131_ _1064_ _1565_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__or2_1
X_5062_ _1038_ _1587_ _1589_ _1592_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__o211a_1
X_4013_ _0661_ seq.encode.keys_edge_det\[10\] seq.tempo_select.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _0663_ sky130_fd_sc_hd__or3_1
X_5964_ _2398_ sound1.divisor_m\[6\] sound1.divisor_m\[5\] _2399_ vssd1 vssd1 vccd1
+ vccd1 _2400_ sky130_fd_sc_hd__a22o_1
X_7703_ _2005_ _3749_ _3750_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4915_ _1025_ _1345_ _1462_ _1465_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__o211a_1
X_5895_ sound4.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4846_ sound2.count\[7\] _1368_ _1396_ sound2.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _1397_ sky130_fd_sc_hd__a2bb2o_1
X_7634_ _3702_ _2135_ vssd1 vssd1 vccd1 vccd1 _3703_ sky130_fd_sc_hd__or2b_1
X_7565_ _3659_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6516_ sound1.divisor_m\[0\] sound1.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4777_ _1198_ _1323_ _1327_ _1204_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7496_ sound3.sdiv.C\[1\] sound3.sdiv.C\[0\] sound3.sdiv.C\[2\] vssd1 vssd1 vccd1
+ vccd1 _3644_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6447_ sound1.count\[11\] _2201_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6378_ _0632_ _0643_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8117_ net112 sound2.osc.next_count\[18\] net73 vssd1 vssd1 vccd1 vccd1 sound2.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_5329_ _0959_ _1833_ _1834_ _1835_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__o2111a_1
X_8048_ net112 _0190_ net73 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4700_ sound1.count\[4\] _1263_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__or2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _2159_ _2161_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4631_ _0939_ _1200_ _1189_ _0990_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7350_ sound3.divisor_m\[10\] _3516_ vssd1 vssd1 vccd1 vccd1 _3517_ sky130_fd_sc_hd__xnor2_1
X_4562_ _0674_ _0681_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7281_ sound3.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _3455_ sky130_fd_sc_hd__inv_2
X_6301_ sound3.sdiv.Q\[6\] _0577_ _2731_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4493_ _0674_ _0684_ _0683_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6232_ _2659_ _2663_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6163_ _2439_ _2504_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ sound3.divisor_m\[14\] _2521_ _2529_ sound3.count_m\[14\] vssd1 vssd1 vccd1
+ vccd1 _2530_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5114_ _1015_ _1562_ _1570_ _0952_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__o221a_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _1095_ _1567_ _1570_ _1097_ _1575_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__o221a_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6996_ _3259_ _3260_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5947_ sound1.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7617_ _2110_ _2128_ vssd1 vssd1 vccd1 vccd1 _3691_ sky130_fd_sc_hd__or2_1
X_5878_ sound4.divisor_m\[5\] _2312_ _2313_ sound4.divisor_m\[4\] vssd1 vssd1 vccd1
+ vccd1 _2314_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4829_ _1125_ _1321_ _1327_ _1127_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7548_ sound4.count_m\[9\] _3403_ _2196_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__a21o_1
X_7479_ sound3.sdiv.A\[24\] _3595_ vssd1 vssd1 vccd1 vccd1 _3631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xsass_synth_146 vssd1 vssd1 vccd1 vccd1 sass_synth_146/HI multi[3] sky130_fd_sc_hd__conb_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6850_ _3140_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
X_5801_ wave_comb.u1.A\[7\] _2224_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__or2_1
X_6781_ sound1.sdiv.Q\[8\] _2894_ _2890_ sound1.sdiv.Q\[7\] _2837_ vssd1 vssd1 vccd1
+ vccd1 _0149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3993_ _0649_ _0650_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_91_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5732_ sound4.count\[10\] _2186_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7402_ _3560_ _3563_ vssd1 vssd1 vccd1 vccd1 _3564_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4614_ _0958_ _1141_ _1179_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5594_ sound4.sdiv.A\[9\] _2076_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7333_ sound3.divisor_m\[8\] _3501_ vssd1 vssd1 vccd1 vccd1 _3502_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4545_ _0695_ net64 _1040_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7264_ _3437_ _3438_ _3439_ _3440_ sound3.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _0306_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4476_ _0950_ _0996_ _1046_ _0994_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7195_ sound3.count_m\[11\] _3132_ _3398_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6215_ _2645_ _2647_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6146_ wave_comb.u1.next_start _2580_ _2581_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__a21o_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ sound3.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__inv_2
X_5028_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__buf_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ sound2.divisor_m\[9\] sound2.divisor_m\[8\] sound2.divisor_m\[7\] _3221_ vssd1
+ vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ select1.sequencer_on _0897_ _0899_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a31oi_2
X_4261_ _0843_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6000_ _2435_ sound1.sdiv.next_start vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4192_ seq.tempo_select.state\[0\] _0781_ _0784_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_
+ sky130_fd_sc_hd__o22ai_1
X_7951_ net131 _0114_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7882_ net108 net11 net69 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6902_ sound2.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__inv_2
X_6833_ sound2.count\[16\] _2855_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6764_ _0565_ _3106_ sound1.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3976_ inputcont.INTERNAL_SYNCED_I\[9\] _0624_ _0622_ vssd1 vssd1 vccd1 vccd1 _0639_
+ sky130_fd_sc_hd__a21oi_1
X_6695_ _3050_ _3051_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5715_ sound4.sdiv.Q\[9\] _2184_ _2185_ sound4.sdiv.Q\[8\] _2188_ vssd1 vssd1 vccd1
+ vccd1 _0009_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5646_ _2110_ _2128_ _2107_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8365_ net118 rate_clk.next_count\[2\] net79 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5577_ sound4.divisor_m\[13\] _2059_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7316_ _3482_ _3485_ vssd1 vssd1 vccd1 vccd1 _3487_ sky130_fd_sc_hd__nand2_1
X_4528_ _0939_ _1095_ _1056_ _0958_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8296_ net122 _0396_ net83 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[10\] sky130_fd_sc_hd__dfrtp_4
X_7247_ _3429_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_1
X_4459_ _1000_ _1025_ _1027_ _0976_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__o221a_1
X_7178_ sound3.count\[3\] _2863_ vssd1 vssd1 vccd1 vccd1 _3390_ sky130_fd_sc_hd__and2_1
X_6129_ _2564_ _2530_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__or2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nor2b_2
X_3761_ inputcont.INTERNAL_SYNCED_I\[9\] inputcont.INTERNAL_SYNCED_I\[8\] _0443_ _0444_
+ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__or4_4
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5500_ _1994_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ sound1.divisor_m\[5\] _1186_ _2864_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5431_ sound4.count\[0\] sound4.count\[1\] sound4.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1940_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8150_ net131 _0271_ net92 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[3\] sky130_fd_sc_hd__dfrtp_1
X_5362_ _0677_ _1083_ _1784_ _1777_ _1064_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__o32a_1
XFILLER_0_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8081_ net116 _0223_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[16\] sky130_fd_sc_hd__dfrtp_1
X_7101_ _3349_ _3353_ _3354_ _3174_ sound2.sdiv.A\[22\] vssd1 vssd1 vccd1 vccd1 _0229_
+ sky130_fd_sc_hd__a32o_1
X_4313_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__and3b_1
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7032_ sound2.divisor_m\[15\] _3292_ vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__xnor2_1
X_5293_ sound4.count\[10\] _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4244_ _0829_ _0813_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__and3b_1
X_4175_ seq.player_1.state\[2\] seq.player_1.state\[3\] _0772_ _0773_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_1.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7934_ net127 _0097_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[8\] sky130_fd_sc_hd__dfrtp_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7865_ net110 seq.tempo_select.next_state\[0\] net71 vssd1 vssd1 vccd1 vccd1 seq.tempo_select.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_7796_ net138 net7 net99 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6816_ sound2.count_m\[7\] _2857_ _3122_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__a21o_1
X_6747_ sound1.sdiv.A\[25\] _3055_ vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3959_ inputcont.INTERNAL_SYNCED_I\[7\] _0621_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nor2_1
X_6678_ sound1.divisor_m\[16\] _3028_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5629_ sound4.divisor_m\[2\] sound4.divisor_m\[1\] sound4.divisor_m\[0\] _2036_ vssd1
+ vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8348_ net120 sound4.osc.next_count\[6\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_8279_ net122 _0379_ net83 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5980_ sound1.count_m\[1\] sound1.divisor_m\[2\] vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4931_ _1035_ _1323_ _1322_ _1039_ _1481_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__o221a_1
X_4862_ sound2.count\[1\] _1404_ _1412_ sound2.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _1413_ sky130_fd_sc_hd__a2bb2o_1
X_7650_ sound4.sdiv.A\[13\] _2183_ sound4.sdiv.next_dived _3714_ vssd1 vssd1 vccd1
+ vccd1 _0418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6601_ _2395_ _2957_ sound1.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ inputcont.INTERNAL_SYNCED_I\[10\] _0445_ _0488_ _0491_ vssd1 vssd1 vccd1 vccd1
+ _0492_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4793_ _1331_ _1334_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__or2_1
X_7581_ _2005_ _1840_ _3668_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6532_ sound1.divisor_m\[2\] _2904_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6463_ sound1.count\[18\] _2855_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8202_ net142 _0323_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5414_ sound4.count\[12\] _1924_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__xor2_1
X_6394_ _2623_ _2655_ _2805_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8133_ net109 _0254_ net70 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5345_ _0993_ _1012_ _1790_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8064_ net117 _0206_ net78 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[18\] sky130_fd_sc_hd__dfrtp_1
X_5276_ _1125_ _1784_ _1786_ _1127_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__o22a_1
X_7015_ _3273_ _3276_ vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__nand2_1
X_4227_ seq.clk_div.count\[4\] _0815_ _0818_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
X_4158_ seq.player_2.state\[0\] _0761_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__and2_1
X_4089_ seq.player_8.state\[1\] _0713_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__nor2_1
X_7917_ net126 _0080_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7848_ net108 seq.clk_div.next_count\[5\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_7779_ net139 _0053_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 piano_keys[4] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5130_ _0687_ _1001_ _1578_ _1572_ _1116_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__o32a_1
XFILLER_0_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5061_ _1026_ _1559_ _1572_ _1064_ _1591_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__o221a_1
X_4012_ _0661_ seq.encode.keys_edge_det\[10\] seq.tempo_select.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _0662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5963_ sound1.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__inv_2
X_7702_ _0556_ _3747_ sound4.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 _3750_ sky130_fd_sc_hd__a21oi_1
X_4914_ _1005_ _1338_ _1336_ _1027_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__o221a_1
X_5894_ sound4.divisor_m\[13\] _2324_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4845_ _1390_ _1392_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7633_ _2136_ _2083_ vssd1 vssd1 vccd1 vccd1 _3702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7564_ sound4.divisor_m\[2\] _3658_ _3419_ vssd1 vssd1 vccd1 vccd1 _3659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4776_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6515_ _0867_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__buf_8
XFILLER_0_99_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7495_ _1545_ vssd1 vssd1 vccd1 vccd1 _3643_ sky130_fd_sc_hd__clkbuf_8
X_6446_ sound1.count_m\[10\] _2836_ _2848_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6377_ wave_comb.u1.Q\[11\] _0573_ wave_comb.u1.next_dived wave_comb.u1.Q\[10\] vssd1
+ vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8116_ net112 sound2.osc.next_count\[17\] net73 vssd1 vssd1 vccd1 vccd1 sound2.count\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_5328_ _1077_ _1769_ _1836_ _1838_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__o211a_1
X_8047_ net111 _0189_ net72 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[1\] sky130_fd_sc_hd__dfrtp_4
X_5259_ _0673_ _1765_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4630_ _0686_ _0950_ _0994_ _1146_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6300_ sound3.sdiv.Q\[5\] _2632_ _2699_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__a21o_1
X_4561_ _0967_ _1123_ _1125_ _0958_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7280_ _3447_ _3450_ vssd1 vssd1 vccd1 vccd1 _3454_ sky130_fd_sc_hd__or2_1
X_4492_ _0964_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6231_ _2659_ _2663_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6162_ _2439_ _2504_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5113_ _1079_ _1580_ _1574_ _0680_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ sound3.divisor_m\[15\] vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__inv_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _1572_ _1574_ _0960_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__a21o_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6995_ _3255_ _3258_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5946_ sound1.count_m\[15\] _2381_ sound1.count_m\[14\] _2375_ vssd1 vssd1 vccd1
+ vccd1 _2382_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5877_ sound4.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7616_ _3689_ vssd1 vssd1 vccd1 vccd1 _3690_ sky130_fd_sc_hd__inv_2
X_4828_ sound2.count\[6\] _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4759_ _0575_ _0560_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nor2_4
X_7547_ sound4.count_m\[8\] _3403_ _2195_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a21o_1
X_7478_ sound3.sdiv.A\[24\] _3595_ vssd1 vssd1 vccd1 vccd1 _3630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6429_ sound1.count_m\[2\] _2836_ _2839_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3992_ pm.count\[3\] _0647_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__nor2_1
X_5800_ wave_comb.u1.A\[7\] _2224_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__nand2_1
X_6780_ sound1.sdiv.Q\[7\] _2894_ _2890_ sound1.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1
+ _0148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5731_ sound4.sdiv.Q\[17\] _2182_ _2185_ sound4.sdiv.Q\[16\] _2196_ vssd1 vssd1 vccd1
+ vccd1 _0017_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5662_ sound4.sdiv.A\[14\] _2144_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__nand2_1
X_7401_ sound3.divisor_m\[15\] _3562_ vssd1 vssd1 vccd1 vccd1 _3563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4613_ _0969_ _1180_ _1181_ _0967_ _1183_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5593_ _2075_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7332_ sound3.divisor_m\[7\] _3492_ _3448_ vssd1 vssd1 vccd1 vccd1 _3501_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4544_ _0976_ _1112_ _1113_ _1000_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7263_ _0577_ vssd1 vssd1 vccd1 vccd1 _3440_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6214_ _2645_ _2647_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__nor2_1
X_4475_ _0674_ _0945_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nor2_4
X_7194_ sound3.count\[11\] _2863_ vssd1 vssd1 vccd1 vccd1 _3398_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6145_ wave_comb.u1.Q\[2\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ sound3.divisor_m\[5\] _2511_ _2508_ sound3.divisor_m\[4\] vssd1 vssd1 vccd1
+ vccd1 _2512_ sky130_fd_sc_hd__o22a_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _1556_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__or2_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6978_ sound2.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5929_ _2364_ _2332_ _2342_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _0841_ _0813_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4191_ seq.tempo_select.state\[0\] seq.tempo_select.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7950_ net130 _0113_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6901_ _3170_ sound2.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__or2b_1
X_7881_ net118 net10 net79 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_6832_ sound2.count_m\[15\] _2857_ _3130_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6763_ sound1.sdiv.C\[3\] _0565_ _3106_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3975_ _0633_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6694_ _3041_ _3043_ _3040_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__a21boi_1
X_5714_ sound4.count\[1\] _2186_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5645_ _2116_ _2127_ _2114_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8364_ net118 rate_clk.next_count\[1\] net79 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5576_ _2036_ _2032_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__and2_1
X_7315_ _3482_ _3485_ vssd1 vssd1 vccd1 vccd1 _3486_ sky130_fd_sc_hd__or2_1
X_4527_ _0969_ _1096_ _1097_ _1000_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8295_ net122 _0395_ net83 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[9\] sky130_fd_sc_hd__dfrtp_2
X_7246_ sound3.divisor_m\[13\] _1667_ _3419_ vssd1 vssd1 vccd1 vccd1 _3429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4458_ _0969_ _1025_ _1028_ _1005_ _0943_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__o32a_1
X_7177_ sound3.count_m\[2\] _3132_ _3389_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__a21o_1
X_6128_ _2562_ _2527_ _2528_ _2563_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__o31a_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ _0959_ _0944_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__or2_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _2474_ sound2.divisor_m\[4\] _2476_ _2494_ _2469_ vssd1 vssd1 vccd1 vccd1
+ _2495_ sky130_fd_sc_hd__o221a_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3760_ inputcont.INTERNAL_SYNCED_I\[5\] inputcont.INTERNAL_SYNCED_I\[4\] inputcont.INTERNAL_SYNCED_I\[7\]
+ inputcont.INTERNAL_SYNCED_I\[6\] vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__or4_4
XFILLER_0_82_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5430_ _1939_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _0997_ _1792_ _1796_ _1112_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8080_ net116 _0222_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7100_ _3351_ _3352_ _3350_ vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__a21o_1
X_5292_ _1053_ _1781_ _1787_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__o211ai_4
X_4312_ _0881_ _0882_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__nand2_1
X_7031_ sound2.divisor_m\[14\] _3283_ _3177_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__o21a_1
X_4243_ seq.clk_div.count\[8\] _0824_ seq.clk_div.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _0830_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4174_ seq.player_1.state\[1\] _0770_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7933_ net127 _0096_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[7\] sky130_fd_sc_hd__dfrtp_2
X_7864_ net110 seq.clk_div.next_count\[21\] net71 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7795_ net110 net6 net71 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_6815_ sound2.count\[7\] _2855_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__and2_1
X_6746_ sound1.sdiv.A\[25\] _2895_ sound1.sdiv.next_dived _3095_ vssd1 vssd1 vccd1
+ vccd1 _0133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3958_ inputcont.INTERNAL_SYNCED_I\[7\] _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__and2_1
X_6677_ _2890_ _3034_ _3035_ _2894_ sound1.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 _0124_
+ sky130_fd_sc_hd__a32o_1
X_3889_ sound2.sdiv.C\[4\] sound2.sdiv.C\[3\] sound2.sdiv.C\[2\] _0558_ sound2.sdiv.C\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__a311oi_4
X_5628_ sound4.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5559_ _2040_ _2041_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__or2_1
X_8347_ net121 sound4.osc.next_count\[5\] net82 vssd1 vssd1 vccd1 vccd1 sound4.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_8278_ net118 _0378_ net79 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7229_ _3418_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__clkbuf_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4930_ _1043_ _1339_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__or2_1
X_4861_ _1405_ _1408_ _1411_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6600_ _2960_ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3812_ _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__clkbuf_4
X_4792_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__buf_4
X_7580_ sound4.divisor_m\[9\] _2005_ vssd1 vssd1 vccd1 vccd1 _3668_ sky130_fd_sc_hd__nor2_1
X_6531_ sound1.divisor_m\[1\] sound1.divisor_m\[0\] _2903_ vssd1 vssd1 vccd1 vccd1
+ _2904_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6462_ _0554_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__buf_6
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8201_ net142 _0322_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[16\] sky130_fd_sc_hd__dfrtp_1
X_6393_ _2815_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
X_5413_ _1079_ _1842_ _1919_ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__a211o_2
XFILLER_0_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8132_ net112 _0253_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[13\] sky130_fd_sc_hd__dfrtp_1
X_5344_ _0977_ _0996_ _1784_ _1854_ _0960_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__o32a_1
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8063_ net117 _0205_ net78 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[17\] sky130_fd_sc_hd__dfrtp_2
X_5275_ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7014_ _3273_ _3276_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__or2_1
X_4226_ seq.clk_div.count\[4\] _0815_ _0813_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__o21ai_1
X_4157_ _0449_ seq.encode.keys_edge_det\[3\] vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4088_ seq.player_8.state\[0\] seq.player_8.state\[1\] _0712_ vssd1 vssd1 vccd1 vccd1
+ _0715_ sky130_fd_sc_hd__and3_1
X_7916_ net126 _0079_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7847_ net108 seq.clk_div.next_count\[4\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ net139 _0052_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6729_ sound1.sdiv.A\[22\] _3055_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 piano_keys[5] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5060_ _1556_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__or2_4
X_4011_ seq.encode.keys_sync\[10\] vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__inv_2
X_5962_ sound1.count_m\[5\] vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7701_ sound4.sdiv.C\[3\] _0556_ _3747_ vssd1 vssd1 vccd1 vccd1 _3749_ sky130_fd_sc_hd__and3_1
X_4913_ _0997_ _1323_ _1343_ _1010_ _1463_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__o221a_1
X_5893_ _2326_ sound4.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4844_ _0985_ _1322_ _1339_ _1181_ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7632_ _3700_ _3701_ sound4.sdiv.A\[8\] _2183_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_62_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7563_ _1903_ vssd1 vssd1 vccd1 vccd1 _3658_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4775_ _0499_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__or2_1
X_6514_ _2889_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7494_ _3437_ _3641_ _3642_ _3440_ sound3.sdiv.C\[1\] vssd1 vssd1 vccd1 vccd1 _0334_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6445_ sound1.count\[10\] _2201_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6376_ _0645_ _2801_ _2802_ _2803_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8115_ net112 sound2.osc.next_count\[16\] net73 vssd1 vssd1 vccd1 vccd1 sound2.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_5327_ _1020_ _1777_ _1792_ _1014_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__o221a_1
X_8046_ net111 _0188_ net72 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[0\] sky130_fd_sc_hd__dfrtp_4
X_5258_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5189_ _1621_ _1719_ _1591_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__o21a_1
X_4209_ seq.clk_div.count\[7\] seq.clk_div.count\[11\] _0802_ seq.clk_div.count\[21\]
+ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire60 _2541_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4560_ _0992_ _1126_ _1127_ _0990_ _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__o221a_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4491_ _0676_ _0685_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6230_ sound2.sdiv.Q\[5\] _2295_ _2662_ _2292_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6161_ _2590_ _2595_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5112_ net64 _1077_ _1567_ _1553_ _0946_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__o32a_1
XFILLER_0_20_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ sound3.divisor_m\[13\] _2522_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5043_ _1573_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__buf_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6994_ _3255_ _3258_ vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__nor2_1
X_5945_ sound1.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__inv_2
X_5876_ sound4.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7615_ _2110_ _2128_ vssd1 vssd1 vccd1 vccd1 _3689_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4827_ _0983_ _1338_ _1371_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4758_ _1310_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7546_ sound4.count_m\[7\] _3403_ _2194_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__a21o_1
X_7477_ _3621_ _3627_ _3622_ vssd1 vssd1 vccd1 vccd1 _3629_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4689_ _1256_ _1257_ _1258_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6428_ sound1.count\[2\] _2201_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6359_ wave_comb.u1.Q\[7\] _0569_ _2787_ _2788_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__a22o_1
X_8029_ net111 _0171_ net72 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3991_ pm.count\[3\] _0647_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5730_ sound4.count\[9\] _2186_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7400_ _3448_ _3561_ vssd1 vssd1 vccd1 vccd1 _3562_ sky130_fd_sc_hd__and2_1
X_5661_ sound4.divisor_m\[15\] _2143_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4612_ _1182_ _1000_ _1003_ _0985_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5592_ sound4.divisor_m\[10\] _2074_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__xnor2_1
X_7331_ sound3.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 _3500_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4543_ _0687_ _1001_ _0943_ _0997_ _0939_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o32a_1
XFILLER_0_53_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7262_ sound3.divisor_m\[0\] sound3.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3439_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6213_ _2585_ _2606_ _2646_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__a21oi_1
X_4474_ _1003_ _1039_ _1041_ _0939_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7193_ sound3.count_m\[10\] _3132_ _3397_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6144_ wave_comb.u1.Q\[1\] _0569_ _2578_ _2579_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__a22o_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ sound3.count_m\[4\] vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__inv_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _0698_ net56 vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _3164_ _3242_ _3243_ _3174_ sound2.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 _0216_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5928_ _2362_ _2329_ _2330_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__o31a_1
X_5859_ _2276_ _2292_ _2295_ sound2.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7529_ sound3.sdiv.Q\[18\] _3654_ _3643_ sound3.sdiv.Q\[17\] _3397_ vssd1 vssd1 vccd1
+ vccd1 _0357_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ seq.clk_div.count\[19\] _0782_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__a21oi_1
X_7880_ net130 net4 net91 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6900_ _3164_ _3172_ _3173_ _3174_ sound2.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _0208_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6831_ sound2.count\[15\] _2855_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6762_ _2890_ _3105_ _3107_ _2894_ sound1.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3974_ _0634_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6693_ _3048_ _3049_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__nand2_1
X_5713_ sound4.sdiv.Q\[8\] _2184_ _2185_ sound4.sdiv.Q\[7\] _2187_ vssd1 vssd1 vccd1
+ vccd1 _0008_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5644_ _2120_ _2125_ _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8363_ net118 rate_clk.next_count\[0\] net79 vssd1 vssd1 vccd1 vccd1 rate_clk.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7314_ sound3.divisor_m\[6\] _3484_ vssd1 vssd1 vccd1 vccd1 _3485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5575_ sound4.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4526_ _0952_ _0972_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__nor2_2
X_8294_ net123 _0394_ net84 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7245_ _3428_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
X_4457_ _0695_ _0946_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nor2_8
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7176_ sound3.count\[2\] _2863_ vssd1 vssd1 vccd1 vccd1 _3389_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6127_ _2523_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__inv_2
X_4388_ _0951_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__buf_8
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _2481_ _2483_ _2475_ sound2.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2494_
+ sky130_fd_sc_hd__o2bb2a_1
X_5009_ sound2.count\[18\] _1539_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__or2_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5360_ _1016_ _1786_ _1781_ _1116_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5291_ _1012_ _1790_ _1798_ _1801_ _1778_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__o2111a_1
X_4311_ seq.player_3.state\[0\] seq.player_3.state\[1\] seq.player_3.state\[2\] seq.player_3.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7030_ sound2.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__inv_2
X_4242_ seq.clk_div.count\[8\] seq.clk_div.count\[9\] _0824_ vssd1 vssd1 vccd1 vccd1
+ _0829_ sky130_fd_sc_hd__and3_1
X_4173_ seq.player_1.state\[0\] seq.player_1.state\[1\] _0769_ vssd1 vssd1 vccd1 vccd1
+ _0772_ sky130_fd_sc_hd__and3_1
X_7932_ net127 _0095_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7863_ net110 seq.clk_div.next_count\[20\] net71 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7794_ net139 net5 net100 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6814_ sound2.count_m\[6\] _2857_ _3121_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a21o_1
X_6745_ _3091_ _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__xnor2_1
X_3957_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6676_ _3022_ _3026_ _3033_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__a21o_1
X_3888_ sound2.sdiv.start vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5627_ _2109_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__inv_2
X_5558_ sound4.sdiv.A\[19\] _2038_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8346_ net120 sound4.osc.next_count\[4\] net81 vssd1 vssd1 vccd1 vccd1 sound4.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4509_ _0956_ _1078_ _1079_ _0992_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8277_ net118 _0377_ net79 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[10\] sky130_fd_sc_hd__dfrtp_1
X_7228_ sound3.divisor_m\[6\] _1594_ _3142_ vssd1 vssd1 vccd1 vccd1 _3418_ sky130_fd_sc_hd__mux2_1
X_5489_ sound4.count\[12\] sound4.count\[13\] _1973_ sound4.count\[14\] vssd1 vssd1
+ vccd1 vccd1 _1986_ sky130_fd_sc_hd__a31o_1
X_7159_ sound2.sdiv.Q\[15\] _3167_ _3349_ sound2.sdiv.Q\[14\] _3122_ vssd1 vssd1 vccd1
+ vccd1 _0255_ sky130_fd_sc_hd__a221o_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4860_ _1317_ _1409_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__and3_1
X_3811_ _0479_ _0478_ _0485_ _0489_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6530_ sound1.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4791_ net40 _1330_ _1324_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6461_ sound1.count_m\[17\] _2836_ _2856_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8200_ net142 _0321_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6392_ pm.current_waveform\[3\] _2814_ _2808_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5412_ _1025_ _1920_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8131_ net112 _0252_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _1780_ _1832_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5274_ _0719_ _0587_ _0672_ _0673_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__or4_2
X_8062_ net116 _0204_ net77 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[16\] sky130_fd_sc_hd__dfrtp_1
X_7013_ sound2.divisor_m\[13\] _3275_ vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__xnor2_1
X_4225_ _0817_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_4156_ _0758_ _0757_ _0760_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_3.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4087_ seq.player_8.state\[0\] _0712_ _0714_ vssd1 vssd1 vccd1 vccd1 seq.player_8.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_7915_ net126 _0078_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[8\] sky130_fd_sc_hd__dfrtp_1
X_7846_ net108 seq.clk_div.next_count\[3\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7777_ net139 _0051_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[6\] sky130_fd_sc_hd__dfrtp_1
X_4989_ _1527_ _1528_ _1504_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__and3b_1
X_6728_ _3079_ _3080_ sound1.sdiv.A\[22\] _2895_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6659_ sound1.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8329_ net124 _0429_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 piano_keys[6] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4010_ wave.mode\[1\] _0659_ vssd1 vssd1 vccd1 vccd1 wave.next_state\[1\] sky130_fd_sc_hd__xor2_1
X_5961_ sound1.count_m\[7\] _2395_ _2396_ sound1.divisor_m\[7\] vssd1 vssd1 vccd1
+ vccd1 _2397_ sky130_fd_sc_hd__a2bb2o_1
X_7700_ _3681_ _3746_ _3748_ _2184_ sound4.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 _0434_
+ sky130_fd_sc_hd__a32o_1
X_4912_ _1020_ _1347_ _1333_ _0973_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5892_ _2326_ sound4.divisor_m\[12\] _2327_ sound4.divisor_m\[11\] vssd1 vssd1 vccd1
+ vccd1 _2328_ sky130_fd_sc_hd__a22o_1
X_7631_ _2089_ _2134_ _1764_ vssd1 vssd1 vccd1 vccd1 _3701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4843_ _1026_ _1343_ _1333_ _1174_ _1393_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7562_ _3657_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4774_ _0504_ _1324_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__or2_2
X_7493_ sound3.sdiv.C\[1\] sound3.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3642_ sky130_fd_sc_hd__or2_1
X_6513_ sound1.divisor_m\[18\] _1223_ _2864_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6444_ sound1.count_m\[9\] _2836_ _2847_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6375_ _2796_ net53 vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8114_ net112 sound2.osc.next_count\[15\] net73 vssd1 vssd1 vccd1 vccd1 sound2.count\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_5326_ _1158_ _1790_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__or2_1
X_8045_ net120 _0187_ net81 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[18\] sky130_fd_sc_hd__dfrtp_1
X_5257_ _1765_ _1767_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__or2_1
X_4208_ seq.clk_div.count\[13\] vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__inv_2
X_5188_ _1629_ _1657_ _1692_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4139_ seq.player_4.state\[2\] seq.player_4.state\[3\] _0748_ _0749_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_4.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire61 net62 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7829_ net113 seq.player_2.next_state\[3\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4490_ _0939_ _1057_ _1058_ _0958_ _1060_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6160_ _2292_ _2592_ _2593_ _2594_ _2279_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__o32ai_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5111_ sound3.count\[7\] vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__inv_2
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _2524_ sound3.divisor_m\[12\] vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__nor2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5042_ _1560_ _1568_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__or2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6993_ sound2.divisor_m\[11\] _3257_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__xnor2_1
X_5944_ sound1.count_m\[10\] _2378_ _2379_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5875_ _2306_ _2307_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7614_ _3681_ _3687_ _3688_ _2184_ sound4.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _0408_
+ sky130_fd_sc_hd__a32o_1
X_4826_ _0676_ _1372_ _1373_ _1375_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7545_ sound4.count_m\[6\] _3403_ _2193_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__a21o_1
X_4757_ _1256_ _1308_ _1309_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7476_ sound3.sdiv.A\[24\] _3463_ sound3.sdiv.next_dived _3628_ vssd1 vssd1 vccd1
+ vccd1 _0330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4688_ sound1.count\[0\] sound1.count\[1\] vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6427_ sound1.count_m\[1\] _2836_ _2838_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6358_ _2783_ _2786_ _0569_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__a21oi_1
X_5309_ _1010_ _1772_ _1778_ _1819_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__o211a_1
X_6289_ sound2.sdiv.Q\[6\] _0578_ _2718_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__a21o_1
X_8028_ net120 _0170_ net81 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ _0647_ _0648_ vssd1 vssd1 vccd1 vccd1 pm.next_count\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_0_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _2142_ _2054_ sound4.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4611_ _0959_ _0944_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5591_ _2036_ _2030_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__and2_1
X_7330_ _3437_ _3498_ _3499_ _3440_ sound3.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 _0313_
+ sky130_fd_sc_hd__a32o_1
X_4542_ _1015_ _1062_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7261_ sound3.divisor_m\[0\] sound3.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3438_ sky130_fd_sc_hd__nand2_1
X_4473_ _0958_ _1042_ _1043_ _0967_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6212_ _2605_ _2600_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7192_ sound3.count\[10\] _2863_ vssd1 vssd1 vccd1 vccd1 _3397_ sky130_fd_sc_hd__and2_1
X_6143_ _2311_ _2577_ _0569_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__a21oi_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _2508_ sound3.divisor_m\[4\] _2509_ sound3.divisor_m\[3\] vssd1 vssd1 vccd1
+ vccd1 _2510_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _1555_ _1546_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__or2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6976_ _3233_ _3237_ _3240_ _3241_ vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__a211o_1
X_5927_ _2325_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5858_ sound2.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5789_ wave_comb.u1.A\[5\] _2224_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4809_ _1354_ _1356_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__and3_2
X_7528_ sound3.sdiv.Q\[17\] _3654_ _3643_ sound3.sdiv.Q\[16\] _3396_ vssd1 vssd1 vccd1
+ vccd1 _0356_ sky130_fd_sc_hd__a221o_1
X_7459_ sound3.sdiv.A\[20\] sound3.sdiv.A\[19\] _3595_ vssd1 vssd1 vccd1 vccd1 _3614_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6830_ sound2.count_m\[14\] _2857_ _3129_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__a21o_1
X_6761_ _3106_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5712_ sound4.count\[0\] _2186_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ inputcont.INTERNAL_SYNCED_I\[11\] _0635_ _0619_ vssd1 vssd1 vccd1 vccd1 _0636_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6692_ _3045_ _3047_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5643_ _2117_ _2119_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8362_ net145 wave.next_state\[1\] net106 vssd1 vssd1 vccd1 vccd1 wave.mode\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5574_ sound4.sdiv.A\[13\] _2056_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__xnor2_1
X_7313_ _3448_ _3483_ vssd1 vssd1 vccd1 vccd1 _3484_ sky130_fd_sc_hd__and2_1
X_4525_ _0983_ _0978_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__or2_2
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8293_ net122 _0393_ net83 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[7\] sky130_fd_sc_hd__dfrtp_2
X_7244_ sound3.divisor_m\[12\] _3427_ _3419_ vssd1 vssd1 vccd1 vccd1 _3428_ sky130_fd_sc_hd__mux2_1
X_4456_ _0964_ _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nand2_2
X_7175_ sound3.count_m\[1\] _3132_ _3388_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__a21o_1
X_4387_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__buf_4
X_6126_ _2533_ _2561_ _2526_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__a21oi_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6057_ _2467_ _2492_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5008_ _1541_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6959_ _3215_ _3219_ _3226_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _1151_ _1769_ _1800_ _0983_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4310_ select1.sequencer_on _0880_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _0828_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_4172_ seq.player_1.state\[0\] _0769_ _0771_ vssd1 vssd1 vccd1 vccd1 seq.player_1.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_117_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7931_ net127 _0094_ net88 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[5\] sky130_fd_sc_hd__dfrtp_2
X_7862_ net110 seq.clk_div.next_count\[19\] net71 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_7793_ net130 net18 net91 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6813_ sound2.count\[6\] _2855_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6744_ _3092_ _3093_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__and2_1
X_3956_ _0611_ _0618_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6675_ _3022_ _3026_ _3033_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__nand3_1
XFILLER_0_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3887_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__inv_2
X_5626_ _2107_ _2108_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5557_ sound4.sdiv.A\[20\] _2038_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__xnor2_1
X_8345_ net121 sound4.osc.next_count\[3\] net82 vssd1 vssd1 vccd1 vccd1 sound4.count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_4508_ _0970_ _0869_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nand2_4
X_8276_ net122 _0376_ net83 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[9\] sky130_fd_sc_hd__dfrtp_1
X_5488_ _1984_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7227_ _3417_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_1
X_4439_ _0685_ _0681_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__nand2_8
X_7158_ sound2.sdiv.Q\[14\] _3167_ _3349_ sound2.sdiv.Q\[13\] _3121_ vssd1 vssd1 vccd1
+ vccd1 _0254_ sky130_fd_sc_hd__a221o_1
X_6109_ sound3.count_m\[16\] vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__inv_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _3342_ _3344_ sound2.sdiv.A\[20\] _3168_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3810_ inputcont.INTERNAL_SYNCED_I\[6\] _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__o31ai_2
X_4790_ _1340_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ sound1.count\[17\] _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6391_ _2590_ _2616_ _2805_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5411_ _1245_ _1800_ _1796_ _1110_ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8130_ net112 _0251_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[11\] sky130_fd_sc_hd__dfrtp_1
X_5342_ _1096_ _1786_ _1794_ _1097_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__o22a_1
X_8061_ net116 _0203_ net77 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7012_ _3177_ _3274_ vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__and2_1
X_5273_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__buf_4
X_4224_ _0815_ _0816_ _0813_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__and3b_1
X_4155_ seq.player_3.state\[1\] seq.player_3.state\[2\] _0754_ seq.player_3.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__a31o_1
X_4086_ seq.player_8.state\[1\] seq.player_8.state\[2\] seq.player_8.state\[3\] _0713_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a311o_1
X_7914_ net127 _0077_ net88 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7845_ net108 seq.clk_div.next_count\[2\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7776_ net139 _0050_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[5\] sky130_fd_sc_hd__dfrtp_1
X_4988_ sound2.count\[10\] _1524_ sound2.count\[11\] vssd1 vssd1 vccd1 vccd1 _1528_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6727_ _3078_ _3076_ _3077_ _0866_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3939_ _0587_ _0597_ _0596_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6658_ _2890_ _3017_ _3018_ _2894_ sound1.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _0122_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5609_ _2091_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__inv_2
X_6589_ sound1.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__inv_2
X_8328_ net138 _0428_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[23\] sky130_fd_sc_hd__dfrtp_1
X_8259_ net132 _0359_ net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[20\] sky130_fd_sc_hd__dfrtp_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 piano_keys[7] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5960_ sound1.count_m\[6\] vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__inv_2
X_5891_ sound4.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__inv_2
X_4911_ _1017_ _1321_ _1341_ _1016_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7630_ _2089_ _2134_ vssd1 vssd1 vccd1 vccd1 _3700_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4842_ _0996_ _1321_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7561_ sound4.divisor_m\[1\] _3656_ _3419_ vssd1 vssd1 vccd1 vccd1 _3657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4773_ _0698_ _0507_ net42 vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__or3_2
X_7492_ sound3.sdiv.C\[1\] sound3.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6512_ _2888_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6443_ sound1.count\[9\] _2201_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6374_ _0569_ _2794_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8113_ net110 sound2.osc.next_count\[14\] net71 vssd1 vssd1 vccd1 vccd1 sound2.count\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_5325_ _1028_ _1800_ _1794_ _1083_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8044_ net117 _0186_ net78 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[17\] sky130_fd_sc_hd__dfrtp_1
X_5256_ _0673_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4207_ _0796_ _0797_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5187_ sound3.count\[11\] _1699_ _1707_ _1716_ _1717_ vssd1 vssd1 vccd1 vccd1 _1718_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4138_ seq.player_4.state\[1\] _0746_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nor2_1
X_4069_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire62 _2344_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7828_ net113 seq.player_2.next_state\[2\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7759_ net143 _0044_ net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6090_ _2524_ sound3.divisor_m\[12\] _2525_ sound3.divisor_m\[11\] vssd1 vssd1 vccd1
+ vccd1 _2526_ sky130_fd_sc_hd__a22o_1
X_5110_ _0688_ _1559_ _1578_ _1014_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__o221a_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _1571_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__buf_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6992_ _3177_ _3256_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__and2_1
X_5943_ sound1.divisor_m\[10\] sound1.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2379_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ wave_comb.u1.next_start _2309_ _2310_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7613_ _2116_ _2127_ vssd1 vssd1 vccd1 vccd1 _3688_ sky130_fd_sc_hd__nand2_1
X_4825_ _0677_ _1038_ _1336_ _1339_ _1026_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7544_ sound4.count_m\[5\] _3403_ _2192_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4756_ sound1.count\[18\] _1305_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7475_ _3623_ _3627_ vssd1 vssd1 vccd1 vccd1 _3628_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4687_ sound1.count\[0\] sound1.count\[1\] vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__or2_1
X_6426_ sound1.count\[1\] _2201_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6357_ _2783_ _2786_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__or2_1
X_5308_ _1773_ _1777_ _1055_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__a21o_1
X_6288_ sound2.sdiv.Q\[6\] _2718_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__nand2_1
X_5239_ _1753_ _1754_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[15\] sky130_fd_sc_hd__nor2_1
X_8027_ net120 _0169_ net81 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4610_ _0952_ _1004_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5590_ _2070_ _2072_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4541_ _1015_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nand2_4
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7260_ _1545_ vssd1 vssd1 vccd1 vccd1 _3437_ sky130_fd_sc_hd__buf_6
X_4472_ _0679_ _0944_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nor2_2
XFILLER_0_123_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7191_ sound3.count_m\[9\] _3132_ _3396_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__a21o_1
X_6211_ _2638_ _2644_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6142_ _2311_ _2577_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ sound3.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__inv_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _0698_ _0546_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nor2_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6975_ _3240_ _3241_ _3233_ _3237_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5926_ _2335_ _2361_ _2328_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5857_ _2277_ _2292_ _2293_ sound1.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5788_ wave_comb.u1.A\[5\] _2224_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__or2_1
X_4808_ _1242_ _1321_ _1327_ _1101_ _1358_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__o221a_1
X_7527_ sound3.sdiv.Q\[16\] _3654_ _3643_ sound3.sdiv.Q\[15\] _3395_ vssd1 vssd1 vccd1
+ vccd1 _0355_ sky130_fd_sc_hd__a221o_1
X_4739_ sound1.count\[13\] sound1.count\[14\] _1290_ vssd1 vssd1 vccd1 vccd1 _1296_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_43_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7458_ sound3.sdiv.A\[20\] _3595_ _3607_ vssd1 vssd1 vccd1 vccd1 _3613_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6409_ _2826_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__inv_2
X_7389_ sound3.divisor_m\[13\] _3543_ vssd1 vssd1 vccd1 vccd1 _3552_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6760_ sound1.sdiv.C\[2\] sound1.sdiv.C\[1\] sound1.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3106_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3972_ _0617_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__inv_2
X_5711_ _0575_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__buf_4
X_6691_ _3045_ _3047_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5642_ sound4.divisor_m\[0\] sound4.sdiv.Q\[27\] _2123_ _2124_ vssd1 vssd1 vccd1
+ vccd1 _2125_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8361_ net145 wave.next_state\[0\] net106 vssd1 vssd1 vccd1 vccd1 wave.mode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5573_ sound4.divisor_m\[14\] _2055_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7312_ sound3.divisor_m\[5\] sound3.divisor_m\[4\] _3465_ vssd1 vssd1 vccd1 vccd1
+ _3483_ sky130_fd_sc_hd__or3_1
X_4524_ _0685_ _0677_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nand2_4
XFILLER_0_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8292_ net121 _0392_ net82 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7243_ _1681_ vssd1 vssd1 vccd1 vccd1 _3427_ sky130_fd_sc_hd__inv_2
X_4455_ _0695_ _0677_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__nand2_4
X_7174_ sound3.count\[1\] _2863_ vssd1 vssd1 vccd1 vccd1 _3388_ sky130_fd_sc_hd__and2_1
X_4386_ _0909_ _0956_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6125_ _2534_ _2535_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__nor2_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _2465_ _2466_ _2462_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__a21o_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _1539_ _1540_ _1504_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__and3b_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6958_ _3215_ _3219_ _3226_ vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5909_ _2315_ sound4.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__or2_1
X_6889_ sound2.divisor_m\[0\] sound2.sdiv.Q\[27\] vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4240_ _0813_ _0826_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__and3_1
X_4171_ seq.player_1.state\[1\] seq.player_1.state\[2\] seq.player_1.state\[3\] _0770_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__a311o_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7930_ net128 _0093_ net89 vssd1 vssd1 vccd1 vccd1 sound1.divisor_m\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ net111 seq.clk_div.next_count\[18\] net72 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6812_ sound2.count_m\[5\] _2857_ _3120_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__a21o_1
X_7792_ net144 net17 net105 vssd1 vssd1 vccd1 vccd1 inputcont.u1.ff_intermediate\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_6743_ sound1.sdiv.A\[24\] _3055_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__nand2_1
X_3955_ _0611_ _0618_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6674_ _3031_ _3032_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3886_ sound4.sdiv.C\[4\] sound4.sdiv.C\[3\] sound4.sdiv.C\[2\] _0555_ sound4.sdiv.C\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5625_ _2104_ _2106_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5556_ sound4.sdiv.A\[25\] _2038_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__nand2_1
X_8344_ net121 sound4.osc.next_count\[2\] net82 vssd1 vssd1 vccd1 vccd1 sound4.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4507_ _0695_ _0680_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nand2_2
X_5487_ sound4.count\[13\] sound4.count\[14\] _1977_ vssd1 vssd1 vccd1 vccd1 _1984_
+ sky130_fd_sc_hd__and3_2
X_8275_ net120 _0375_ net81 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7226_ sound3.divisor_m\[5\] _3416_ _3142_ vssd1 vssd1 vccd1 vccd1 _3417_ sky130_fd_sc_hd__mux2_1
X_4438_ sound1.count\[1\] _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ _0699_ net35 _0917_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__a21bo_2
X_7157_ sound2.sdiv.Q\[13\] _3167_ _3349_ sound2.sdiv.Q\[12\] _3120_ vssd1 vssd1 vccd1
+ vccd1 _0253_ sky130_fd_sc_hd__a221o_1
X_6108_ sound3.count_m\[17\] _2543_ sound3.count_m\[18\] vssd1 vssd1 vccd1 vccd1 _2544_
+ sky130_fd_sc_hd__a21o_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _1311_ _3343_ vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__nand2_1
X_6039_ sound2.count_m\[2\] vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6390_ _2813_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5410_ _1101_ _1786_ _1790_ _1240_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5341_ _1830_ _1831_ _1841_ _1851_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8060_ net116 _0202_ net77 vssd1 vssd1 vccd1 vccd1 sound2.divisor_m\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7011_ sound2.divisor_m\[12\] sound2.divisor_m\[11\] _3256_ vssd1 vssd1 vccd1 vccd1
+ _3274_ sky130_fd_sc_hd__or3_1
X_5272_ _1782_ _1770_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__or2_1
X_4223_ seq.clk_div.count\[1\] seq.clk_div.count\[0\] seq.clk_div.count\[2\] seq.clk_div.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4154_ _0758_ _0757_ _0759_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_3.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4085_ seq.player_8.state\[0\] _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7913_ net127 _0076_ net88 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7844_ net108 seq.clk_div.next_count\[1\] net69 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_7775_ net139 _0049_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6726_ _3076_ _3077_ _3078_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4987_ sound2.count\[10\] sound2.count\[11\] _1524_ vssd1 vssd1 vccd1 vccd1 _1527_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3938_ _0599_ _0602_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nor2_1
X_6657_ _3005_ _3008_ _3016_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3869_ _0520_ _0541_ _0512_ _0532_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__a211oi_1
X_6588_ _2954_ _2955_ sound1.sdiv.A\[7\] _2895_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__a2bb2o_1
X_5608_ sound4.divisor_m\[7\] _2090_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__xnor2_1
X_5539_ _0657_ pm.current_waveform\[7\] _2008_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_
+ sky130_fd_sc_hd__o22a_1
X_8327_ net138 _0427_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8258_ net132 _0358_ net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[19\] sky130_fd_sc_hd__dfrtp_1
X_8189_ net142 _0310_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[4\] sky130_fd_sc_hd__dfrtp_1
X_7209_ sound3.count\[18\] _2863_ vssd1 vssd1 vccd1 vccd1 _3406_ sky130_fd_sc_hd__and2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 piano_keys[8] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4910_ sound2.count\[18\] _1445_ _1448_ _1455_ _1460_ vssd1 vssd1 vccd1 vccd1 _1461_
+ sky130_fd_sc_hd__a2111o_1
X_5890_ sound4.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _1176_ _1323_ _1338_ _1028_ _1391_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4772_ _0504_ _1320_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__nand2_8
X_7560_ _1931_ vssd1 vssd1 vccd1 vccd1 _3656_ sky130_fd_sc_hd__inv_2
X_7491_ _3640_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6511_ sound1.divisor_m\[17\] _1225_ _2864_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6442_ sound1.count_m\[8\] _2836_ _2846_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6373_ wave_comb.u1.Q\[9\] wave_comb.u1.Q\[10\] _0571_ vssd1 vssd1 vccd1 vccd1 _2801_
+ sky130_fd_sc_hd__mux2_1
X_8112_ net110 sound2.osc.next_count\[13\] net71 vssd1 vssd1 vccd1 vccd1 sound2.count\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5324_ _1004_ _1784_ _1786_ _1189_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8043_ net117 _0185_ net78 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[16\] sky130_fd_sc_hd__dfrtp_1
X_5255_ _0699_ net47 vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__and2_1
X_4206_ _0782_ _0798_ _0799_ seq.clk_div.count\[21\] seq.clk_div.count\[20\] vssd1
+ vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5186_ sound3.count\[3\] _1641_ _1681_ sound3.count\[12\] vssd1 vssd1 vccd1 vccd1
+ _1717_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ seq.player_4.state\[0\] seq.player_4.state\[1\] _0745_ vssd1 vssd1 vccd1 vccd1
+ _0748_ sky130_fd_sc_hd__and3_1
X_4068_ _0703_ _0705_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__nor2_2
XFILLER_0_66_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7827_ net113 seq.player_2.next_state\[1\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7758_ net139 _0043_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6709_ _3050_ _3058_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__or2_1
X_7689_ _3681_ _3740_ _3741_ _2184_ sound4.sdiv.A\[25\] vssd1 vssd1 vccd1 vccd1 _0430_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ net43 _1548_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__or2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6991_ sound2.divisor_m\[10\] _3245_ vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__or2_1
X_5942_ sound1.divisor_m\[11\] vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__inv_2
X_5873_ wave_comb.u1.Q\[1\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7612_ _2116_ _2127_ vssd1 vssd1 vccd1 vccd1 _3687_ sky130_fd_sc_hd__or2_1
X_4824_ _1053_ _1341_ _1345_ _1063_ _1374_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__o221a_1
X_4755_ sound1.count\[18\] _1305_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__or2_1
X_7543_ sound4.count_m\[4\] _3403_ _2191_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7474_ _3607_ _3618_ _3625_ _3626_ vssd1 vssd1 vccd1 vccd1 _3627_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4686_ sound1.count\[0\] _1256_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[0\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6425_ sound1.count_m\[0\] _2836_ _2837_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6356_ _2784_ _2745_ _2785_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__a21o_1
X_5307_ sound4.count\[14\] _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__xnor2_1
X_8026_ net128 _0168_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[27\] sky130_fd_sc_hd__dfrtp_1
X_6287_ sound2.sdiv.Q\[5\] _2660_ _2686_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5238_ sound3.count\[15\] _1750_ _1721_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__o21ai_1
X_5169_ _1154_ _1550_ _1570_ _1077_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4540_ _0685_ _0970_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nand2_4
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4471_ _0944_ _0947_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7190_ sound3.count\[9\] _2863_ vssd1 vssd1 vccd1 vccd1 _3396_ sky130_fd_sc_hd__and2_1
X_6210_ _2639_ _2279_ _2292_ _2643_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6141_ _2575_ _2576_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__xnor2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ sound3.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__inv_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _0977_ _0996_ _1550_ _1553_ _1096_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o32a_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6974_ sound2.sdiv.A\[8\] _3239_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _2336_ _2337_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5856_ sound1.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4807_ _1110_ _1336_ _1345_ _1238_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__o221a_1
X_5787_ wave_comb.u1.next_dived _2235_ _2236_ _0573_ wave_comb.u1.A\[5\] vssd1 vssd1
+ vccd1 vccd1 _0033_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7526_ sound3.sdiv.Q\[15\] _3654_ _3643_ sound3.sdiv.Q\[14\] _3394_ vssd1 vssd1 vccd1
+ vccd1 _0354_ sky130_fd_sc_hd__a221o_1
X_4738_ _1295_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7457_ sound3.sdiv.A\[21\] _3595_ vssd1 vssd1 vccd1 vccd1 _3612_ sky130_fd_sc_hd__xnor2_1
X_4669_ _0683_ _0959_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6408_ _2755_ _2790_ _2805_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7388_ sound3.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _3551_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6339_ _2767_ _2768_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__xnor2_1
X_8009_ net128 _0151_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3971_ inputcont.INTERNAL_SYNCED_I\[4\] _0512_ _0615_ _0502_ vssd1 vssd1 vccd1 vccd1
+ _0634_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_128_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5710_ _1764_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__clkbuf_8
X_6690_ sound1.divisor_m\[18\] _3046_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5641_ _2122_ sound4.sdiv.A\[0\] vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8360_ net136 sound4.osc.next_count\[18\] net97 vssd1 vssd1 vccd1 vccd1 sound4.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5572_ sound4.sdiv.A\[26\] _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7311_ sound3.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _3482_ sky130_fd_sc_hd__inv_2
X_4523_ _0996_ _1090_ _1091_ _1092_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o2111a_1
X_8291_ net123 _0391_ net84 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7242_ _3426_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4454_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__buf_8
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7173_ sound3.count_m\[0\] _3132_ _3387_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__a21o_1
X_4385_ _0940_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6124_ _2559_ _2515_ _2548_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__a21o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _2447_ _2490_ _2454_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__a21o_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ sound2.count\[15\] sound2.count\[16\] _1533_ sound2.count\[17\] vssd1 vssd1
+ vccd1 vccd1 _1540_ sky130_fd_sc_hd__a31o_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _3224_ _3225_ vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6888_ _1311_ vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__buf_6
XFILLER_0_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5908_ _2325_ _2328_ _2339_ _2343_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5839_ sound1.sdiv.Q\[0\] _0579_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7509_ _3634_ _3639_ _3652_ _0563_ _2005_ vssd1 vssd1 vccd1 vccd1 _3653_ sky130_fd_sc_hd__a311o_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4170_ seq.player_1.state\[0\] _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7860_ net107 seq.clk_div.next_count\[17\] net68 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_6811_ sound2.count\[5\] _2855_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7791_ net118 inputcont.u1.ff_intermediate\[13\] net79 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_OCTAVE_INPUT
+ sky130_fd_sc_hd__dfrtp_1
X_6742_ sound1.sdiv.A\[24\] _3055_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__or2_1
X_3954_ inputcont.INTERNAL_SYNCED_I\[11\] _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6673_ _3027_ _3030_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3885_ sound4.sdiv.start vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5624_ _2104_ _2106_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8343_ net121 sound4.osc.next_count\[1\] net82 vssd1 vssd1 vccd1 vccd1 sound4.count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_5555_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4506_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5486_ _1983_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
X_8274_ net122 _0374_ net83 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[7\] sky130_fd_sc_hd__dfrtp_1
X_7225_ _1635_ vssd1 vssd1 vccd1 vccd1 _3416_ sky130_fd_sc_hd__inv_2
X_4437_ _0962_ _0987_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nand3_1
X_7156_ sound2.sdiv.Q\[12\] _3167_ _3349_ sound2.sdiv.Q\[11\] _3119_ vssd1 vssd1 vccd1
+ vccd1 _0252_ sky130_fd_sc_hd__a221o_1
X_6107_ sound3.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4368_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__clkbuf_8
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _3339_ _3341_ _3337_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__a21o_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nor3_1
X_6038_ sound2.count_m\[3\] vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7989_ net125 sound1.osc.next_count\[10\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5340_ sound4.count\[3\] _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5271_ _1766_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__inv_2
X_7010_ sound2.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__inv_2
X_4222_ seq.clk_div.count\[2\] seq.clk_div.count\[3\] _0777_ vssd1 vssd1 vccd1 vccd1
+ _0815_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4153_ seq.player_3.state\[2\] _0756_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4084_ seq.encode.keys_edge_det\[9\] inputcont.INTERNAL_SYNCED_I\[7\] vssd1 vssd1
+ vccd1 vccd1 _0712_ sky130_fd_sc_hd__and2b_1
X_7912_ net127 _0075_ net88 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7843_ net107 seq.clk_div.next_count\[0\] net68 vssd1 vssd1 vccd1 vccd1 seq.clk_div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7774_ net139 _0048_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4986_ sound2.count\[10\] _1524_ _1526_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[10\]
+ sky130_fd_sc_hd__a21oi_1
X_6725_ sound1.sdiv.A\[21\] _3055_ vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__xnor2_1
X_3937_ _0600_ _0590_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6656_ _3005_ _3008_ _3016_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__nand3_1
X_3868_ _0521_ _0523_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6587_ _2946_ _2953_ _0866_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3799_ inputcont.INTERNAL_SYNCED_I\[4\] _0443_ inputcont.INTERNAL_SYNCED_I\[5\] vssd1
+ vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__o21ai_4
X_5607_ _2036_ _2028_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__and2_1
X_5538_ _2007_ pm.current_waveform\[6\] _2010_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8326_ net138 _0426_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[21\] sky130_fd_sc_hd__dfrtp_2
X_8257_ net132 _0357_ net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7208_ sound3.count_m\[17\] _3403_ _3405_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__a21o_1
X_5469_ sound4.count\[10\] _1966_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__nand2_1
X_8188_ net142 _0309_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7139_ _3383_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 piano_keys[9] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4840_ _1180_ _1327_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6510_ _2887_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _0499_ _1316_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__nand2_4
X_7490_ _1545_ _0577_ sound3.sdiv.C\[0\] vssd1 vssd1 vccd1 vccd1 _3640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6441_ sound1.count\[8\] _2201_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6372_ _0645_ _2798_ _2799_ _2800_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8111_ net110 sound2.osc.next_count\[12\] net71 vssd1 vssd1 vccd1 vccd1 sound2.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_5323_ net47 _1129_ _1770_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8042_ net116 _0184_ net77 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[15\] sky130_fd_sc_hd__dfrtp_1
X_5254_ _0698_ _0606_ net49 vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__or3_4
X_5185_ _1642_ _1649_ _1714_ sound3.count\[9\] _1715_ vssd1 vssd1 vccd1 vccd1 _1716_
+ sky130_fd_sc_hd__o221ai_1
X_4205_ seq.clk_div.count\[11\] seq.clk_div.count\[19\] vssd1 vssd1 vccd1 vccd1 _0799_
+ sky130_fd_sc_hd__nand2_1
X_4136_ seq.player_4.state\[0\] _0745_ _0747_ vssd1 vssd1 vccd1 vccd1 seq.player_4.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
X_4067_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__or3b_4
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7826_ net113 seq.player_2.next_state\[0\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_2.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7757_ net143 _0042_ net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4969_ sound2.count\[4\] sound2.count\[5\] _1511_ vssd1 vssd1 vccd1 vccd1 _1515_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6708_ _3050_ _3061_ _3058_ _3062_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__o31a_1
XFILLER_0_74_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7688_ _2173_ _2174_ _3739_ vssd1 vssd1 vccd1 vccd1 _3741_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6639_ sound1.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8309_ net123 _0409_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[4\] sky130_fd_sc_hd__dfrtp_1
Xfanout140 net145 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6990_ sound2.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ sound1.count_m\[14\] _2375_ sound1.count_m\[13\] _2376_ vssd1 vssd1 vccd1
+ vccd1 _2377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5872_ wave_comb.u1.Q\[0\] _2308_ _0645_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7611_ _3681_ _3685_ _3686_ _2184_ sound4.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _0407_
+ sky130_fd_sc_hd__a32o_1
X_4823_ _1057_ _1343_ _1333_ _1056_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4754_ _1307_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_7542_ sound4.count_m\[3\] _3403_ _2190_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7473_ sound3.sdiv.A\[22\] sound3.sdiv.A\[21\] sound3.sdiv.A\[20\] sound3.sdiv.A\[19\]
+ _3595_ vssd1 vssd1 vccd1 vccd1 _3626_ sky130_fd_sc_hd__o41a_1
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4685_ _1173_ _1255_ _1070_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__o21a_4
XFILLER_0_43_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6424_ sound1.count\[0\] _2201_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6355_ _2740_ _2742_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6286_ sound2.sdiv.Q\[7\] _0578_ _2286_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__and3_1
X_5306_ _1062_ _1777_ _1813_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__o211a_2
X_5237_ sound3.count\[15\] _1750_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__and2_1
X_8025_ net127 _0167_ net88 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[26\] sky130_fd_sc_hd__dfrtp_1
X_5168_ _1043_ _1559_ _1580_ _1033_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__o221a_2
XFILLER_0_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5099_ _1180_ _1553_ _1565_ _1174_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__o22a_1
X_4119_ seq.player_6.state\[1\] seq.player_6.state\[2\] _0730_ seq.player_6.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ net107 seq.player_7.next_state\[3\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_7.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _1019_ net63 vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__nor2_8
XFILLER_0_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6140_ _2291_ _2305_ _2303_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _2505_ _2506_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ net43 _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__nand2_8
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6973_ sound2.sdiv.A\[8\] _3239_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5924_ _2347_ _2359_ _2317_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__a21o_1
X_5855_ net30 net31 vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__nand2_8
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4806_ _1004_ _1133_ _1339_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5786_ _2228_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7525_ sound3.sdiv.Q\[14\] _3654_ _3643_ sound3.sdiv.Q\[13\] _3393_ vssd1 vssd1 vccd1
+ vccd1 _0353_ sky130_fd_sc_hd__a221o_1
X_4737_ _1256_ _1293_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7456_ sound3.sdiv.A\[21\] _3463_ sound3.sdiv.next_dived _3611_ vssd1 vssd1 vccd1
+ vccd1 _0327_ sky130_fd_sc_hd__a22o_1
X_4668_ _1004_ _1003_ _1028_ _1238_ _1000_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__o32a_1
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6407_ _2825_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
X_7387_ _3437_ _3549_ _3550_ _3440_ sound3.sdiv.A\[13\] vssd1 vssd1 vccd1 vccd1 _0319_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4599_ _1070_ _1161_ _1163_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__and4_2
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6338_ sound3.sdiv.Q\[7\] _0577_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6269_ sound3.sdiv.Q\[5\] _0577_ _2699_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__a21o_1
X_8008_ net128 _0150_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ inputcont.INTERNAL_SYNCED_I\[10\] _0610_ _0608_ vssd1 vssd1 vccd1 vccd1 _0633_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5640_ sound4.sdiv.A\[0\] _2122_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5571_ sound4.divisor_m\[13\] _2032_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nor2_1
X_7310_ _3437_ _3480_ _3481_ _3440_ sound3.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _0311_
+ sky130_fd_sc_hd__a32o_1
X_4522_ _0992_ _1003_ _0948_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__a21o_1
X_8290_ net121 _0390_ net82 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7241_ sound3.divisor_m\[11\] _3425_ _3419_ vssd1 vssd1 vccd1 vccd1 _3426_ sky130_fd_sc_hd__mux2_1
X_4453_ _0685_ _0681_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7172_ sound3.count\[0\] _2855_ vssd1 vssd1 vccd1 vccd1 _3387_ sky130_fd_sc_hd__and2_1
X_4384_ _0926_ _0936_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__nor2b_2
X_6123_ _2558_ _2512_ _2549_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__a21o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _2449_ _2489_ _2442_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__a21o_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ sound2.count\[16\] sound2.count\[17\] _1536_ vssd1 vssd1 vccd1 vccd1 _1539_
+ sky130_fd_sc_hd__and3_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _3220_ _3223_ vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5907_ _2340_ sound4.divisor_m\[16\] sound4.divisor_m\[9\] _2334_ _2342_ vssd1 vssd1
+ vccd1 vccd1 _2343_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6887_ _2843_ _1445_ _3163_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5838_ sound2.sdiv.Q\[0\] _0578_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5769_ _2219_ _2215_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7508_ sound3.divisor_m\[18\] sound3.divisor_m\[17\] sound3.sdiv.A\[26\] _3578_ vssd1
+ vssd1 vccd1 vccd1 _3652_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7439_ _3590_ _3592_ _3589_ vssd1 vssd1 vccd1 vccd1 _3597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6810_ sound2.count_m\[4\] _2857_ _3119_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7790_ net122 inputcont.u1.ff_intermediate\[12\] net83 vssd1 vssd1 vccd1 vccd1 inputcont.INTERNAL_SYNCED_I\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_6741_ sound1.sdiv.A\[23\] _3055_ _3089_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3953_ _0615_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6672_ _3027_ _3030_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__or2_1
X_3884_ rate_clk.count\[7\] _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__nand2_8
XFILLER_0_42_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5623_ sound4.divisor_m\[4\] _2105_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8342_ net121 sound4.osc.next_count\[0\] net82 vssd1 vssd1 vccd1 vccd1 sound4.count\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5554_ sound4.divisor_m\[18\] _2035_ _2036_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4505_ _0679_ _1046_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__or2_1
X_5485_ _1779_ _1936_ _1981_ _1982_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__and4_1
X_8273_ net122 _0373_ net83 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7224_ _3415_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
X_4436_ _0990_ _0978_ _0944_ _0998_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__o311a_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4367_ _0909_ _0918_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__or3_1
X_7155_ sound2.sdiv.Q\[11\] _3167_ _3349_ sound2.sdiv.Q\[10\] _3118_ vssd1 vssd1 vccd1
+ vccd1 _0251_ sky130_fd_sc_hd__a221o_1
X_6106_ net59 vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _3337_ _3339_ _3341_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__and3_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__buf_6
X_6037_ _2472_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__inv_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ net125 sound1.osc.next_count\[9\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6939_ _3197_ _3200_ _3208_ vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__or3b_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _1780_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4221_ seq.clk_div.count\[2\] _0777_ _0814_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[2\]
+ sky130_fd_sc_hd__a21oi_1
X_4152_ seq.player_3.state\[2\] seq.player_3.state\[3\] vssd1 vssd1 vccd1 vccd1 _0758_
+ sky130_fd_sc_hd__nand2_1
X_4083_ _0711_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7911_ net126 _0074_ net87 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[4\] sky130_fd_sc_hd__dfrtp_1
X_7842_ net143 _0065_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7773_ net143 _0047_ net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4985_ sound2.count\[10\] _1524_ _1504_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__o21ai_1
X_6724_ sound1.sdiv.A\[20\] sound1.sdiv.A\[19\] _3055_ vssd1 vssd1 vccd1 vccd1 _3077_
+ sky130_fd_sc_hd__o21ai_1
X_3936_ _0473_ _0486_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6655_ _3014_ _3015_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__nand2_1
X_3867_ _0540_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__inv_2
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6586_ _2946_ _2953_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3798_ inputcont.INTERNAL_SYNCED_I\[10\] _0445_ _0474_ _0475_ _0476_ vssd1 vssd1
+ vccd1 vccd1 _0477_ sky130_fd_sc_hd__a2111o_1
X_5606_ _2087_ _2088_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nand2_1
X_5537_ _2009_ pm.current_waveform\[5\] _2011_ _2020_ vssd1 vssd1 vccd1 vccd1 _2021_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8325_ net124 _0425_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8256_ net131 _0356_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7207_ sound3.count\[17\] _2863_ vssd1 vssd1 vccd1 vccd1 _3405_ sky130_fd_sc_hd__and2_1
X_5468_ _1969_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_8187_ net142 _0308_ net103 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[2\] sky130_fd_sc_hd__dfrtp_1
X_4419_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5399_ sound4.count\[2\] _1903_ _1909_ sound4.count\[11\] vssd1 vssd1 vccd1 vccd1
+ _1910_ sky130_fd_sc_hd__a2bb2o_1
X_7138_ _2843_ _3382_ vssd1 vssd1 vccd1 vccd1 _3383_ sky130_fd_sc_hd__and2_1
X_7069_ sound2.sdiv.A\[18\] _3168_ sound2.sdiv.next_dived _3326_ vssd1 vssd1 vccd1
+ vccd1 _0225_ sky130_fd_sc_hd__a22o_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 seq_play vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ net40 _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nand2_4
XFILLER_0_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6440_ sound1.count_m\[7\] _2836_ _2845_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6371_ wave_comb.u1.Q\[9\] _0573_ _0646_ wave_comb.u1.Q\[8\] vssd1 vssd1 vccd1 vccd1
+ _2800_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8110_ net110 sound2.osc.next_count\[11\] net71 vssd1 vssd1 vccd1 vccd1 sound2.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_5322_ _0677_ _1832_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8041_ net109 _0183_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[14\] sky130_fd_sc_hd__dfrtp_1
X_5253_ _1764_ vssd1 vssd1 vccd1 vccd1 sound4.sdiv.next_dived sky130_fd_sc_hd__buf_4
X_5184_ sound3.count\[9\] _1714_ _1699_ sound3.count\[11\] vssd1 vssd1 vccd1 vccd1
+ _1715_ sky130_fd_sc_hd__o2bb2a_1
X_4204_ seq.clk_div.count\[3\] seq.clk_div.count\[17\] _0785_ seq.clk_div.count\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__or4bb_1
X_4135_ seq.player_4.state\[1\] seq.player_4.state\[2\] seq.player_4.state\[3\] _0746_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__a311o_1
X_4066_ _0703_ _0704_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__nor2_1
Xwire54 _2797_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7825_ net113 seq.player_3.next_state\[3\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_3.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7756_ net143 _0041_ net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4968_ sound2.count\[4\] _1511_ _1514_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6707_ _3048_ _3056_ _3057_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7687_ _2173_ _2174_ _3739_ vssd1 vssd1 vccd1 vccd1 _3740_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4899_ _0499_ _1315_ _1319_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__a21oi_1
X_3919_ _0529_ _0525_ _0549_ _0582_ _0526_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__a41o_1
XFILLER_0_104_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6638_ _2890_ _2999_ _3000_ _2894_ sound1.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _0120_
+ sky130_fd_sc_hd__a32o_1
X_6569_ _2903_ _2937_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__and2_1
X_8308_ net123 _0408_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[3\] sky130_fd_sc_hd__dfrtp_1
X_8239_ net143 _0339_ net104 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[0\] sky130_fd_sc_hd__dfrtp_1
Xfanout130 net134 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_8
Xfanout141 net145 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5940_ sound1.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5871_ _2306_ _2307_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__xnor2_1
X_7610_ _2120_ _2125_ vssd1 vssd1 vccd1 vccd1 _3686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4822_ _1064_ _1347_ _1322_ _0979_ _1317_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__o221a_1
X_4753_ _1305_ _1306_ _1256_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7541_ sound4.count_m\[2\] _3403_ _2189_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7472_ _3624_ _3612_ vssd1 vssd1 vccd1 vccd1 _3625_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6423_ _0554_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__buf_4
X_4684_ _1187_ _1197_ _1209_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6354_ _2742_ _2740_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__or2b_1
X_6285_ wave_comb.u1.next_start _2714_ _2715_ _2716_ vssd1 vssd1 vccd1 vccd1 _0051_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5305_ _1814_ _1815_ _0695_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a21o_1
X_5236_ _1752_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_8024_ net127 _0166_ net88 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5167_ _1004_ _1693_ _1694_ _1001_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__o221a_1
X_5098_ sound3.count\[14\] _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__xor2_1
X_4118_ _0734_ _0733_ _0735_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_6.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_4049_ _0682_ _0683_ _0687_ _0689_ _0681_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o32a_1
XFILLER_0_79_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7808_ net108 seq.player_7.next_state\[2\] net69 vssd1 vssd1 vccd1 vccd1 seq.player_7.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7739_ net137 _0024_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _2281_ _2299_ _2297_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__a21o_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ net56 _1551_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__nor2_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6972_ sound2.divisor_m\[9\] _3238_ vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5923_ _2314_ _2358_ _2319_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5854_ _2181_ _2289_ _2290_ sound4.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4805_ _1025_ _1323_ _1338_ _1240_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__o221a_1
X_7524_ sound3.sdiv.Q\[13\] _3654_ _3643_ sound3.sdiv.Q\[12\] _3392_ vssd1 vssd1 vccd1
+ vccd1 _0352_ sky130_fd_sc_hd__a221o_1
X_5785_ _2228_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4736_ sound1.count\[13\] _1290_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__or2_1
X_7455_ _3609_ _3610_ vssd1 vssd1 vccd1 vccd1 _3611_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4667_ _0681_ _0944_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7386_ _3537_ _3541_ _3548_ vssd1 vssd1 vccd1 vccd1 _3550_ sky130_fd_sc_hd__nand3_1
X_6406_ pm.current_waveform\[7\] _2824_ _2808_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6337_ sound3.sdiv.Q\[6\] _2632_ _2731_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__a21o_1
X_4598_ _1003_ _1164_ _1165_ _0943_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__o221a_1
X_6268_ sound3.sdiv.Q\[5\] _2699_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6199_ sound3.sdiv.Q\[2\] _2632_ _2602_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__a21o_1
X_5219_ sound3.count\[9\] _1738_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__and2_1
X_8007_ net128 _0149_ net89 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5570_ _2050_ _2052_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__nor2_1
X_4521_ _0993_ _0943_ _1012_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7240_ _1699_ vssd1 vssd1 vccd1 vccd1 _3425_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4452_ _1011_ _0967_ _1003_ _1014_ _1022_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4383_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7171_ sound2.sdiv.Q\[27\] _3168_ _3164_ sound2.sdiv.Q\[26\] vssd1 vssd1 vccd1 vccd1
+ _0267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6122_ _2553_ _2557_ _2510_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _2452_ _2488_ _2451_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__a21bo_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ sound2.count\[16\] _1536_ _1538_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[16\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6955_ _3220_ _3223_ vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ sound4.count_m\[15\] _2341_ sound4.count_m\[14\] _2331_ vssd1 vssd1 vccd1
+ vccd1 _2342_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6886_ _2470_ _2005_ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5837_ sound3.sdiv.Q\[0\] _0577_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5768_ wave_comb.u1.A\[2\] _0573_ wave_comb.u1.next_dived _2220_ vssd1 vssd1 vccd1
+ vccd1 _0030_ sky130_fd_sc_hd__a22o_1
X_7507_ _3651_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__clkbuf_1
X_4719_ sound1.count\[9\] _1278_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__and2_1
X_7438_ sound3.sdiv.A\[18\] _3595_ vssd1 vssd1 vccd1 vccd1 _3596_ sky130_fd_sc_hd__xnor2_1
X_5699_ _1763_ _2180_ _2181_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7369_ sound3.sdiv.A\[11\] vssd1 vssd1 vccd1 vccd1 _3534_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ sound1.sdiv.A\[24\] _2895_ _3088_ _3090_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3952_ _0612_ _0614_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__and2_1
X_6671_ sound1.divisor_m\[16\] _3029_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__xnor2_1
X_3883_ rate_clk.count\[6\] _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__and2_2
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5622_ _2036_ _2026_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8341_ net138 sound4.sdiv.next_start net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.start
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5553_ sound4.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4504_ _0688_ _0958_ _0943_ _0971_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5484_ sound4.count\[13\] _1977_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8272_ net123 _0372_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[5\] sky130_fd_sc_hd__dfrtp_1
X_7223_ sound3.divisor_m\[4\] _3414_ _3142_ vssd1 vssd1 vccd1 vccd1 _3415_ sky130_fd_sc_hd__mux2_1
X_4435_ _1000_ _1001_ _1003_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4366_ _0926_ _0936_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7154_ sound2.sdiv.Q\[10\] _3167_ _3349_ sound2.sdiv.Q\[9\] _3117_ vssd1 vssd1 vccd1
+ vccd1 _0250_ sky130_fd_sc_hd__a221o_1
X_6105_ _2523_ _2526_ _2537_ _2540_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _3321_ _3330_ _3331_ _3340_ vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__o211a_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _0674_ _0677_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__or2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ sound2.count_m\[17\] _2470_ sound2.count_m\[16\] _2471_ vssd1 vssd1 vccd1
+ vccd1 _2472_ sky130_fd_sc_hd__o22a_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ net125 sound1.osc.next_count\[8\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _3197_ _3200_ _3208_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__o21bai_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6869_ _1488_ vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4220_ seq.clk_div.count\[2\] _0777_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ seq.player_3.state\[2\] seq.player_3.state\[3\] _0756_ _0757_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_3.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_4082_ net1 pm.pwm_o vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7910_ net128 _0073_ net89 vssd1 vssd1 vccd1 vccd1 sound1.count_m\[3\] sky130_fd_sc_hd__dfrtp_1
X_7841_ net143 _0064_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7772_ net139 _0046_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[1\] sky130_fd_sc_hd__dfrtp_1
X_4984_ _1524_ _1525_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[9\] sky130_fd_sc_hd__nor2_1
X_6723_ sound1.sdiv.A\[20\] _3055_ _3069_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3935_ _0547_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6654_ _3010_ _3013_ vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3866_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5605_ sound4.sdiv.A\[7\] _2086_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6585_ _2951_ _2952_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3797_ inputcont.INTERNAL_SYNCED_I\[6\] _0443_ _0463_ inputcont.INTERNAL_SYNCED_I\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__o31a_1
X_5536_ _0651_ pm.current_waveform\[4\] _2013_ _2019_ vssd1 vssd1 vccd1 vccd1 _2020_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8324_ net124 _0424_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[19\] sky130_fd_sc_hd__dfrtp_4
X_8255_ net131 _0355_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[16\] sky130_fd_sc_hd__dfrtp_1
X_5467_ _1779_ _1936_ _1967_ _1968_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__and4_1
XFILLER_0_112_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7206_ sound3.count_m\[16\] _3403_ _3404_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a21o_1
X_4418_ _0926_ _0936_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__or3_1
X_8186_ net141 _0307_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[1\] sky130_fd_sc_hd__dfrtp_1
X_5398_ _1035_ _1769_ _1792_ _1041_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__o221a_2
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7137_ sound2.sdiv.C\[3\] _0559_ _3378_ sound2.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1
+ _3382_ sky130_fd_sc_hd__a31o_1
X_4349_ seq.player_6.state\[2\] _0894_ _0896_ _0919_ vssd1 vssd1 vccd1 vccd1 _0920_
+ sky130_fd_sc_hd__a22o_1
X_7068_ _3323_ _3325_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__xnor2_1
X_6019_ sound2.count_m\[8\] sound2.divisor_m\[9\] vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__or2b_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6370_ _2794_ net54 _2796_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5321_ _1782_ _1771_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__nor2_1
X_8040_ net109 _0182_ net70 vssd1 vssd1 vccd1 vccd1 sound2.count_m\[13\] sky130_fd_sc_hd__dfrtp_1
X_5252_ _1763_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5183_ _1709_ _1711_ _1713_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__and3_1
X_4203_ seq.clk_div.count\[20\] _0664_ _0665_ seq.clk_div.count\[21\] vssd1 vssd1
+ vccd1 vccd1 _0797_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4134_ seq.player_4.state\[0\] _0745_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4065_ seq.beat\[0\] seq.beat\[2\] seq.beat\[1\] vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__or3b_4
Xwire55 _3086_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_7824_ net113 seq.player_3.next_state\[2\] net74 vssd1 vssd1 vccd1 vccd1 seq.player_3.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7755_ net143 _0040_ net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4967_ sound2.count\[4\] _1511_ _1504_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6706_ _3031_ _3040_ _3041_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__a21bo_1
X_7686_ sound4.sdiv.A\[24\] _2038_ vssd1 vssd1 vccd1 vccd1 _3739_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4898_ _1333_ _1325_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__nand2_1
X_3918_ _0549_ _0582_ _0529_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6637_ _2987_ _2991_ _2998_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__o21bai_2
X_3849_ _0488_ _0491_ _0441_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__a211oi_4
X_6568_ sound1.divisor_m\[5\] sound1.divisor_m\[4\] _2919_ vssd1 vssd1 vccd1 vccd1
+ _2937_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8307_ net123 _0407_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5519_ _0553_ _2004_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[6\] sky130_fd_sc_hd__nor2_1
X_6499_ _2880_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8238_ net137 sound4.sdiv.next_dived net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.dived
+ sky130_fd_sc_hd__dfrtp_1
X_8169_ net140 _0290_ net101 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout131 net133 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_4
Xfanout120 net2 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_4
Xfanout142 net145 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_4
XFILLER_0_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5870_ _2181_ _2286_ _2284_ _2283_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4821_ _0944_ _1327_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4752_ sound1.count\[15\] sound1.count\[16\] _1296_ sound1.count\[17\] vssd1 vssd1
+ vccd1 vccd1 _1306_ sky130_fd_sc_hd__a31o_1
X_7540_ sound4.count_m\[1\] _3403_ _2188_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7471_ _3609_ vssd1 vssd1 vccd1 vccd1 _3624_ sky130_fd_sc_hd__inv_2
X_4683_ _1228_ _1236_ _1251_ _1253_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__or4b_1
XFILLER_0_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6422_ seq.beat\[3\] _2834_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6353_ _2779_ _2782_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6284_ wave_comb.u1.Q\[6\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5304_ _0680_ _1784_ _1792_ _0684_ _1800_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__o221a_1
X_5235_ _1750_ _1751_ _1721_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__and3b_1
X_8023_ net134 _0165_ net95 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _1041_ _1567_ _1565_ _1129_ _1696_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__o221a_1
X_5097_ _1624_ _1627_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__nand2_1
X_4117_ seq.player_6.state\[2\] _0732_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__xor2_1
X_4048_ _0691_ vssd1 vssd1 vccd1 vccd1 oct.next_state\[0\] sky130_fd_sc_hd__clkbuf_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ sound1.sdiv.Q\[1\] vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7807_ net107 seq.player_7.next_state\[1\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_7.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_7738_ net122 _0023_ net83 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7669_ _2168_ _2041_ vssd1 vssd1 vccd1 vccd1 _3727_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _0698_ _0546_ net46 vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__or3_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6971_ _2460_ _3230_ sound2.sdiv.A\[26\] vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5922_ _2313_ sound4.divisor_m\[4\] _2348_ _2357_ _2320_ vssd1 vssd1 vccd1 vccd1
+ _2358_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5853_ sound4.sdiv.next_start _2279_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5784_ wave_comb.u1.A\[4\] _2224_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4804_ _1004_ _1028_ _1322_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__or3_1
X_7523_ sound3.sdiv.Q\[12\] _3654_ _3643_ sound3.sdiv.Q\[11\] _3391_ vssd1 vssd1 vccd1
+ vccd1 _0351_ sky130_fd_sc_hd__a221o_1
X_4735_ sound1.count\[13\] _1290_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7454_ sound3.sdiv.A\[19\] _3595_ _3607_ vssd1 vssd1 vccd1 vccd1 _3610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ sound1.count\[6\] vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7385_ _3537_ _3541_ _3548_ vssd1 vssd1 vccd1 vccd1 _3549_ sky130_fd_sc_hd__a21o_1
X_6405_ _2725_ _2748_ _2805_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__mux2_1
X_4597_ _0990_ _0997_ _0992_ _1166_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__o221a_1
X_6336_ _2764_ _2765_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6267_ sound3.sdiv.Q\[4\] _2632_ _2669_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__a21o_1
X_6198_ sound3.sdiv.next_start _2570_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__nor2_1
X_5218_ _1740_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_8006_ net135 _0148_ net96 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[7\] sky130_fd_sc_hd__dfrtp_2
X_5149_ _1101_ _1553_ _1678_ _1679_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4520_ _0976_ _0994_ _0960_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4451_ _0979_ _0958_ _0992_ _1016_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__o221a_1
XFILLER_0_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7170_ sound2.sdiv.Q\[26\] _3167_ _1311_ sound2.sdiv.Q\[25\] _3134_ vssd1 vssd1 vccd1
+ vccd1 _0266_ sky130_fd_sc_hd__a221o_1
X_6121_ _2518_ _2520_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__nand2_1
X_4382_ _0951_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__or2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6052_ sound2.count_m\[10\] _2443_ _2455_ _2456_ _2444_ vssd1 vssd1 vccd1 vccd1 _2488_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ sound2.count\[16\] _1536_ _1504_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__o21ai_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6954_ sound2.divisor_m\[7\] _3222_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5905_ sound4.divisor_m\[16\] vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6885_ _3162_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5836_ wave_comb.u1.Q\[0\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5767_ _2215_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7506_ sound3.sdiv.C\[5\] _0554_ vssd1 vssd1 vccd1 vccd1 _3651_ sky130_fd_sc_hd__and2_1
X_4718_ _1280_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_5698_ sound4.sdiv.Q\[0\] _0576_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__and2_2
XFILLER_0_8_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7437_ _3594_ vssd1 vssd1 vccd1 vccd1 _3595_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4649_ sound1.count\[15\] _1215_ _1219_ sound1.count\[16\] vssd1 vssd1 vccd1 vccd1
+ _1220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7368_ _3532_ _3533_ sound3.sdiv.A\[11\] _3463_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7299_ _3458_ _3461_ _3470_ vssd1 vssd1 vccd1 vccd1 _3472_ sky130_fd_sc_hd__or3b_1
X_6319_ sound1.sdiv.Q\[6\] _2656_ _2722_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3951_ _0612_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6670_ _2903_ _3028_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__and2_1
X_3882_ rate_clk.count\[5\] rate_clk.count\[4\] _0551_ vssd1 vssd1 vccd1 vccd1 _0552_
+ sky130_fd_sc_hd__and3_1
X_5621_ sound4.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__inv_2
X_8340_ net145 _0440_ net106 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.M\[2\] sky130_fd_sc_hd__dfrtp_1
X_5552_ sound4.divisor_m\[17\] _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4503_ _1015_ _0981_ _0969_ _0946_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__o22a_1
X_8271_ net123 _0371_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5483_ sound4.count\[13\] _1977_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7222_ _1601_ vssd1 vssd1 vccd1 vccd1 _3414_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4434_ _0944_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__nor2_2
XFILLER_0_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4365_ _0699_ net38 _0934_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7153_ sound2.sdiv.Q\[9\] _3174_ _3349_ sound2.sdiv.Q\[8\] _3116_ vssd1 vssd1 vccd1
+ vccd1 _0249_ sky130_fd_sc_hd__a221o_1
X_6104_ _2538_ sound3.divisor_m\[16\] sound3.divisor_m\[9\] _2532_ _2539_ vssd1 vssd1
+ vccd1 vccd1 _2540_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7084_ _3323_ _3330_ _3331_ _3324_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__or4bb_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _0867_ vssd1 vssd1 vccd1 vccd1 sound1.sdiv.next_dived sky130_fd_sc_hd__buf_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ sound2.divisor_m\[17\] vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__inv_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7986_ net125 sound1.osc.next_count\[7\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _3206_ _3207_ vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__nand2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6868_ _3152_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5819_ _0646_ _0573_ wave_comb.u1.C\[0\] vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6799_ sound1.sdiv.Q\[26\] _2893_ _0867_ sound1.sdiv.Q\[25\] _2858_ vssd1 vssd1 vccd1
+ vccd1 _0167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ seq.player_3.state\[1\] _0754_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4081_ _0710_ vssd1 vssd1 vccd1 vccd1 tempo_select_on sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7840_ net143 _0063_ net104 vssd1 vssd1 vccd1 vccd1 pm.current_waveform\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7771_ net139 _0045_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.Q\[0\] sky130_fd_sc_hd__dfrtp_1
X_4983_ sound2.count\[9\] _1522_ _1504_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6722_ _3074_ _3075_ sound1.sdiv.A\[21\] _2895_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3934_ _0514_ _0533_ _0510_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6653_ _3010_ _3013_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__or2_1
X_3865_ _0534_ _0535_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5604_ sound4.sdiv.A\[7\] _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__nand2_1
X_6584_ _2947_ _2950_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3796_ inputcont.INTERNAL_SYNCED_I\[8\] _0443_ _0444_ inputcont.INTERNAL_SYNCED_I\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__o31a_2
X_5535_ _2012_ pm.current_waveform\[3\] pm.current_waveform\[2\] _2014_ _2018_ vssd1
+ vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__o221a_1
X_8323_ net123 _0423_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8254_ net131 _0354_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5466_ sound4.count\[9\] _1962_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7205_ sound3.count\[16\] _2863_ vssd1 vssd1 vccd1 vccd1 _3404_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4417_ _0909_ _0940_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__or2_2
XFILLER_0_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8185_ net140 _0306_ net101 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.A\[0\] sky130_fd_sc_hd__dfrtp_1
X_5397_ _1129_ _1777_ _1905_ _1906_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__o2111a_1
X_4348_ seq.player_7.state\[2\] _0898_ _0901_ seq.player_8.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _0919_ sky130_fd_sc_hd__a22o_1
X_7136_ _2005_ _3380_ _3381_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__nor3_1
X_7067_ _3306_ _3315_ _3324_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__a21o_1
X_4279_ _0855_ _0813_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__and3b_1
X_6018_ sound2.count_m\[15\] _2446_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__and2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ net134 _0132_ net95 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[24\] sky130_fd_sc_hd__dfrtp_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5320_ sound4.count\[8\] _1829_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__nor2_1
X_5251_ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4202_ seq.clk_div.count\[7\] vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__inv_2
X_5182_ _1189_ _1553_ _1580_ _1028_ _1712_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__o221a_1
X_4133_ _0607_ seq.encode.keys_edge_det\[5\] vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nor2_1
X_4064_ _0701_ _0703_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__nor2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7823_ net114 seq.player_3.next_state\[1\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_3.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_7754_ net143 _0039_ net104 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.C\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6705_ sound1.sdiv.A\[19\] _2895_ sound1.sdiv.next_dived _3060_ vssd1 vssd1 vccd1
+ vccd1 _0127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4966_ _1513_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7685_ _1763_ _2174_ _3737_ _3738_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__o31ai_1
X_4897_ sound2.count\[18\] _1445_ _1447_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3917_ _0510_ _0513_ _0533_ _0530_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__o31a_2
X_6636_ _2987_ _2991_ _2998_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3848_ inputcont.INTERNAL_SYNCED_I\[9\] _0454_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6567_ sound1.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3779_ inputcont.INTERNAL_SYNCED_I\[10\] _0445_ inputcont.INTERNAL_SYNCED_I\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__or3b_1
X_8306_ net138 _0406_ net99 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[1\] sky130_fd_sc_hd__dfrtp_1
X_5518_ rate_clk.count\[6\] _0552_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6498_ sound1.divisor_m\[12\] _2879_ _2864_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8237_ net135 sound3.osc.next_count\[18\] net96 vssd1 vssd1 vccd1 vccd1 sound3.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_5449_ _1954_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
X_8168_ net140 _0289_ net101 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[2\] sky130_fd_sc_hd__dfrtp_2
Xfanout121 net2 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
Xfanout110 net115 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__buf_4
Xfanout143 net144 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_4
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
X_7119_ sound2.sdiv.A\[25\] _3168_ sound2.sdiv.next_dived _3369_ vssd1 vssd1 vccd1
+ vccd1 _0232_ sky130_fd_sc_hd__a22o_1
X_8099_ net111 sound2.osc.next_count\[0\] net72 vssd1 vssd1 vccd1 vccd1 sound2.count\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4820_ _0679_ _1040_ _1321_ _1323_ _1059_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__o32a_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ sound1.count\[16\] sound1.count\[17\] _1299_ vssd1 vssd1 vccd1 vccd1 _1305_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_8_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7470_ _3621_ _3622_ vssd1 vssd1 vccd1 vccd1 _3623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4682_ _1073_ _1089_ _1104_ sound1.count\[0\] _1252_ vssd1 vssd1 vccd1 vccd1 _1253_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6421_ _2835_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6352_ _2780_ _2739_ _2781_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6283_ wave_comb.u1.Q\[5\] _0645_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5303_ _1769_ _1781_ _0687_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__a21o_1
X_5234_ sound3.count\[12\] sound3.count\[13\] _1744_ sound3.count\[14\] vssd1 vssd1
+ vccd1 vccd1 _1751_ sky130_fd_sc_hd__a31o_1
X_8022_ net125 _0164_ net86 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[23\] sky130_fd_sc_hd__dfrtp_1
X_5165_ _0947_ _1611_ _1695_ _1035_ _1562_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__o32a_1
X_4116_ seq.player_6.state\[2\] seq.player_6.state\[3\] vssd1 vssd1 vccd1 vccd1 _0734_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5096_ _1095_ _1550_ _1626_ _0695_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__o22a_1
X_4047_ _0679_ _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__or2_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ net107 seq.player_7.next_state\[0\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_7.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _2394_ _2404_ _2422_ _2433_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__a31o_2
XFILLER_0_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4949_ _1497_ _1499_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__nand2_1
X_7737_ net122 _0022_ net83 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7668_ sound4.sdiv.A\[19\] _2183_ _3681_ _3726_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6619_ sound1.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__inv_2
X_7599_ sound4.divisor_m\[17\] _0554_ vssd1 vssd1 vccd1 vccd1 _3679_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6970_ _3164_ _3236_ _3237_ _3174_ sound2.sdiv.A\[8\] vssd1 vssd1 vccd1 vccd1 _0215_
+ sky130_fd_sc_hd__a32o_1
X_5921_ _2351_ _2353_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__or2b_1
X_5852_ _2288_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__buf_4
X_5783_ _2229_ _2231_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4803_ _1245_ _1341_ _1343_ _0985_ _1353_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__o221a_1
X_7522_ sound3.sdiv.Q\[11\] _3654_ _3643_ sound3.sdiv.Q\[10\] _3390_ vssd1 vssd1 vccd1
+ vccd1 _0350_ sky130_fd_sc_hd__a221o_1
X_4734_ _1292_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7453_ sound3.sdiv.A\[20\] _3595_ vssd1 vssd1 vccd1 vccd1 _3609_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4665_ sound1.count\[14\] _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7384_ _3546_ _3547_ vssd1 vssd1 vccd1 vccd1 _3548_ sky130_fd_sc_hd__nand2_1
X_6404_ _2823_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4596_ _0994_ _1126_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6335_ _2728_ _2729_ _2726_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__o21a_1
X_6266_ _2696_ _2697_ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__xor2_1
X_8005_ net135 _0147_ net96 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[6\] sky130_fd_sc_hd__dfrtp_2
X_6197_ _2619_ _2630_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__xnor2_1
X_5217_ _1738_ _1739_ _1721_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__and3b_1
X_5148_ _1240_ _1578_ _1550_ _1242_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__o22a_1
X_5079_ _1562_ _1548_ _0869_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4450_ _0950_ _1017_ _1020_ _0994_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4381_ _0674_ _0684_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nor2_8
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6120_ _2520_ _2542_ _2550_ _2555_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__or4b_1
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _2473_ _2476_ _2477_ _2486_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__nor4_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5002_ _1536_ _1537_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[15\] sky130_fd_sc_hd__nor2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6953_ _3177_ _3221_ vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6884_ sound2.divisor_m\[17\] _1446_ _3142_ vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__mux2_1
X_5904_ sound4.count_m\[15\] vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__inv_2
X_5835_ wave_comb.u1.A\[9\] _2224_ _2261_ _2272_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5766_ _2216_ _2218_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7505_ _3650_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__clkbuf_1
X_4717_ _1278_ _1279_ _1256_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__and3b_1
X_5697_ sound4.divisor_m\[18\] sound4.sdiv.A\[26\] _2035_ _2039_ _2179_ vssd1 vssd1
+ vccd1 vccd1 _2180_ sky130_fd_sc_hd__o311a_1
XFILLER_0_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7436_ sound3.divisor_m\[18\] sound3.divisor_m\[17\] _3578_ _3448_ vssd1 vssd1 vccd1
+ vccd1 _3594_ sky130_fd_sc_hd__o31a_1
X_4648_ _0688_ _1216_ _1070_ _1217_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_114_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7367_ _3518_ _3524_ _3531_ _0563_ _2005_ vssd1 vssd1 vccd1 vccd1 _3533_ sky130_fd_sc_hd__a311o_1
X_4579_ _0680_ _0959_ _0958_ _1149_ _1070_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__o311a_1
X_7298_ _3458_ _3461_ _3470_ vssd1 vssd1 vccd1 vccd1 _3471_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6318_ wave_comb.u1.next_start _2747_ _2748_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a21o_1
X_6249_ wave_comb.u1.Q\[5\] _0572_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3950_ _0496_ _0613_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3881_ rate_clk.count\[3\] _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5620_ sound4.sdiv.A\[4\] _2102_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5551_ sound4.divisor_m\[16\] _2033_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__or2_1
X_4502_ sound1.count\[7\] vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__inv_2
X_8270_ net123 _0370_ net84 vssd1 vssd1 vccd1 vccd1 sound4.count_m\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7221_ _3413_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
X_5482_ _1980_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4433_ _0972_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__buf_8
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4364_ _0698_ seq.player_1.state\[3\] _0871_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7152_ sound2.sdiv.Q\[8\] _3174_ _3349_ sound2.sdiv.Q\[7\] _3115_ vssd1 vssd1 vccd1
+ vccd1 _0248_ sky130_fd_sc_hd__a221o_1
X_6103_ _2538_ sound3.divisor_m\[16\] sound3.count_m\[14\] _2529_ vssd1 vssd1 vccd1
+ vccd1 _2539_ sky130_fd_sc_hd__o2bb2a_1
X_4295_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__inv_4
X_7083_ _3294_ _3298_ _3323_ _3338_ _3332_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ sound2.divisor_m\[18\] vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__inv_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7985_ net134 sound1.osc.next_count\[6\] net95 vssd1 vssd1 vccd1 vccd1 sound1.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _3203_ _3205_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6867_ sound2.divisor_m\[10\] _3151_ _3142_ vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5818_ _2261_ _2262_ wave_comb.u1.A\[10\] _0573_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a2bb2o_1
X_6798_ sound1.sdiv.Q\[25\] _2893_ _0867_ sound1.sdiv.Q\[24\] _2856_ vssd1 vssd1 vccd1
+ vccd1 _0166_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5749_ sound4.count\[18\] _2201_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7419_ _3448_ _3578_ vssd1 vssd1 vccd1 vccd1 _3579_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4080_ net1 net21 vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7770_ net133 pm.next_pwm_o net94 vssd1 vssd1 vccd1 vccd1 pm.pwm_o sky130_fd_sc_hd__dfrtp_1
X_4982_ sound2.count\[8\] sound2.count\[9\] _1520_ vssd1 vssd1 vccd1 vccd1 _1524_
+ sky130_fd_sc_hd__and3_1
X_6721_ _3067_ _3069_ _3073_ _0866_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3933_ _0595_ _0596_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__and3b_1
X_6652_ _2376_ _3012_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3864_ _0530_ _0536_ net57 _0512_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5603_ _2085_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__inv_2
X_6583_ _2947_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3795_ _0443_ _0444_ inputcont.INTERNAL_SYNCED_I\[8\] vssd1 vssd1 vccd1 vccd1 _0474_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8322_ net123 _0422_ net84 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[17\] sky130_fd_sc_hd__dfrtp_1
X_5534_ pm.next_count\[0\] pm.current_waveform\[0\] _2016_ _2017_ vssd1 vssd1 vccd1
+ vccd1 _2018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8253_ net131 _0353_ net92 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[14\] sky130_fd_sc_hd__dfrtp_1
X_5465_ _1966_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__inv_2
X_8184_ net140 _0305_ net101 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[18\] sky130_fd_sc_hd__dfrtp_2
X_4416_ _0964_ _0967_ _0969_ _0973_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__o221a_1
X_7204_ _0554_ vssd1 vssd1 vccd1 vccd1 _3403_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7135_ _0559_ _3378_ sound2.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 _3381_ sky130_fd_sc_hd__a21oi_1
X_5396_ _1125_ _1780_ _1800_ _1033_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__o2bb2a_1
X_4347_ _0699_ net35 _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__a21boi_4
X_7066_ _3302_ _3313_ _3314_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__o21ba_1
X_4278_ seq.clk_div.count\[18\] _0853_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6017_ _2447_ _2449_ _2451_ _2452_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__and4_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ net130 _0131_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[23\] sky130_fd_sc_hd__dfrtp_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7899_ net107 inputcont.INTERNAL_SYNCED_I\[6\] net68 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6919_ _3190_ _3191_ vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5250_ _0575_ _0557_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4201_ _0787_ _0788_ _0790_ _0793_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__o32a_1
X_5181_ _1077_ _1562_ _1565_ _1020_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__o22a_1
X_4132_ _0742_ _0741_ _0744_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_5.next_state\[3\]
+ sky130_fd_sc_hd__o211a_1
X_4063_ _0702_ net52 vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nand2_4
XFILLER_0_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire57 _0537_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
X_7822_ net114 seq.player_3.next_state\[0\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_3.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7753_ net139 _0038_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4965_ _1511_ _1512_ _1504_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__and3b_1
X_6704_ _3058_ _3059_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__xnor2_1
X_3916_ _0512_ _0533_ _0580_ _0502_ inputcont.INTERNAL_SYNCED_I\[3\] vssd1 vssd1 vccd1
+ vccd1 _0581_ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7684_ sound4.sdiv.A\[24\] _2182_ vssd1 vssd1 vccd1 vccd1 _3738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4896_ sound2.count\[17\] _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6635_ _2996_ _2997_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3847_ _0500_ _0491_ _0475_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_116_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6566_ _2890_ _2934_ _2935_ _2894_ sound1.sdiv.A\[5\] vssd1 vssd1 vccd1 vccd1 _0113_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ inputcont.INTERNAL_SYNCED_I\[2\] _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8305_ net137 _0405_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5517_ _0552_ _2003_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8236_ net135 sound3.osc.next_count\[17\] net96 vssd1 vssd1 vccd1 vccd1 sound3.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_6497_ _1249_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5448_ _1779_ _1936_ _1952_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8167_ net140 _0288_ net101 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout100 net106 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_8
Xfanout111 net115 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_4
Xfanout122 net124 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_4
X_5379_ _1775_ _1888_ _1889_ _1774_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__o2bb2a_1
Xfanout144 net145 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_8
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
X_8098_ net136 sound2.sdiv.next_start net97 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.start
+ sky130_fd_sc_hd__dfrtp_1
X_7118_ _3365_ _3368_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__xnor2_1
X_7049_ sound2.divisor_m\[16\] sound2.divisor_m\[15\] sound2.divisor_m\[14\] _3283_
+ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _1304_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4681_ sound1.count\[12\] _1249_ _1170_ sound1.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _1252_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6420_ _2833_ _2834_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6351_ _2730_ _2734_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5302_ _1058_ _1771_ _1788_ _1111_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__o22a_1
X_6282_ _2712_ _2713_ _0569_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5233_ sound3.count\[13\] sound3.count\[14\] _1747_ vssd1 vssd1 vccd1 vccd1 _1750_
+ sky130_fd_sc_hd__and3_1
X_8021_ net126 _0163_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5164_ _0540_ _1213_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__nor2_1
X_4115_ seq.player_6.state\[2\] seq.player_6.state\[3\] _0732_ _0733_ _0700_ vssd1
+ vssd1 vccd1 vccd1 seq.player_6.next_state\[1\] sky130_fd_sc_hd__a2111oi_1
X_5095_ net64 _1567_ _1625_ _0687_ _1580_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__o221a_1
X_4046_ _0681_ _0682_ _0683_ _0684_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__o32a_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7805_ net107 seq.player_8.next_state\[3\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_8.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5997_ _2407_ _2432_ _2412_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4948_ sound2.count\[8\] _1412_ _1469_ _1470_ _1498_ vssd1 vssd1 vccd1 vccd1 _1499_
+ sky130_fd_sc_hd__o221a_1
X_7736_ net122 _0021_ net83 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[21\] sky130_fd_sc_hd__dfrtp_1
X_7667_ _3725_ _2165_ vssd1 vssd1 vccd1 vccd1 _3726_ sky130_fd_sc_hd__xnor2_1
X_4879_ _0997_ _1343_ _1333_ _1064_ _1429_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6618_ _2890_ _2981_ _2982_ _2894_ sound1.sdiv.A\[10\] vssd1 vssd1 vccd1 vccd1 _0118_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7598_ _2843_ _1820_ _3678_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__o21ai_1
X_6549_ _2903_ _2919_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__nand2_1
X_8219_ net135 sound3.osc.next_count\[0\] net96 vssd1 vssd1 vccd1 vccd1 sound3.count\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _2323_ net61 _2345_ _2355_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5851_ net30 net31 vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5782_ wave_comb.u1.A\[4\] _0573_ wave_comb.u1.next_dived _2232_ vssd1 vssd1 vccd1
+ vccd1 _0032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4802_ _1025_ _1038_ _1347_ _1333_ _0954_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__o32a_1
X_7521_ sound3.sdiv.Q\[10\] _3654_ _3643_ sound3.sdiv.Q\[9\] _3389_ vssd1 vssd1 vccd1
+ vccd1 _0349_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4733_ _1290_ _1291_ _1256_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7452_ sound3.sdiv.A\[20\] _3463_ sound3.sdiv.next_dived _3608_ vssd1 vssd1 vccd1
+ vccd1 _0326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6403_ pm.current_waveform\[6\] _2822_ _2808_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__mux2_1
X_4664_ _0958_ _1112_ _1231_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7383_ _3542_ _3545_ vssd1 vssd1 vccd1 vccd1 _3547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4595_ _1107_ _0996_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6334_ _2762_ _2763_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__or2_1
X_6265_ _2665_ _2667_ _2664_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8004_ net136 _0146_ net97 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[5\] sky130_fd_sc_hd__dfrtp_2
X_5216_ sound3.count\[6\] sound3.count\[7\] _1732_ sound3.count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1739_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6196_ _2628_ _2629_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__and2b_1
X_5147_ _1038_ _1562_ _1625_ _1025_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a211o_1
X_5078_ sound3.count\[16\] _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__xnor2_1
X_4029_ _0606_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__inv_2
XFILLER_0_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7719_ net137 _0004_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4380_ _0686_ _0675_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ sound2.count_m\[2\] _2478_ _2479_ _2483_ _2485_ vssd1 vssd1 vccd1 vccd1 _2486_
+ sky130_fd_sc_hd__a2111o_1
X_5001_ sound2.count\[15\] _1533_ _1504_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__o21ai_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6952_ sound2.divisor_m\[6\] _3212_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6883_ _3161_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
X_5903_ _2329_ _2330_ _2332_ _2338_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5834_ wave_comb.u1.M\[0\] wave_comb.u1.M\[1\] wave_comb.u1.M\[2\] wave_comb.u1.A\[10\]
+ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__nor4_1
XFILLER_0_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5765_ wave_comb.u1.M\[2\] _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7504_ _2843_ _3649_ vssd1 vssd1 vccd1 vccd1 _3650_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4716_ sound1.count\[6\] sound1.count\[7\] _1269_ sound1.count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1279_ sky130_fd_sc_hd__a31o_1
X_5696_ _2175_ _2176_ _2178_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7435_ sound3.sdiv.A\[18\] _3463_ sound3.sdiv.next_dived _3593_ vssd1 vssd1 vccd1
+ vccd1 _0324_ sky130_fd_sc_hd__a22o_1
X_4647_ _0974_ _1210_ _1010_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7366_ _3518_ _3524_ _3531_ vssd1 vssd1 vccd1 vccd1 _3532_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6317_ wave_comb.u1.Q\[7\] _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__and3_1
X_4578_ _0943_ _1012_ _1127_ _0969_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__o221a_1
X_7297_ _3468_ _3469_ vssd1 vssd1 vccd1 vccd1 _3470_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6248_ wave_comb.u1.Q\[4\] _2680_ _0645_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__mux2_1
X_6179_ _2610_ _2612_ _0569_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3880_ rate_clk.count\[1\] rate_clk.count\[0\] rate_clk.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _0550_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5550_ sound4.divisor_m\[15\] sound4.divisor_m\[14\] sound4.divisor_m\[13\] _2032_
+ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__or4_1
X_4501_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5481_ _1779_ _1936_ _1978_ _1979_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7220_ sound3.divisor_m\[3\] _3412_ _3142_ vssd1 vssd1 vccd1 vccd1 _3413_ sky130_fd_sc_hd__mux2_1
X_4432_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__buf_4
X_7151_ sound2.sdiv.Q\[7\] _3168_ _3164_ sound2.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1
+ _0247_ sky130_fd_sc_hd__a22o_1
X_4363_ seq.player_2.state\[3\] _0878_ _0932_ _0933_ _0873_ vssd1 vssd1 vccd1 vccd1
+ _0934_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6102_ sound3.count_m\[15\] vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__inv_2
X_4294_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__clkbuf_8
X_7082_ _3304_ _3313_ _3314_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__or3_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _2462_ _2465_ _2466_ _2468_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__and4bb_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7984_ net134 sound1.osc.next_count\[5\] net95 vssd1 vssd1 vccd1 vccd1 sound1.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6935_ _3203_ _3205_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6866_ _1387_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__inv_2
X_5817_ _2254_ _2260_ _2259_ _0573_ _0645_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__a311o_1
X_6797_ sound1.sdiv.Q\[24\] _2893_ _0867_ sound1.sdiv.Q\[23\] _2854_ vssd1 vssd1 vccd1
+ vccd1 _0165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5748_ sound4.sdiv.Q\[25\] _2182_ _2185_ sound4.sdiv.Q\[24\] _2205_ vssd1 vssd1 vccd1
+ vccd1 _0025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ _2159_ _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__nor2_1
X_7418_ sound3.divisor_m\[16\] sound3.divisor_m\[15\] _3561_ vssd1 vssd1 vccd1 vccd1
+ _3578_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7349_ _3448_ _3515_ vssd1 vssd1 vccd1 vccd1 _3516_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _1522_ _1523_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[8\] sky130_fd_sc_hd__nor2_1
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6720_ _3067_ _3069_ _3073_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3932_ _0545_ _0543_ _0582_ _0489_ _0508_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a311o_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6651_ _2903_ _3011_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__nand2_1
X_3863_ _0500_ _0491_ _0519_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__nor3_1
XFILLER_0_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6582_ sound1.divisor_m\[7\] _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5602_ sound4.divisor_m\[8\] _2084_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5533_ _2014_ pm.current_waveform\[2\] pm.current_waveform\[1\] _2015_ vssd1 vssd1
+ vccd1 vccd1 _2017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3794_ inputcont.INTERNAL_SYNCED_I\[11\] _0461_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__nand2_1
X_8321_ net124 _0421_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8252_ net132 _0352_ net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[13\] sky130_fd_sc_hd__dfrtp_1
X_5464_ sound4.count\[9\] _1962_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7203_ sound3.count_m\[15\] _3132_ _3402_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a21o_1
X_8183_ net135 _0304_ net96 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4415_ _0976_ _0979_ _0981_ _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5395_ net47 net63 _1788_ _0947_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__a211o_1
X_4346_ _0698_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_1
X_7134_ sound2.sdiv.C\[3\] net66 _3378_ vssd1 vssd1 vccd1 vccd1 _3380_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7065_ _3321_ _3322_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__nand2_1
X_4277_ seq.clk_div.count\[17\] seq.clk_div.count\[18\] _0850_ vssd1 vssd1 vccd1 vccd1
+ _0855_ sky130_fd_sc_hd__and3_1
X_6016_ _2450_ sound2.divisor_m\[12\] sound2.count_m\[10\] _2443_ vssd1 vssd1 vccd1
+ vccd1 _2452_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ net134 _0130_ net95 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6918_ _3183_ _3181_ _3189_ vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__a21oi_1
X_7898_ net107 inputcont.INTERNAL_SYNCED_I\[5\] net68 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6849_ sound2.divisor_m\[4\] _1441_ _2864_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4200_ seq.tempo_select.state\[0\] seq.clk_div.count\[4\] seq.clk_div.count\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__or3b_1
X_5180_ _1193_ _1559_ _1572_ _1129_ _1710_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__o221a_1
X_4131_ seq.player_5.state\[1\] seq.player_5.state\[2\] _0738_ seq.player_5.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__a31o_1
X_4062_ seq.beat\[3\] vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ net114 seq.player_4.next_state\[3\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_7752_ net139 _0037_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4964_ sound2.count\[3\] _1508_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__or2_1
X_6703_ _3050_ _3051_ _3048_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3915_ _0510_ _0514_ _0533_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__nor3_1
XFILLER_0_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7683_ _2173_ _2172_ _2169_ _2170_ _2171_ vssd1 vssd1 vccd1 vccd1 _3737_ sky130_fd_sc_hd__o2111a_1
X_4895_ _1018_ _1314_ _1316_ _0971_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6634_ _2993_ _2995_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3846_ _0515_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nor2_1
X_6565_ _2932_ _2933_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3777_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] vssd1 vssd1
+ vccd1 vccd1 _0459_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6496_ _2878_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8304_ net121 _0404_ net82 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5516_ rate_clk.count\[4\] _0551_ rate_clk.count\[5\] vssd1 vssd1 vccd1 vccd1 _2003_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8235_ net135 sound3.osc.next_count\[16\] net96 vssd1 vssd1 vccd1 vccd1 sound3.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_5447_ sound4.count\[3\] sound4.count\[4\] _1940_ sound4.count\[5\] vssd1 vssd1 vccd1
+ vccd1 _1953_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout101 net106 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_8
X_8166_ net135 _0287_ net96 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout112 net115 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_4
X_5378_ _0688_ _1771_ _1773_ _1138_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout134 net2 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_8
Xfanout145 net2 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_8
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_8
X_7117_ _3366_ _3367_ vssd1 vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__and2b_1
X_4329_ seq.beat\[3\] seq.encode.play _0884_ inputcont.INTERNAL_SYNCED_I\[7\] vssd1
+ vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__a31oi_1
X_8097_ net118 _0239_ net79 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[5\] sky130_fd_sc_hd__dfrtp_1
X_7048_ sound2.sdiv.A\[16\] _3168_ sound2.sdiv.next_dived _3307_ vssd1 vssd1 vccd1
+ vccd1 _0223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4680_ _1237_ _1071_ _1157_ sound1.count\[10\] _1250_ vssd1 vssd1 vccd1 vccd1 _1251_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6350_ _2730_ _2734_ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5301_ sound4.count\[5\] _1810_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6281_ _2684_ _2711_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5232_ sound3.count\[13\] _1747_ _1749_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[13\]
+ sky130_fd_sc_hd__a21oi_1
X_8020_ net126 _0162_ net87 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[21\] sky130_fd_sc_hd__dfrtp_1
X_5163_ _1046_ _1572_ _1550_ _0996_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__o22a_1
X_4114_ seq.player_6.state\[1\] _0730_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__nor2_1
X_5094_ _1562_ _1572_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__and2_1
X_4045_ _0682_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7804_ net107 seq.player_8.next_state\[2\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_8.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _2426_ _2431_ _2414_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__a21o_1
X_4947_ sound2.count\[11\] _1488_ _1495_ sound2.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _1498_ sky130_fd_sc_hd__a22oi_1
X_7735_ net122 _0020_ net83 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7666_ _2158_ _2163_ _2162_ vssd1 vssd1 vccd1 vccd1 _3725_ sky130_fd_sc_hd__a21o_1
X_4878_ _1116_ _1347_ _1345_ _1113_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6617_ _2970_ _2980_ _2976_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _0479_ _0478_ _0480_ net67 _0502_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__a41o_1
X_7597_ _2341_ _2005_ vssd1 vssd1 vccd1 vccd1 _3678_ sky130_fd_sc_hd__or2_1
X_6548_ sound1.divisor_m\[3\] sound1.divisor_m\[2\] sound1.divisor_m\[1\] sound1.divisor_m\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479_ _2868_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
X_8218_ net141 sound3.sdiv.next_start net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.start
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8149_ net135 _0270_ net96 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap1 _0562_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5850_ wave_comb.u1.next_dived _2273_ _2274_ _2287_ vssd1 vssd1 vccd1 vccd1 _0045_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5781_ _2229_ _2231_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4801_ _1329_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nand2_1
X_7520_ sound3.sdiv.Q\[9\] _3654_ _3643_ sound3.sdiv.Q\[8\] _3388_ vssd1 vssd1 vccd1
+ vccd1 _0348_ sky130_fd_sc_hd__a221o_1
X_4732_ sound1.count\[12\] _1287_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7451_ _3606_ _3607_ vssd1 vssd1 vccd1 vccd1 _3608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4663_ _0990_ _1062_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6402_ _2693_ _2716_ _2805_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7382_ _3542_ _3545_ vssd1 vssd1 vccd1 vccd1 _3546_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4594_ _0952_ _1019_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6333_ _2755_ _2761_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6264_ _2694_ _2695_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8003_ net135 _0145_ net96 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[4\] sky130_fd_sc_hd__dfrtp_1
X_5215_ sound3.count\[7\] sound3.count\[8\] _1735_ vssd1 vssd1 vccd1 vccd1 _1738_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_86_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6195_ _2623_ _2627_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5146_ _1245_ _1580_ _1574_ _1110_ _1676_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__o221a_1
X_5077_ _0688_ _1559_ _1591_ _1606_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__o2111a_1
X_4028_ _0587_ _0605_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__nand2_2
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ sound1.count_m\[0\] vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7718_ net137 _0003_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7649_ _3712_ _3713_ vssd1 vssd1 vccd1 vccd1 _3714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ sound2.count\[15\] _1533_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__and2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6951_ sound2.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6882_ sound2.divisor_m\[16\] _1459_ _3142_ vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__mux2_1
X_5902_ _2335_ _2336_ _2337_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__or3_1
X_5833_ _2271_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7503_ sound3.sdiv.C\[3\] _0562_ _3645_ sound3.sdiv.C\[4\] vssd1 vssd1 vccd1 vccd1
+ _3649_ sky130_fd_sc_hd__a31o_1
X_5764_ wave_comb.u1.M\[0\] wave_comb.u1.M\[1\] _2209_ vssd1 vssd1 vccd1 vccd1 _2217_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4715_ sound1.count\[7\] sound1.count\[8\] _1272_ vssd1 vssd1 vccd1 vccd1 _1278_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_71_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5695_ _2039_ _2177_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7434_ _3591_ _3592_ vssd1 vssd1 vccd1 vccd1 _3593_ sky130_fd_sc_hd__xnor2_1
X_4646_ _0990_ _0937_ _1055_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7365_ _3529_ _3530_ vssd1 vssd1 vccd1 vccd1 _3531_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4577_ _0983_ _0992_ _1146_ _0990_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6316_ wave_comb.u1.Q\[6\] _2746_ _0645_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__mux2_1
X_7296_ _3464_ _3467_ vssd1 vssd1 vccd1 vccd1 _3469_ sky130_fd_sc_hd__and2_1
X_6247_ _2678_ _2679_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__xor2_1
X_6178_ _2610_ _2612_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__nor2_1
X_5129_ _0677_ _1083_ _1550_ _1659_ _1107_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__o32a_1
XFILLER_0_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4500_ _0676_ _1052_ _1068_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5480_ sound4.count\[12\] _1973_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _1111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4431_ _0940_ _0965_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7150_ sound2.sdiv.Q\[6\] _3168_ _3164_ sound2.sdiv.Q\[5\] vssd1 vssd1 vccd1 vccd1
+ _0246_ sky130_fd_sc_hd__a22o_1
X_4362_ _0876_ _0877_ _0881_ seq.player_3.state\[3\] vssd1 vssd1 vccd1 vccd1 _0933_
+ sky130_fd_sc_hd__a22o_1
X_6101_ _2527_ _2528_ _2530_ _2536_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__or4_1
X_4293_ _0575_ _0566_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__or2_1
X_7081_ _3335_ _3336_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__nand2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ sound2.divisor_m\[5\] _2464_ _2467_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__o21a_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7983_ net134 sound1.osc.next_count\[4\] net95 vssd1 vssd1 vccd1 vccd1 sound1.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6934_ sound2.divisor_m\[5\] _3204_ vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__xnor2_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6865_ _3150_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5816_ _2254_ _2259_ _2260_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__a21oi_1
X_6796_ sound1.sdiv.Q\[23\] _2893_ _0867_ sound1.sdiv.Q\[22\] _2853_ vssd1 vssd1 vccd1
+ vccd1 _0164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5747_ sound4.count\[17\] _2201_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7417_ sound3.sdiv.A\[16\] vssd1 vssd1 vccd1 vccd1 _3577_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5678_ sound4.divisor_m\[18\] _2160_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4629_ _1165_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__inv_2
X_7348_ sound3.divisor_m\[9\] sound3.divisor_m\[8\] sound3.divisor_m\[7\] _3492_ vssd1
+ vssd1 vccd1 vccd1 _3515_ sky130_fd_sc_hd__or4_1
X_7279_ _3437_ _3452_ _3453_ _3440_ sound3.sdiv.A\[2\] vssd1 vssd1 vccd1 vccd1 _0308_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ sound2.count\[8\] _1520_ _1504_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3931_ _0515_ _0590_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__nand2_1
X_6650_ sound1.divisor_m\[13\] _3002_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__or2_1
X_3862_ _0525_ _0517_ _0513_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6581_ _2903_ _2948_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5601_ sound4.divisor_m\[7\] _2028_ _2036_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__o21a_1
X_5532_ _2015_ pm.current_waveform\[1\] vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3793_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
X_8320_ net124 _0420_ net85 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.A\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8251_ net132 _0351_ net93 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5463_ _1965_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_8182_ net140 _0303_ net101 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[16\] sky130_fd_sc_hd__dfrtp_2
X_7202_ sound3.count\[15\] _2863_ vssd1 vssd1 vccd1 vccd1 _3402_ sky130_fd_sc_hd__and2_1
X_4414_ _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__buf_4
X_5394_ _1001_ _0996_ _1784_ _1904_ _1004_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__o32a_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4345_ seq.player_1.state\[0\] _0871_ _0873_ _0915_ vssd1 vssd1 vccd1 vccd1 _0916_
+ sky130_fd_sc_hd__a22o_1
X_7133_ _3349_ _3377_ _3379_ _3174_ sound2.sdiv.C\[2\] vssd1 vssd1 vccd1 vccd1 _0236_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7064_ sound2.sdiv.A\[17\] _3320_ vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__or2_1
X_4276_ seq.clk_div.count\[17\] _0850_ _0854_ _0813_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[17\]
+ sky130_fd_sc_hd__o211a_1
X_6015_ _2448_ sound2.count_m\[12\] _2450_ sound2.divisor_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2451_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ net134 _0129_ net95 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6917_ _3183_ _3181_ _3189_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__and3_1
X_7897_ net107 inputcont.INTERNAL_SYNCED_I\[4\] net68 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6848_ _3139_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6779_ sound1.sdiv.Q\[6\] _2894_ _2890_ sound1.sdiv.Q\[5\] vssd1 vssd1 vccd1 vccd1
+ _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4130_ _0742_ _0741_ _0743_ _0719_ vssd1 vssd1 vccd1 vccd1 seq.player_5.next_state\[2\]
+ sky130_fd_sc_hd__o211a_1
X_4061_ seq.beat\[1\] seq.beat\[0\] seq.beat\[2\] vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__or3_4
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7820_ net114 seq.player_4.next_state\[2\] net75 vssd1 vssd1 vccd1 vccd1 seq.player_4.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_7751_ net139 _0036_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ sound2.count\[3\] _1508_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__and2_1
X_6702_ _3056_ _3057_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__or2b_1
X_3914_ _0579_ vssd1 vssd1 vccd1 vccd1 sound1.sdiv.next_start sky130_fd_sc_hd__inv_2
X_7682_ sound4.sdiv.A\[23\] _2184_ _3681_ _3736_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6633_ _2993_ _2995_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__or2_1
X_4894_ _0695_ _0964_ _1418_ _1317_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3845_ _0514_ _0516_ _0517_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__or4_2
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6564_ _2932_ _2933_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3776_ _0455_ _0458_ _0453_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__nand3b_2
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6495_ sound1.divisor_m\[11\] _2877_ _2864_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__mux2_1
X_8303_ net121 _0403_ net82 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[17\] sky130_fd_sc_hd__dfrtp_4
X_5515_ rate_clk.count\[4\] _0551_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8234_ net135 sound3.osc.next_count\[15\] net96 vssd1 vssd1 vccd1 vccd1 sound3.count\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ _1951_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout102 net106 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_4
X_8165_ net140 _0286_ net101 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5377_ _0869_ _1765_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__nor2_1
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_4
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_4
X_7116_ sound2.sdiv.A\[24\] _3329_ vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__nand2_1
X_4328_ seq.player_7.state\[0\] seq.player_7.state\[1\] seq.player_7.state\[2\] seq.player_7.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__or4_1
X_8096_ net118 _0238_ net79 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[4\] sky130_fd_sc_hd__dfrtp_1
Xfanout124 net2 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_4
X_7047_ _3305_ _3306_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__nor2_1
X_4259_ seq.clk_div.count\[13\] _0838_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ net131 _0112_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5300_ sound4.count\[5\] _1810_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6280_ _2684_ _2711_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5231_ sound3.count\[13\] _1747_ _1721_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__o21ai_1
X_5162_ _0944_ _1574_ _1570_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5093_ _1062_ _1565_ _1617_ _1622_ _1623_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__o221a_1
X_4113_ seq.player_6.state\[0\] seq.player_6.state\[1\] _0729_ vssd1 vssd1 vccd1 vccd1
+ _0732_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _0685_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nand2_8
X_7803_ net107 seq.player_8.next_state\[1\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_8.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5995_ _2428_ _2430_ _2394_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7734_ net118 _0019_ net79 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4946_ _1318_ _1352_ _1396_ sound2.count\[5\] _1496_ vssd1 vssd1 vccd1 vccd1 _1497_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7665_ sound4.sdiv.A\[18\] _2183_ _3681_ _3724_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__a22o_1
X_4877_ _0677_ _1083_ _1321_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6616_ _2970_ _2976_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3828_ _0472_ _0473_ _0486_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__a21boi_1
X_7596_ _3677_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__clkbuf_1
X_6547_ sound1.sdiv.A\[3\] vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3759_ _0442_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__clkbuf_8
X_6478_ sound1.divisor_m\[4\] _2867_ _2864_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__mux2_1
X_8217_ net144 _0338_ net105 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5429_ _1779_ _1936_ _1937_ _1938_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8148_ net140 _0269_ net101 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8079_ net116 _0221_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _1189_ _1333_ _1336_ _1125_ _1350_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__o221a_1
X_5780_ wave_comb.u1.A\[2\] _2224_ _2230_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__a21bo_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ sound1.count\[12\] _1287_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__and2_1
X_7450_ _3602_ _3605_ _3599_ vssd1 vssd1 vccd1 vccd1 _3607_ sky130_fd_sc_hd__a21oi_2
X_4662_ _0974_ _1058_ _1111_ _0941_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6401_ _2821_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7381_ sound3.divisor_m\[13\] _3544_ vssd1 vssd1 vccd1 vccd1 _3545_ sky130_fd_sc_hd__xnor2_1
X_4593_ _0683_ _0947_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6332_ _2755_ _2761_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6263_ _2693_ _2685_ _2689_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nand3b_1
X_8002_ net135 _0144_ net96 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[3\] sky130_fd_sc_hd__dfrtp_1
X_5214_ sound3.count\[7\] _1735_ _1737_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_6194_ _2623_ _2627_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__nor2_1
X_5145_ _0985_ _1567_ _1570_ _1238_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5076_ _1551_ _1565_ _1055_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__a21o_1
X_4027_ _0673_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__inv_2
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5978_ sound1.count_m\[16\] _2406_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__and2_1
X_7717_ net137 _0002_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4929_ _1046_ _1347_ _1393_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7648_ _2058_ _2060_ vssd1 vssd1 vccd1 vccd1 _3713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7579_ _3667_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6950_ _3164_ _3218_ _3219_ _3174_ sound2.sdiv.A\[6\] vssd1 vssd1 vccd1 vccd1 _0213_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5901_ sound4.divisor_m\[11\] sound4.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2337_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6881_ _3160_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5832_ wave_comb.u1.C\[5\] _0569_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5763_ wave_comb.u1.A\[1\] vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__inv_2
X_7502_ _2005_ _3647_ _3648_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nor3_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4714_ _1277_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5694_ sound4.sdiv.A\[25\] _2038_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7433_ _3582_ _3584_ _3581_ vssd1 vssd1 vccd1 vccd1 _3592_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4645_ _0988_ _0955_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__nand2_1
X_7364_ _3525_ _3528_ vssd1 vssd1 vccd1 vccd1 _3530_ sky130_fd_sc_hd__and2_1
X_4576_ _0994_ _1053_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6315_ _2743_ _2745_ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7295_ _3464_ _3467_ vssd1 vssd1 vccd1 vccd1 _3468_ sky130_fd_sc_hd__nor2_1
X_6246_ _2649_ _2652_ _2648_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__a21oi_1
X_6177_ _2311_ _2577_ _2611_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__o21ai_2
X_5128_ _0683_ _1562_ _1580_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__o21a_1
X_5059_ _1557_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_2 inputcont.u1.ff_intermediate\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _0685_ _0680_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__nor2_8
XFILLER_0_13_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6100_ _2533_ _2534_ _2535_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__or3_1
X_4361_ seq.player_4.state\[3\] _0888_ _0930_ _0931_ _0883_ vssd1 vssd1 vccd1 vccd1
+ _0932_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4292_ _0700_ _0864_ vssd1 vssd1 vccd1 vccd1 seq.encode.next_sequencer_on sky130_fd_sc_hd__xnor2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7080_ sound2.sdiv.A\[19\] _3329_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__nand2_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ sound2.divisor_m\[8\] sound2.count_m\[7\] vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__or2b_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7982_ net125 sound1.osc.next_count\[3\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6933_ sound2.divisor_m\[4\] _3194_ _3177_ vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__o21a_1
X_6864_ sound2.divisor_m\[9\] _3149_ _3142_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__mux2_1
X_5815_ wave_comb.u1.A\[9\] _2224_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6795_ sound1.sdiv.Q\[22\] _2893_ _0867_ sound1.sdiv.Q\[21\] _2852_ vssd1 vssd1 vccd1
+ vccd1 _0163_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5746_ sound4.sdiv.Q\[24\] _2182_ _2185_ sound4.sdiv.Q\[23\] _2204_ vssd1 vssd1 vccd1
+ vccd1 _0024_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5677_ _2036_ _2035_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7416_ sound3.sdiv.A\[16\] _3463_ sound3.sdiv.next_dived _3576_ vssd1 vssd1 vccd1
+ vccd1 _0322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4628_ _0970_ _1078_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__nand2_2
X_7347_ sound3.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 _3514_ sky130_fd_sc_hd__inv_2
X_4559_ _0994_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7278_ _3446_ _3444_ _3451_ vssd1 vssd1 vccd1 vccd1 _3453_ sky130_fd_sc_hd__nand3_1
X_6229_ _2624_ _2661_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 note4[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _0592_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or2_2
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3861_ _0515_ _0519_ _0521_ _0523_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__or4b_1
XFILLER_0_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6580_ sound1.divisor_m\[6\] _2937_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3792_ _0467_ _0470_ inputcont.INTERNAL_SYNCED_I\[12\] vssd1 vssd1 vccd1 vccd1 _0471_
+ sky130_fd_sc_hd__o21a_1
X_5600_ sound4.sdiv.A\[8\] _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__or2_1
X_5531_ pm.count\[1\] vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8250_ net129 _0350_ net90 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.Q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7201_ sound3.count_m\[14\] _3132_ _3401_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a21o_1
X_5462_ _1779_ _1936_ _1963_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8181_ net142 _0302_ net103 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4413_ _0983_ _0951_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__or2_1
X_5393_ _0869_ _1832_ _1842_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4344_ seq.player_2.state\[0\] _0876_ _0878_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7132_ _3378_ vssd1 vssd1 vccd1 vccd1 _3379_ sky130_fd_sc_hd__inv_2
X_7063_ sound2.sdiv.A\[17\] _3320_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__nand2_1
X_6014_ sound2.count_m\[11\] vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__inv_2
X_4275_ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__inv_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7965_ net130 _0128_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6916_ _3187_ _3188_ vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__or2_1
X_7896_ net114 inputcont.INTERNAL_SYNCED_I\[3\] net75 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6847_ sound2.divisor_m\[3\] _1352_ _2864_ vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6778_ sound1.sdiv.Q\[5\] _2894_ sound1.sdiv.next_dived sound1.sdiv.Q\[4\] vssd1
+ vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5729_ sound4.sdiv.Q\[16\] _2182_ _2185_ sound4.sdiv.Q\[15\] _2195_ vssd1 vssd1 vccd1
+ vccd1 _0016_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4060_ _0700_ net1 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__nor2_8
XFILLER_0_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7750_ net139 _0035_ net100 vssd1 vssd1 vccd1 vccd1 wave_comb.u1.A\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4962_ _1510_ vssd1 vssd1 vccd1 vccd1 sound2.osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_6701_ sound1.sdiv.A\[18\] _3055_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__nand2_1
X_3913_ _0575_ net65 vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nor2_4
X_7681_ _2043_ _3735_ vssd1 vssd1 vccd1 vccd1 _3736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4893_ sound2.count\[13\] _1434_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6632_ sound1.divisor_m\[12\] _2994_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3844_ _0479_ _0478_ _0485_ _0489_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6563_ _2923_ _2925_ _2922_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3775_ _0456_ inputcont.INTERNAL_SYNCED_I\[4\] _0443_ _0457_ inputcont.INTERNAL_SYNCED_I\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__o32a_1
X_6494_ _1050_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__inv_2
X_5514_ _0551_ _2002_ vssd1 vssd1 vccd1 vccd1 rate_clk.next_count\[3\] sky130_fd_sc_hd__nor2_1
X_8302_ net122 _0402_ net83 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8233_ net129 sound3.osc.next_count\[14\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_5445_ sound4.count\[4\] sound4.count\[5\] _1944_ vssd1 vssd1 vccd1 vccd1 _1951_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8164_ net135 _0285_ net96 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout103 net106 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__buf_8
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7115_ sound2.sdiv.A\[24\] _3329_ vssd1 vssd1 vccd1 vccd1 _3366_ sky130_fd_sc_hd__nor2_1
X_5376_ _1777_ _1788_ _1213_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__a21o_1
Xfanout136 net145 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_4
Xfanout125 net134 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_4
X_4327_ select1.sequencer_on _0897_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__and2_1
X_8095_ net119 _0237_ net80 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[3\] sky130_fd_sc_hd__dfrtp_2
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_4
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7046_ _3294_ _3298_ _3304_ vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__a21oi_2
X_4258_ seq.clk_div.count\[11\] seq.clk_div.count\[12\] seq.clk_div.count\[13\] _0832_
+ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4189_ seq.clk_div.count\[5\] seq.clk_div.count\[15\] seq.clk_div.count\[17\] seq.clk_div.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_69_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ net131 _0111_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7879_ net130 seq_power_on net91 vssd1 vssd1 vccd1 vccd1 seq.encode.inter_keys\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5230_ _1747_ _1748_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[12\] sky130_fd_sc_hd__nor2_1
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5161_ _1658_ _1667_ _1674_ _1683_ _1691_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__o2111ai_1
X_5092_ _1111_ _1611_ _1568_ _1058_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__o22a_1
X_4112_ seq.player_6.state\[0\] _0729_ _0731_ vssd1 vssd1 vccd1 vccd1 seq.player_6.next_state\[0\]
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4043_ _0686_ _0677_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__nor2_8
XFILLER_0_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5994_ _2409_ sound1.divisor_m\[4\] _2411_ _2429_ _2404_ vssd1 vssd1 vccd1 vccd1
+ _2430_ sky130_fd_sc_hd__o221a_1
X_7802_ net107 seq.player_8.next_state\[0\] net68 vssd1 vssd1 vccd1 vccd1 seq.player_8.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4945_ sound2.count\[11\] _1488_ _1495_ sound2.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _1496_ sky130_fd_sc_hd__o22a_1
X_7733_ net117 _0018_ net78 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7664_ _2158_ _2164_ vssd1 vssd1 vccd1 vccd1 _3724_ sky130_fd_sc_hd__xnor2_1
X_4876_ _0676_ _1322_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6615_ _2974_ _2979_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3827_ _0504_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__inv_2
X_7595_ sound4.divisor_m\[15\] _3676_ _2186_ vssd1 vssd1 vccd1 vccd1 _3677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6546_ sound1.sdiv.A\[3\] _2895_ _2916_ _2917_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a22o_1
X_3758_ inputcont.INTERNAL_SYNCED_I\[0\] inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[3\]
+ inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6477_ _1145_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__inv_2
X_8216_ net141 _0337_ net102 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[4\] sky130_fd_sc_hd__dfrtp_1
X_5428_ sound4.count\[0\] sound4.count\[1\] vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8147_ net140 _0268_ net101 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5359_ _0687_ _1001_ _1790_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8078_ net116 _0220_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[13\] sky130_fd_sc_hd__dfrtp_1
X_7029_ _3164_ _3289_ _3290_ _3174_ sound2.sdiv.A\[14\] vssd1 vssd1 vccd1 vccd1 _0221_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4730_ _1289_ vssd1 vssd1 vccd1 vccd1 sound1.osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ _0685_ _0940_ _0965_ _0964_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7380_ _3448_ _3543_ vssd1 vssd1 vccd1 vccd1 _3544_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6400_ pm.current_waveform\[5\] _2820_ _2808_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6331_ _2289_ _2758_ _2760_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__a21oi_1
X_4592_ _0677_ _0976_ _1046_ _1090_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6262_ _2685_ _2689_ _2693_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8001_ net135 _0143_ net96 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[2\] sky130_fd_sc_hd__dfrtp_1
X_5213_ sound3.count\[7\] _1735_ _1721_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__o21ai_1
X_6193_ _2279_ _2624_ _2626_ _2292_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__o22a_1
X_5144_ _1004_ _1133_ _1559_ _1565_ _0954_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__o32a_1
X_5075_ _1562_ _1548_ _1568_ _1010_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4026_ _0604_ _0595_ _0589_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ sound1.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7716_ net137 _0001_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[1\] sky130_fd_sc_hd__dfrtp_2
X_4928_ sound2.count\[1\] _1404_ _1469_ _1470_ _1478_ vssd1 vssd1 vccd1 vccd1 _1479_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7647_ _2066_ _3710_ vssd1 vssd1 vccd1 vccd1 _3712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _1004_ _1038_ _1327_ _1321_ _1154_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__o32a_1
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7578_ sound4.divisor_m\[8\] _3666_ _3419_ vssd1 vssd1 vccd1 vccd1 _3667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6529_ sound1.sdiv.A\[1\] vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5900_ sound4.divisor_m\[10\] sound4.count_m\[9\] vssd1 vssd1 vccd1 vccd1 _2336_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6880_ sound2.divisor_m\[15\] _1454_ _3142_ vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831_ _2270_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5762_ wave_comb.u1.A\[0\] _2211_ _2213_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7501_ _0562_ _3645_ sound3.sdiv.C\[3\] vssd1 vssd1 vccd1 vccd1 _3648_ sky130_fd_sc_hd__a21oi_1
X_4713_ _1256_ _1275_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5693_ sound4.sdiv.A\[24\] sound4.sdiv.A\[23\] _2038_ vssd1 vssd1 vccd1 vccd1 _2176_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7432_ _3589_ _3590_ vssd1 vssd1 vccd1 vccd1 _3591_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4644_ _0958_ _1058_ _1212_ _1214_ _1070_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7363_ _3525_ _3528_ vssd1 vssd1 vccd1 vccd1 _3529_ sky130_fd_sc_hd__nor2_1
X_4575_ _0683_ _0694_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__or2_4
X_7294_ sound3.divisor_m\[4\] _3466_ vssd1 vssd1 vccd1 vccd1 _3467_ sky130_fd_sc_hd__xor2_1
X_6314_ _2684_ _2711_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6245_ _2676_ _2677_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__xor2_1
X_6176_ _2575_ _2576_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__or2_1
X_5127_ sound3.count\[13\] vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__inv_2
X_5058_ _1059_ _1562_ _1570_ _1063_ _1588_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o221a_1
X_4009_ _0659_ _0660_ vssd1 vssd1 vccd1 vccd1 wave.next_state\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_0_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_3 inputcont.u1.ff_intermediate\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ _0886_ _0887_ _0890_ seq.player_5.state\[3\] vssd1 vssd1 vccd1 vccd1 _0931_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4291_ seq.encode.keys_edge_det\[1\] seq.encode.keys_sync\[1\] vssd1 vssd1 vccd1
+ vccd1 _0864_ sky130_fd_sc_hd__and2b_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _2461_ sound2.divisor_m\[7\] _2463_ sound2.divisor_m\[6\] vssd1 vssd1 vccd1
+ vccd1 _2466_ sky130_fd_sc_hd__o22a_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7981_ net125 sound1.osc.next_count\[2\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6932_ sound2.sdiv.A\[4\] vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6863_ _1495_ vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__inv_2
X_5814_ wave_comb.u1.A\[8\] _2224_ _2257_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__o21bai_1
X_6794_ sound1.sdiv.Q\[21\] _2893_ _0867_ sound1.sdiv.Q\[20\] _2851_ vssd1 vssd1 vccd1
+ vccd1 _0162_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5745_ sound4.count\[16\] _2201_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5676_ sound4.sdiv.A\[17\] vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7415_ _3569_ _3575_ vssd1 vssd1 vccd1 vccd1 _3576_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4627_ _0685_ _0964_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7346_ _3437_ _3512_ _3513_ _3440_ sound3.sdiv.A\[9\] vssd1 vssd1 vccd1 vccd1 _0315_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4558_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__clkbuf_8
X_7277_ _3446_ _3444_ _3451_ vssd1 vssd1 vccd1 vccd1 _3452_ sky130_fd_sc_hd__a21o_1
X_4489_ _0956_ _1026_ _1059_ _0981_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__o22a_1
X_6228_ sound2.sdiv.Q\[3\] _2660_ _2625_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__a21oi_1
X_6159_ sound2.sdiv.Q\[3\] _0578_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__nand2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 pwm_o sky130_fd_sc_hd__clkbuf_4
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 note2[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3860_ _0510_ _0514_ _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__or3_2
X_3791_ _0464_ _0443_ _0461_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or3b_1
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ pm.count\[2\] vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__inv_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5461_ sound4.count\[6\] sound4.count\[7\] _1951_ sound4.count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1964_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7200_ sound3.count\[14\] _2863_ vssd1 vssd1 vccd1 vccd1 _3401_ sky130_fd_sc_hd__and2_1
X_4412_ _0674_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__nor2_8
XFILLER_0_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8180_ net140 _0301_ net101 vssd1 vssd1 vccd1 vccd1 sound3.divisor_m\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5392_ _0993_ _1837_ _1900_ _1902_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7131_ sound2.sdiv.C\[2\] sound2.sdiv.C\[1\] sound2.sdiv.C\[0\] vssd1 vssd1 vccd1
+ vccd1 _3378_ sky130_fd_sc_hd__and3_1
X_4343_ seq.player_3.state\[0\] _0881_ _0883_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_
+ sky130_fd_sc_hd__a22o_1
X_4274_ seq.clk_div.count\[15\] seq.clk_div.count\[16\] seq.clk_div.count\[17\] _0844_
+ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__and4_1
X_7062_ _3319_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6013_ sound2.count_m\[13\] _2441_ _2448_ sound2.count_m\[12\] vssd1 vssd1 vccd1
+ vccd1 _2449_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7964_ net130 _0127_ net91 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[19\] sky130_fd_sc_hd__dfrtp_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6915_ _3184_ _3186_ vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7895_ net114 inputcont.INTERNAL_SYNCED_I\[2\] net75 vssd1 vssd1 vccd1 vccd1 seq.encode.keys_edge_det\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6846_ _3138_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6777_ sound1.sdiv.Q\[4\] _2894_ sound1.sdiv.next_dived sound1.sdiv.Q\[3\] vssd1
+ vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ pm.count\[1\] pm.count\[0\] pm.count\[2\] vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5728_ sound4.count\[8\] _2186_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5659_ sound4.divisor_m\[14\] vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7329_ _3486_ _3490_ _3497_ vssd1 vssd1 vccd1 vccd1 _3499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _1508_ _1504_ _1509_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__and3b_1
X_6700_ sound1.sdiv.A\[18\] _3055_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7680_ sound4.sdiv.A\[21\] _2038_ _3733_ vssd1 vssd1 vccd1 vccd1 _3735_ sky130_fd_sc_hd__a21oi_1
X_3912_ _0578_ vssd1 vssd1 vccd1 vccd1 sound2.sdiv.next_start sky130_fd_sc_hd__inv_2
X_4892_ _1423_ _1424_ _1434_ sound2.count\[13\] _1442_ vssd1 vssd1 vccd1 vccd1 _1443_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6631_ sound1.divisor_m\[11\] _2984_ _2903_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3843_ _0478_ _0485_ _0479_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6562_ _2930_ _2931_ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3774_ inputcont.INTERNAL_SYNCED_I\[1\] inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1
+ vccd1 vccd1 _0457_ sky130_fd_sc_hd__nor2_1
X_8301_ net122 _0401_ net83 vssd1 vssd1 vccd1 vccd1 sound4.divisor_m\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6493_ _2876_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5513_ rate_clk.count\[3\] _0550_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8232_ net129 sound3.osc.next_count\[13\] net90 vssd1 vssd1 vccd1 vccd1 sound3.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5444_ _1950_ vssd1 vssd1 vccd1 vccd1 sound4.osc.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
X_8163_ net140 _0284_ net101 vssd1 vssd1 vccd1 vccd1 sound3.count_m\[16\] sky130_fd_sc_hd__dfrtp_1
Xfanout104 net105 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__buf_6
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7114_ _3360_ _3363_ _3359_ vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__o21a_1
X_5375_ _1867_ _1868_ _1876_ _1877_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__a221o_1
Xfanout126 net134 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_4
Xfanout137 net145 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_4
Xfanout115 net2 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
X_4326_ seq.beat\[3\] seq.encode.play _0879_ inputcont.INTERNAL_SYNCED_I\[6\] vssd1
+ vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__a31o_1
X_8094_ net119 _0236_ net80 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.C\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7045_ _3294_ _3298_ _3304_ vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__and3_1
X_4257_ _0840_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
X_4188_ seq.tempo_select.state\[1\] seq.tempo_select.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _0782_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7947_ net131 _0110_ net92 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.A\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7878_ net114 seq_play_on net75 vssd1 vssd1 vccd1 vccd1 seq.encode.inter_keys\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6829_ sound2.count\[14\] _2855_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ sound3.count\[10\] _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__xnor2_1
X_5091_ _0695_ _0540_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__nor2_1
X_4111_ seq.player_6.state\[1\] seq.player_6.state\[2\] seq.player_6.state\[3\] _0730_
+ _0700_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__a311o_1
XFILLER_0_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4042_ _0676_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__inv_6
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _2416_ _2418_ _2410_ sound1.divisor_m\[3\] vssd1 vssd1 vccd1 vccd1 _2429_
+ sky130_fd_sc_hd__o2bb2a_1
X_7801_ net113 oct.next_state\[2\] net74 vssd1 vssd1 vccd1 vccd1 oct.state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7732_ net120 _0017_ net81 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[17\] sky130_fd_sc_hd__dfrtp_1
X_4944_ _1490_ _1492_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7663_ sound4.sdiv.A\[17\] _2183_ sound4.sdiv.next_dived _3723_ vssd1 vssd1 vccd1
+ vccd1 _0422_ sky130_fd_sc_hd__a22o_1
X_4875_ _1341_ _1372_ _1425_ _1107_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__a31o_1
X_6614_ sound1.divisor_m\[10\] _2978_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3826_ _0500_ _0475_ _0491_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__a31oi_4
X_7594_ _1891_ vssd1 vssd1 vccd1 vccd1 _3676_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6545_ _2909_ _2915_ _0866_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ inputcont.INTERNAL_SYNCED_I\[10\] vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8215_ net144 _0336_ net105 vssd1 vssd1 vccd1 vccd1 sound3.sdiv.C\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6476_ _2005_ _1208_ _2866_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5427_ sound4.count\[0\] sound4.count\[1\] vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8146_ net117 _0267_ net78 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[27\] sky130_fd_sc_hd__dfrtp_1
X_5358_ _0683_ _1769_ _1794_ _0996_ _1800_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__o221a_1
X_8077_ net116 _0219_ net77 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.A\[12\] sky130_fd_sc_hd__dfrtp_1
X_4309_ _0702_ seq.encode.play _0879_ inputcont.INTERNAL_SYNCED_I\[2\] vssd1 vssd1
+ vccd1 vccd1 _0880_ sky130_fd_sc_hd__a31o_1
X_7028_ _3277_ _3280_ _3288_ vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__a21o_1
X_5289_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _1229_ _1230_ _0695_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6330_ _2759_ _2753_ sound2.sdiv.Q\[8\] _2295_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__a2bb2o_1
X_4591_ _0969_ _1004_ _1038_ _1077_ _1000_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__o32a_1
XFILLER_0_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6261_ _2289_ _2691_ _2692_ _2293_ sound1.sdiv.Q\[6\] vssd1 vssd1 vccd1 vccd1 _2693_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8000_ net140 _0142_ net101 vssd1 vssd1 vccd1 vccd1 sound1.sdiv.Q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5212_ _1735_ _1736_ vssd1 vssd1 vccd1 vccd1 sound3.osc.next_count\[6\] sky130_fd_sc_hd__nor2_1
X_6192_ _2594_ _2625_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__xor2_1
X_5143_ sound3.count\[1\] _1673_ _1635_ sound3.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _1674_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5074_ sound3.count\[17\] _1604_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__xor2_1
X_4025_ _0667_ _0670_ _0672_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__o21ai_4
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ sound1.count_m\[17\] _2405_ sound1.count_m\[18\] vssd1 vssd1 vccd1 vccd1 _2412_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7715_ net137 _0000_ net98 vssd1 vssd1 vccd1 vccd1 sound4.sdiv.Q\[0\] sky130_fd_sc_hd__dfrtp_1
X_4927_ sound2.count\[0\] _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4858_ _1025_ _1046_ _1339_ _1322_ _1164_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__o32a_1
XFILLER_0_51_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7646_ _3681_ _3710_ _3711_ _2184_ sound4.sdiv.A\[12\] vssd1 vssd1 vccd1 vccd1 _0417_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3809_ _0474_ _0475_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nor2_1
X_7577_ _1829_ vssd1 vssd1 vccd1 vccd1 _3666_ sky130_fd_sc_hd__inv_2
X_4789_ _1331_ _1324_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__or2_1
X_6528_ sound1.divisor_m\[0\] sound1.sdiv.Q\[27\] _2898_ _2900_ vssd1 vssd1 vccd1
+ vccd1 _2901_ sky130_fd_sc_hd__a31oi_2
X_6459_ _0575_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__buf_6
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8129_ net112 _0250_ net73 vssd1 vssd1 vccd1 vccd1 sound2.sdiv.Q\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5830_ wave_comb.u1.C\[4\] _0569_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__and2_1
X_5761_ wave_comb.u1.next_dived _2213_ _2214_ _0573_ wave_comb.u1.A\[1\] vssd1 vssd1
+ vccd1 vccd1 _0029_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7500_ sound3.sdiv.C\[3\] _0562_ _3645_ vssd1 vssd1 vccd1 vccd1 _3647_ sky130_fd_sc_hd__and3_1
X_4712_ sound1.count\[7\] _1272_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7431_ _3586_ _3588_ vssd1 vssd1 vccd1 vccd1 _3590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5692_ sound4.sdiv.A\[24\] _2038_ _2174_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4643_ _0990_ _0941_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7362_ sound3.divisor_m\[11\] _3527_ vssd1 vssd1 vccd1 vccd1 _3528_ sky130_fd_sc_hd__xnor2_1
X_4574_ _1070_ _1132_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__and3_2
XFILLER_0_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7293_ _3448_ _3465_ vssd1 vssd1 vccd1 vccd1 _3466_ sky130_fd_sc_hd__nand2_1
X_6313_ _2710_ _2708_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__and2b_1
X_6244_ _2631_ _2637_ _2638_ _2644_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6175_ _2607_ _2609_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5126_ sound3.count\[5\] _1635_ _1641_ sound3.count\[3\] _1656_ vssd1 vssd1 vccd1
+ vccd1 _1657_ sky130_fd_sc_hd__a221o_1
X_5057_ _0679_ net63 _1550_ _1580_ _1053_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__o32a_1
X_4008_ inputcont.INTERNAL_MODE _0658_ wave.mode\[0\] vssd1 vssd1 vccd1 vccd1 _0660_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5959_ sound1.divisor_m\[8\] vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7629_ _3681_ _3698_ _3699_ _2184_ sound4.sdiv.A\[7\] vssd1 vssd1 vccd1 vccd1 _0412_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 inputcont.u1.ff_intermediate\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ seq.encode.play _0863_ vssd1 vssd1 vccd1 vccd1 seq.encode.next_play sky130_fd_sc_hd__xnor2_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7980_ net125 sound1.osc.next_count\[1\] net86 vssd1 vssd1 vccd1 vccd1 sound1.count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6931_ _3200_ _3202_ sound2.sdiv.A\[4\] _3168_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a2bb2o_1
X_6862_ _3148_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5813_ wave_comb.u1.A\[9\] _0573_ wave_comb.u1.next_dived _2258_ vssd1 vssd1 vccd1
+ vccd1 _0037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6793_ sound1.sdiv.Q\[20\] _2893_ _0867_ sound1.sdiv.Q\[19\] _2850_ vssd1 vssd1 vccd1
+ vccd1 _0161_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ sound4.sdiv.Q\[23\] _2182_ _2185_ sound4.sdiv.Q\[22\] _2203_ vssd1 vssd1 vccd1
+ vccd1 _0023_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5675_ _2049_ _2053_ _2152_ _2157_ _2155_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__a221o_1
X_7414_ _3573_ _3574_ vssd1 vssd1 vccd1 vccd1 _3575_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4626_ sound1.count\[9\] _1196_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7345_ _3503_ _3507_ _3510_ _3511_ vssd1 vssd1 vccd1 vccd1 _3513_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4557_ _0995_ _0947_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__or2_1
X_7276_ _3447_ _3450_ vssd1 vssd1 vccd1 vccd1 _3451_ sky130_fd_sc_hd__xnor2_1
X_4488_ _1018_ _0959_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6227_ _0578_ _2499_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__and2_1
X_6158_ sound2.sdiv.Q\[2\] _0578_ _2591_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__a21oi_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _1146_ _1572_ _1574_ _1125_ _1639_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__o221a_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ sound3.count_m\[10\] vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 mode_out[0] sky130_fd_sc_hd__buf_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 note2[2] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 seq_led_on sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3790_ _0469_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5460_ _1962_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4411_ _0676_ _0680_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__nand2_4
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5391_ _0997_ _1769_ _1792_ _1010_ _1901_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7130_ sound2.sdiv.C\[1\] sound2.sdiv.C\[0\] sound2.sdiv.C\[2\] vssd1 vssd1 vccd1
+ vccd1 _3377_ sky130_fd_sc_hd__a21o_1
X_4342_ seq.player_4.state\[0\] _0886_ _0888_ _0912_ vssd1 vssd1 vccd1 vccd1 _0913_
+ sky130_fd_sc_hd__a22o_1
X_4273_ _0852_ vssd1 vssd1 vccd1 vccd1 seq.clk_div.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
X_7061_ sound2.divisor_m\[18\] _3318_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__xnor2_1
X_6012_ sound2.divisor_m\[13\] vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__inv_2
.ends

