* NGSPICE file created from synth.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt synth VGND VPWR clk en keypad_i[0] keypad_i[10] keypad_i[11] keypad_i[12]
+ keypad_i[13] keypad_i[14] keypad_i[1] keypad_i[2] keypad_i[3] keypad_i[4] keypad_i[5]
+ keypad_i[6] keypad_i[7] keypad_i[8] keypad_i[9] n_rst pwm_o sound_series[0] sound_series[1]
+ sound_series[2] sound_series[3]
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1270_ _0583_ _0584_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1606_ _0147_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_0985_ kp_encoder.sync_out\[4\] kp_encoder.sync_out\[5\] kp_encoder.sync_out\[6\]
+ kp_encoder.sync_out\[7\] VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or4b_1
X_1468_ net114 _0632_ _0634_ seq_div.R\[21\] VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1537_ _0106_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
X_1399_ _0709_ seq_div.R\[8\] _0707_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1253_ clk8.count\[19\] clk8.count\[18\] _0567_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__and3_1
X_1322_ _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__clkbuf_8
X_1184_ clk8.count\[3\] clk8.count\[2\] clk8.count\[4\] clk8.count\[5\] VGND VGND
+ VPWR VPWR _0523_ sky130_fd_sc_hd__or4b_1
XFILLER_0_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0968_ kp_encoder.sync_out\[4\] kp_encoder.sync_out\[5\] kp_encoder.sync_out\[6\]
+ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or3b_1
XFILLER_0_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0899_ _0260_ _0272_ _0238_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0822_ _0154_ _0184_ _0196_ SS_FSM.count\[2\] VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1236_ clk8.count\[12\] clk8.count\[13\] _0553_ clk8.count\[14\] VGND VGND VPWR VPWR
+ _0561_ sky130_fd_sc_hd__a31o_1
X_1305_ pwm.count\[5\] _0597_ _0593_ pwm.count\[6\] _0620_ VGND VGND VPWR VPWR _0621_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1167_ _0510_ _0511_ _0331_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__and3b_1
X_1098_ _0463_ VGND VGND VPWR VPWR osc.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ _0375_ _0391_ _0382_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1785_ clknet_4_3_0_clk net55 net30 VGND VGND VPWR VPWR kp_encoder.last_sk sky130_fd_sc_hd__dfrtp_1
X_0805_ SS_FSM.count\[6\] SS_FSM.count\[7\] VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1219_ clk8.count\[9\] _0546_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold63 clk8.count\[13\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 seq_div.Q\[2\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 clk8.count\[3\] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 SS_FSM.count\[7\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold30 seq_div.dividend\[0\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold85 seq_div.dividend\[0\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _0237_ _0214_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__nor2_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _0348_ _0349_ _0350_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1768_ clknet_4_10_0_clk net8 net34 VGND VGND VPWR VPWR kp_encoder.q\[1\] sky130_fd_sc_hd__dfrtp_1
X_1699_ clknet_4_1_0_clk _0055_ net29 VGND VGND VPWR VPWR SS_FSM.count\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR sound_series[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1622_ clknet_4_3_0_clk SS_FSM.next_sound\[1\] net30 VGND VGND VPWR VPWR SS_FSM.sound\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_1484_ _0778_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
X_1553_ _0179_ _0117_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__nand2_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0984_ kp_encoder.sync_out\[2\] kp_encoder.sync_out\[3\] VGND VGND VPWR VPWR _0355_
+ sky130_fd_sc_hd__nor2_1
X_1605_ net130 osc.count\[14\] _0132_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_1
X_1536_ seq_div.D\[11\] _0105_ _0631_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_1
X_1467_ _0765_ seq_div.R\[20\] _0707_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1398_ seq_div.D\[0\] _0695_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1252_ _0572_ VGND VGND VPWR VPWR clk8.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
X_1321_ _0626_ _0631_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__nor2_1
X_1183_ net61 _0519_ _0522_ VGND VGND VPWR VPWR pwm.next_count\[7\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0967_ kp_encoder.sync_out\[10\] VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1519_ _0435_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
X_0898_ _0232_ _0268_ _0271_ _0175_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0821_ SS_FSM.count\[3\] VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1235_ clk8.count\[13\] clk8.count\[14\] _0556_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__and3_1
X_1304_ pwm.count\[4\] _0601_ _0597_ pwm.count\[5\] _0619_ VGND VGND VPWR VPWR _0620_
+ sky130_fd_sc_hd__o221a_1
X_1166_ pwm.count\[0\] pwm.count\[1\] pwm.count\[2\] VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1097_ _0461_ _0417_ _0448_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__and4b_1
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1020_ _0361_ _0377_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1784_ clknet_4_7_0_clk net50 net31 VGND VGND VPWR VPWR kp_encoder.last_mk sky130_fd_sc_hd__dfrtp_1
X_0804_ SS_FSM.count\[0\] VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1218_ _0548_ VGND VGND VPWR VPWR clk8.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_1149_ net93 _0497_ _0499_ VGND VGND VPWR VPWR clk_div.next_count\[4\] sky130_fd_sc_hd__o21a_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold64 clk8.next_count\[13\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0029_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 pwm.count\[0\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 seq_div.dividend\[10\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _0003_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 seq_div.dividend\[1\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 seq_div.dividend\[4\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1003_ _0351_ _0361_ _0370_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_16_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1698_ clknet_4_1_0_clk _0054_ net28 VGND VGND VPWR VPWR SS_FSM.count\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1767_ clknet_4_10_0_clk net2 net34 VGND VGND VPWR VPWR kp_encoder.q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput21 net21 VGND VGND VPWR VPWR sound_series[2] sky130_fd_sc_hd__clkbuf_4
X_1621_ clknet_4_3_0_clk SS_FSM.next_sound\[0\] net30 VGND VGND VPWR VPWR SS_FSM.sound\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_1552_ _0172_ _0173_ _0269_ _0116_ _0236_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__a41o_1
XFILLER_0_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1483_ seq_div.Q\[1\] seq_div.q_out\[1\] _0776_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__mux2_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0983_ kp_encoder.sync_out\[9\] VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__inv_2
X_1604_ _0146_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_1535_ _0395_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
X_1466_ _0671_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__xnor2_1
X_1397_ net68 _0632_ _0634_ seq_div.R\[8\] _0708_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1320_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__buf_6
X_1182_ net61 _0519_ _0331_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__o21ai_1
X_1251_ _0570_ _0531_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and3b_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0897_ _0167_ _0269_ _0270_ _0264_ _0214_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__a2111o_1
X_0966_ kp_encoder.sync_out\[8\] _0334_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1449_ _0749_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1518_ _0094_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0820_ _0179_ _0162_ _0165_ _0183_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__or4_4
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1303_ pwm.count\[3\] _0605_ _0601_ pwm.count\[4\] _0618_ VGND VGND VPWR VPWR _0619_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1234_ net101 _0556_ _0559_ VGND VGND VPWR VPWR clk8.next_count\[13\] sky130_fd_sc_hd__o21a_1
X_1165_ pwm.count\[2\] pwm.count\[0\] pwm.count\[1\] VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1096_ osc.count\[5\] _0458_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0949_ _0159_ _0314_ _0316_ _0320_ _0214_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o311a_1
X_1783_ clknet_4_15_0_clk net7 net38 VGND VGND VPWR VPWR kp_encoder.q\[14\] sky130_fd_sc_hd__dfrtp_1
X_0803_ _0177_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1217_ _0546_ _0531_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__and3b_1
X_1148_ net93 _0497_ _0350_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__a21oi_1
X_1079_ osc.count\[0\] osc.count\[1\] VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold21 seq_div.Q\[7\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 seq_div.Q\[0\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 seq_div.dividend\[13\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 clk_div.count\[3\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 clk8.count\[4\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 seq_div.dividend\[11\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _0013_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 kp_encoder.q\[2\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ net1 _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__and2_2
XFILLER_0_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1766_ clknet_4_15_0_clk net46 net38 VGND VGND VPWR VPWR kp_encoder.sync_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1697_ clknet_4_1_0_clk _0053_ net29 VGND VGND VPWR VPWR SS_FSM.count\[2\] sky130_fd_sc_hd__dfstp_4
XFILLER_0_12_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR sound_series[3] sky130_fd_sc_hd__buf_2
X_1620_ clknet_4_13_0_clk _0002_ net37 VGND VGND VPWR VPWR seq_div.count_div\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1482_ _0777_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
X_1551_ _0196_ _0193_ _0222_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__or3_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1749_ clknet_4_5_0_clk clk8.next_count\[18\] net32 VGND VGND VPWR VPWR clk8.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0982_ net20 _0344_ _0346_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__or3_1
X_1603_ net129 osc.count\[13\] _0132_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
X_1465_ _0701_ _0760_ _0676_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__o21ai_2
X_1534_ _0104_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1396_ _0707_ _0628_ seq_div.D\[0\] VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and3b_1
XFILLER_0_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1250_ clk8.count\[18\] _0567_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or2_1
X_1181_ _0521_ VGND VGND VPWR VPWR pwm.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0965_ _0335_ kp_encoder.sync_out\[11\] kp_encoder.sync_out\[12\] VGND VGND VPWR
+ VPWR _0336_ sky130_fd_sc_hd__or3b_1
X_0896_ _0154_ SS_FSM.count\[5\] VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__nor2_1
X_1448_ _0691_ _0742_ _0661_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1517_ seq_div.D\[4\] _0093_ _0632_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_1
X_1379_ _0640_ _0659_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1233_ clk8.count\[13\] _0556_ _0531_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__a21boi_1
X_1302_ pwm.count\[2\] _0609_ _0605_ pwm.count\[3\] _0617_ VGND VGND VPWR VPWR _0618_
+ sky130_fd_sc_hd__o221a_1
X_1164_ net58 net71 _0509_ VGND VGND VPWR VPWR pwm.next_count\[1\] sky130_fd_sc_hd__a21oi_1
X_1095_ osc.count\[5\] osc.count\[4\] _0455_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0948_ _0317_ _0318_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0879_ SS_FSM.count\[3\] _0162_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0802_ _0157_ _0158_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1782_ clknet_4_7_0_clk net6 net31 VGND VGND VPWR VPWR kp_encoder.q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1216_ clk8.count\[7\] clk8.count\[6\] _0540_ clk8.count\[8\] VGND VGND VPWR VPWR
+ _0547_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1147_ net70 _0494_ _0498_ VGND VGND VPWR VPWR clk_div.next_count\[3\] sky130_fd_sc_hd__o21a_1
X_1078_ _0331_ net97 _0417_ _0448_ VGND VGND VPWR VPWR osc.next_count\[0\] sky130_fd_sc_hd__nand4_1
Xhold22 _0034_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 kp_encoder.q\[0\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 _0028_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 pwm.count\[1\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 clk_div.count\[4\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 seq_div.D\[12\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 seq_div.dividend\[1\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 seq_div.D\[0\] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1001_ _0334_ _0344_ _0346_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a31o_1
X_1765_ clknet_4_7_0_clk net43 net31 VGND VGND VPWR VPWR kp_encoder.sync_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1696_ clknet_4_0_0_clk _0052_ net28 VGND VGND VPWR VPWR SS_FSM.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1481_ net120 seq_div.q_out\[0\] _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__mux2_1
X_1550_ _0240_ _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__nor2_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1748_ clknet_4_5_0_clk clk8.next_count\[17\] net32 VGND VGND VPWR VPWR clk8.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1679_ clknet_4_9_0_clk _0035_ net33 VGND VGND VPWR VPWR seq_div.D\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0981_ _0344_ _0346_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__nand2_2
X_1602_ _0145_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1464_ _0628_ _0762_ _0763_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1533_ net119 _0103_ _0631_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1395_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__buf_6
XFILLER_0_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1180_ _0519_ _0331_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0964_ kp_encoder.sync_out\[8\] kp_encoder.sync_out\[9\] kp_encoder.sync_out\[10\]
+ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1516_ _0381_ _0392_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__nand2_1
X_0895_ SS_FSM.count\[3\] _0190_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__or2_2
X_1447_ _0689_ _0658_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__nor2_1
X_1378_ _0664_ _0689_ _0658_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1232_ _0558_ VGND VGND VPWR VPWR clk8.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
X_1301_ pwm.count\[1\] _0615_ _0609_ pwm.count\[2\] _0616_ VGND VGND VPWR VPWR _0617_
+ sky130_fd_sc_hd__a221o_1
X_1163_ pwm.count\[0\] net71 _0331_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__o21ai_1
X_1094_ _0460_ VGND VGND VPWR VPWR osc.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0947_ _0167_ _0195_ _0213_ _0159_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0878_ _0228_ _0248_ _0251_ _0178_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1781_ clknet_4_5_0_clk net5 net31 VGND VGND VPWR VPWR kp_encoder.q\[12\] sky130_fd_sc_hd__dfrtp_1
X_0801_ _0169_ net25 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1215_ clk8.count\[7\] clk8.count\[8\] _0543_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1146_ _0350_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1077_ _0443_ _0445_ _0405_ _0413_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_7_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold12 kp_encoder.sync_out\[13\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 pwm.count\[7\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 pwm.next_count\[1\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 clk_div.count\[1\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 seq_div.dividend\[4\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 clk8.count\[16\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 SS_FSM.count\[8\] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 seq_div.dividend\[5\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ _0327_ _0329_ _0344_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1764_ clknet_4_6_0_clk net51 net30 VGND VGND VPWR VPWR kp_encoder.sync_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1695_ clknet_4_0_0_clk _0051_ net28 VGND VGND VPWR VPWR SS_FSM.count\[0\] sky130_fd_sc_hd__dfrtp_4
X_1129_ _0485_ _0417_ _0448_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__and4b_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1480_ seq_div.state\[1\] seq_div.state\[0\] VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nand2_4
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1678_ clknet_4_13_0_clk net60 net37 VGND VGND VPWR VPWR seq_div.Q\[7\] sky130_fd_sc_hd__dfrtp_1
X_1747_ clknet_4_5_0_clk clk8.next_count\[16\] net32 VGND VGND VPWR VPWR clk8.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0980_ _0348_ _0349_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a21o_1
X_1601_ seq_div.dividend\[12\] osc.count\[12\] _0132_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__mux2_1
X_1532_ _0411_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1463_ seq_div.dividend\[12\] _0632_ _0634_ seq_div.R\[20\] VGND VGND VPWR VPWR _0763_
+ sky130_fd_sc_hd__a22o_1
X_1394_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0894_ _0178_ _0265_ _0267_ _0176_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a211o_1
X_0963_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or2_1
X_1515_ _0092_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
X_1377_ _0636_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__inv_2
X_1446_ net88 _0712_ _0717_ seq_div.R\[17\] _0748_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1231_ _0556_ _0331_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__and3b_1
X_1300_ pwm.count\[0\] _0592_ _0610_ _0614_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__o31a_1
X_1162_ _0350_ net58 VGND VGND VPWR VPWR pwm.next_count\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1093_ _0458_ _0417_ _0448_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__and4b_1
XFILLER_0_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0877_ _0249_ _0250_ _0228_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o21ai_1
X_0946_ _0205_ _0288_ _0228_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1429_ _0628_ _0733_ _0734_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0800_ SS_FSM.count\[8\] _0171_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__a21o_4
X_1780_ clknet_4_1_0_clk net4 net29 VGND VGND VPWR VPWR kp_encoder.q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ net106 _0543_ _0545_ VGND VGND VPWR VPWR clk8.next_count\[7\] sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1145_ clk_div.count\[3\] _0494_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1076_ _0409_ _0446_ _0412_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__or3b_1
X_0929_ _0178_ _0300_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or2_1
Xhold24 seq_div.Q\[5\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold68 clk8.count\[7\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 seq_div.count_div\[1\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 kp_encoder.q\[12\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 seq_div.state\[1\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 clk_div.next_count\[1\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 seq_div.dividend\[11\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1694_ clknet_4_12_0_clk _0050_ net35 VGND VGND VPWR VPWR seq_div.D\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1763_ clknet_4_3_0_clk net47 net30 VGND VGND VPWR VPWR kp_encoder.sync_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1128_ osc.count\[13\] _0482_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1059_ _0383_ _0378_ _0429_ _0382_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o22ai_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1746_ clknet_4_5_0_clk clk8.next_count\[15\] net32 VGND VGND VPWR VPWR clk8.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1677_ clknet_4_13_0_clk net63 net36 VGND VGND VPWR VPWR seq_div.Q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1462_ _0761_ seq_div.R\[19\] _0707_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__mux2_1
X_1600_ _0144_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_1531_ _0102_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1393_ seq_div.R\[23\] _0681_ _0682_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__and4b_1
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1729_ clknet_4_7_0_clk pwm.next_count\[6\] net31 VGND VGND VPWR VPWR pwm.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0962_ kp_encoder.sync_out\[4\] kp_encoder.sync_out\[5\] kp_encoder.sync_out\[6\]
+ kp_encoder.sync_out\[7\] VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or4_1
X_0893_ _0228_ _0261_ _0253_ _0266_ _0178_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a311oi_1
X_1445_ seq_div.R\[16\] _0707_ _0747_ _0625_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a211o_1
X_1514_ seq_div.D\[3\] _0091_ _0632_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1376_ _0684_ _0686_ _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1230_ clk8.count\[12\] _0553_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or2_1
X_1161_ _0508_ VGND VGND VPWR VPWR clk_div.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1092_ osc.count\[4\] _0455_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0945_ _0189_ _0186_ _0205_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o21a_1
X_0876_ _0154_ _0155_ _0196_ SS_FSM.count\[2\] VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1428_ net78 _0632_ _0634_ seq_div.R\[14\] VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__a22o_1
X_1359_ _0668_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1213_ clk8.count\[7\] clk8.count\[6\] _0540_ _0350_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__a31o_1
X_1144_ _0496_ VGND VGND VPWR VPWR clk_div.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1075_ _0393_ _0407_ osc.count\[8\] VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0859_ _0180_ _0206_ _0178_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__or3_2
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ _0185_ _0270_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nand2_1
Xhold25 _0033_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _0629_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _0076_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 kp_encoder.q\[8\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 seq_div.dividend\[2\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 seq_div.dividend\[5\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1693_ clknet_4_12_0_clk _0049_ net35 VGND VGND VPWR VPWR seq_div.D\[14\] sky130_fd_sc_hd__dfrtp_1
X_1762_ clknet_4_2_0_clk net42 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1127_ osc.count\[13\] _0482_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__and2_1
X_1058_ _0361_ _0377_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1745_ clknet_4_5_0_clk clk8.next_count\[14\] net32 VGND VGND VPWR VPWR clk8.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1676_ clknet_4_15_0_clk _0032_ net37 VGND VGND VPWR VPWR seq_div.Q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1461_ _0701_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__xor2_1
X_1530_ seq_div.D\[9\] _0101_ _0631_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1392_ _0683_ _0688_ _0693_ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1728_ clknet_4_7_0_clk pwm.next_count\[5\] net31 VGND VGND VPWR VPWR pwm.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ clknet_4_1_0_clk clk_div.next_count\[4\] net30 VGND VGND VPWR VPWR clk_div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0961_ kp_encoder.sync_out\[0\] kp_encoder.sync_out\[1\] kp_encoder.sync_out\[2\]
+ kp_encoder.sync_out\[3\] VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0892_ _0184_ SS_FSM.count\[2\] _0166_ _0196_ _0154_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1444_ _0707_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__nor2_1
X_1513_ _0420_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
X_1375_ _0647_ _0651_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1160_ _0331_ _0506_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__and3_1
X_1091_ osc.count\[4\] osc.count\[3\] _0452_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0944_ _0249_ _0315_ _0228_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0875_ _0209_ _0210_ _0165_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a21oi_2
X_1358_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__inv_2
X_1427_ _0732_ seq_div.R\[13\] _0707_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__mux2_1
X_1289_ seq_div.q_out\[3\] _0588_ _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1212_ _0543_ _0544_ VGND VGND VPWR VPWR clk8.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1143_ _0494_ _0331_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and3b_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1074_ _0418_ _0419_ _0441_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0927_ _0179_ _0184_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0789_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[2\] SS_FSM.count\[3\] VGND VGND VPWR
+ VPWR _0164_ sky130_fd_sc_hd__o31a_2
XFILLER_0_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0858_ _0176_ _0227_ _0231_ _0159_ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o221a_1
Xhold37 seq_div.Q\[3\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 clk_div.count\[0\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 seq_div.count_div\[0\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 osc.count\[0\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 kp_encoder.q\[1\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1761_ clknet_4_3_0_clk net54 net30 VGND VGND VPWR VPWR kp_encoder.sync_out\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1692_ clknet_4_12_0_clk _0048_ net35 VGND VGND VPWR VPWR seq_div.D\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1126_ _0484_ VGND VGND VPWR VPWR osc.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1057_ osc.count\[1\] _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1744_ clknet_4_5_0_clk net102 net29 VGND VGND VPWR VPWR clk8.count\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1675_ clknet_4_15_0_clk _0031_ net37 VGND VGND VPWR VPWR seq_div.Q\[4\] sky130_fd_sc_hd__dfrtp_1
X_1109_ _0470_ _0417_ _0448_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1460_ _0693_ _0741_ _0758_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1391_ _0696_ _0700_ _0701_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__or4b_1
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1727_ clknet_4_7_0_clk pwm.next_count\[4\] net31 VGND VGND VPWR VPWR pwm.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_1658_ clknet_4_4_0_clk clk_div.next_count\[3\] net30 VGND VGND VPWR VPWR clk_div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1589_ net78 osc.count\[6\] _0132_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0960_ net1 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1512_ _0090_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0891_ _0167_ _0195_ _0263_ _0264_ _0225_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a32o_1
X_1443_ _0691_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__xor2_1
X_1374_ _0643_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1090_ _0457_ VGND VGND VPWR VPWR osc.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
X_0943_ _0210_ _0262_ _0189_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__a21oi_1
X_0874_ _0165_ _0244_ _0195_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1288_ _0582_ _0602_ _0603_ _0591_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__a31o_1
X_1357_ seq_div.D\[13\] seq_div.R\[20\] VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__and2b_1
X_1426_ _0699_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1142_ clk_div.count\[1\] clk_div.count\[0\] clk_div.count\[2\] VGND VGND VPWR VPWR
+ _0495_ sky130_fd_sc_hd__a21o_1
X_1211_ clk8.count\[6\] _0540_ _0531_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1073_ _0438_ _0436_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__nand2_1
X_0857_ _0171_ _0216_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__nand2_2
X_0926_ _0240_ _0236_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold38 _0030_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 kp_encoder.q\[9\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 clk8.count\[1\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ net96 _0712_ _0716_ _0625_ _0718_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__o221a_1
X_0788_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[3\] SS_FSM.count\[2\] VGND VGND VPWR
+ VPWR _0163_ sky130_fd_sc_hd__nor4_4
Xhold49 seq_div.D\[6\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1691_ clknet_4_14_0_clk _0047_ net37 VGND VGND VPWR VPWR seq_div.D\[12\] sky130_fd_sc_hd__dfrtp_1
X_1760_ clknet_4_3_0_clk net52 net30 VGND VGND VPWR VPWR kp_encoder.sync_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1125_ _0482_ _0417_ _0448_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__and4b_1
XFILLER_0_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ _0375_ _0425_ _0426_ _0420_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a31o_1
X_0909_ _0178_ _0279_ _0281_ _0214_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1743_ clknet_4_7_0_clk clk8.next_count\[12\] net31 VGND VGND VPWR VPWR clk8.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1674_ clknet_4_13_0_clk net76 net37 VGND VGND VPWR VPWR seq_div.Q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1039_ _0375_ _0361_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__nand2_1
X_1108_ osc.count\[8\] _0467_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1390_ seq_div.D\[15\] seq_div.R\[22\] VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1726_ clknet_4_7_0_clk pwm.next_count\[3\] net31 VGND VGND VPWR VPWR pwm.count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_1657_ clknet_4_4_0_clk clk_div.next_count\[2\] net30 VGND VGND VPWR VPWR clk_div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1588_ _0138_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0890_ _0166_ _0249_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1442_ _0660_ _0742_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__nand2_1
X_1511_ seq_div.D\[2\] _0089_ _0632_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1373_ _0645_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1709_ clknet_4_9_0_clk _0065_ net33 VGND VGND VPWR VPWR seq_div.dividend\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 net32 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_6
XFILLER_0_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ _0228_ _0248_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nor2_1
X_0873_ _0241_ _0243_ _0245_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1425_ _0654_ _0727_ _0650_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__a21o_1
X_1287_ _0585_ seq_div.q_out\[2\] VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__nand2_1
X_1356_ seq_div.R\[20\] seq_div.D\[13\] VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1210_ clk8.count\[6\] _0540_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__and2_1
X_1141_ clk_div.count\[1\] clk_div.count\[0\] clk_div.count\[2\] VGND VGND VPWR VPWR
+ _0494_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1072_ _0418_ _0419_ _0424_ _0433_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0925_ _0175_ _0296_ _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0787_ _0160_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__and2_2
X_0856_ _0169_ _0165_ _0228_ _0229_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__o41a_1
Xhold39 seq_div.Q\[4\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 kp_encoder.sync_out\[14\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 clk8.next_count\[1\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ seq_div.R\[10\] _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__or2_1
X_1339_ seq_div.D\[4\] seq_div.R\[11\] VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1690_ clknet_4_12_0_clk _0046_ net37 VGND VGND VPWR VPWR seq_div.D\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1124_ osc.count\[12\] _0479_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__or2_1
X_1055_ _0361_ _0370_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput18 net18 VGND VGND VPWR VPWR pwm_o sky130_fd_sc_hd__clkbuf_4
X_0839_ SS_FSM.count\[6\] net24 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__xnor2_4
X_0908_ _0167_ _0187_ _0192_ _0280_ _0159_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1673_ clknet_4_13_0_clk net80 net36 VGND VGND VPWR VPWR seq_div.Q\[2\] sky130_fd_sc_hd__dfrtp_1
X_1742_ clknet_4_7_0_clk clk8.next_count\[11\] net31 VGND VGND VPWR VPWR clk8.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1038_ osc.count\[8\] _0393_ _0407_ _0408_ osc.count\[9\] VGND VGND VPWR VPWR _0409_
+ sky130_fd_sc_hd__a32o_1
X_1107_ osc.count\[8\] _0467_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1725_ clknet_4_7_0_clk pwm.next_count\[2\] net31 VGND VGND VPWR VPWR pwm.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1656_ clknet_4_6_0_clk net95 net30 VGND VGND VPWR VPWR clk_div.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1587_ net127 osc.count\[5\] _0132_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1510_ _0422_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
X_1441_ net99 _0712_ _0717_ seq_div.R\[16\] _0744_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__o221a_1
X_1372_ _0644_ _0648_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__or2b_1
X_1708_ clknet_4_9_0_clk _0064_ net33 VGND VGND VPWR VPWR seq_div.dividend\[4\] sky130_fd_sc_hd__dfrtp_1
X_1639_ clknet_4_3_0_clk osc.next_count\[0\] net30 VGND VGND VPWR VPWR osc.count\[0\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout31 net32 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_4
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0941_ _0310_ _0312_ _0175_ _0232_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a211o_1
X_0872_ _0167_ _0195_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__nor2_1
X_1355_ _0635_ _0665_ _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__and3_1
X_1424_ _0628_ _0729_ _0730_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a21o_1
X_1286_ _0585_ seq_div.q_out\[2\] VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1140_ net94 net64 _0493_ VGND VGND VPWR VPWR clk_div.next_count\[1\] sky130_fd_sc_hd__o21a_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1071_ _0434_ _0436_ _0438_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__or4bb_1
X_0924_ SS_FSM.count\[3\] SS_FSM.count\[2\] _0234_ _0175_ VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_11_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0786_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[2\] VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__o21ai_2
X_0855_ _0209_ _0210_ _0167_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a21o_1
Xhold29 pwm.count\[7\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 clk8.count\[20\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1407_ _0625_ _0712_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__nand2_2
X_1338_ seq_div.D\[5\] seq_div.R\[12\] VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__and2b_1
X_1269_ seq_div.q_out\[7\] VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1123_ osc.count\[12\] osc.count\[11\] _0476_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and3_1
X_1054_ _0361_ _0370_ _0382_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__o21ai_1
X_0907_ _0189_ _0229_ _0228_ _0209_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__o211a_1
Xoutput19 net19 VGND VGND VPWR VPWR sound_series[0] sky130_fd_sc_hd__clkbuf_4
X_0838_ _0166_ _0212_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2_1
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1741_ clknet_4_5_0_clk clk8.next_count\[10\] net29 VGND VGND VPWR VPWR clk8.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1672_ clknet_4_13_0_clk net82 net36 VGND VGND VPWR VPWR seq_div.Q\[1\] sky130_fd_sc_hd__dfrtp_1
X_1106_ _0469_ VGND VGND VPWR VPWR osc.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1037_ _0374_ _0394_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1724_ clknet_4_6_0_clk net72 net31 VGND VGND VPWR VPWR pwm.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ clknet_4_7_0_clk clk_div.next_count\[0\] net30 VGND VGND VPWR VPWR clk_div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1586_ _0137_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ _0650_ _0654_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__or2b_1
X_1440_ seq_div.R\[15\] _0707_ _0742_ _0743_ _0625_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1638_ clknet_4_12_0_clk _0018_ net37 VGND VGND VPWR VPWR seq_div.R\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1707_ clknet_4_8_0_clk _0063_ net33 VGND VGND VPWR VPWR seq_div.dividend\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1569_ SS_FSM.count\[5\] _0123_ _0127_ _0128_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__o22a_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout32 net17 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
XFILLER_0_44_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0940_ _0201_ _0257_ _0311_ _0187_ _0176_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0871_ _0205_ _0165_ _0159_ _0244_ _0214_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1285_ seq_div.q_out\[4\] _0588_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o21ai_1
X_1354_ seq_div.R\[19\] seq_div.D\[12\] VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or2b_1
X_1423_ net107 _0632_ _0634_ seq_div.R\[13\] VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1070_ _0418_ _0419_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0923_ _0282_ _0287_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0854_ _0179_ _0162_ _0183_ _0190_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__o31a_1
XFILLER_0_11_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0785_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[2\] VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__or3_2
XFILLER_0_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1268_ mode_FSM.mode\[1\] seq_div.q_out\[6\] mode_FSM.mode\[0\] VGND VGND VPWR VPWR
+ _0584_ sky130_fd_sc_hd__o21a_1
Xhold19 seq_div.count_div\[2\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ _0715_ seq_div.R\[9\] _0707_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__mux2_1
X_1337_ _0646_ _0647_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1199_ _0534_ _0331_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ _0481_ VGND VGND VPWR VPWR osc.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
X_1053_ osc.count\[3\] _0420_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0837_ _0196_ _0160_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0906_ _0167_ _0276_ _0277_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1740_ clknet_4_4_0_clk clk8.next_count\[9\] net29 VGND VGND VPWR VPWR clk8.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1671_ clknet_4_13_0_clk _0027_ net35 VGND VGND VPWR VPWR seq_div.Q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ _0467_ _0417_ _0448_ _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__and4b_1
X_1036_ _0379_ _0406_ _0382_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1723_ clknet_4_6_0_clk pwm.next_count\[0\] net36 VGND VGND VPWR VPWR pwm.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1654_ clknet_4_6_0_clk osc.next_count\[15\] net35 VGND VGND VPWR VPWR osc.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1585_ net124 osc.count\[4\] _0132_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1019_ _0375_ _0370_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1370_ _0678_ seq_div.R\[22\] VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1637_ clknet_4_15_0_clk _0017_ net37 VGND VGND VPWR VPWR seq_div.R\[22\] sky130_fd_sc_hd__dfrtp_2
X_1706_ clknet_4_8_0_clk _0062_ net33 VGND VGND VPWR VPWR seq_div.dividend\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1499_ seq_div.Q\[1\] _0628_ _0634_ net79 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a22o_1
X_1568_ _0237_ _0159_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__nor2_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout33 net38 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_6
XFILLER_0_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0870_ _0219_ _0222_ _0223_ _0185_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a31o_1
X_1422_ _0728_ seq_div.R\[12\] _0707_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__mux2_1
X_1284_ _0582_ _0598_ _0599_ _0591_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__a31o_1
X_1353_ _0636_ _0662_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0999_ _0352_ _0362_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ _0176_ _0290_ _0291_ _0294_ _0217_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__o311a_1
X_0853_ _0205_ net26 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__xnor2_4
X_0784_ _0157_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__nor2_8
X_1405_ _0686_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1267_ seq_div.q_out\[6\] _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__nand2_1
Xinput1 en VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
X_1198_ clk8.count\[1\] clk8.count\[0\] clk8.count\[2\] VGND VGND VPWR VPWR _0535_
+ sky130_fd_sc_hd__a21o_1
X_1336_ seq_div.R\[10\] seq_div.D\[3\] VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1121_ _0479_ _0417_ _0448_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__and4b_1
X_1052_ osc.count\[3\] _0420_ _0422_ osc.count\[2\] VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0836_ SS_FSM.count\[4\] net27 _0164_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or4_2
X_0905_ SS_FSM.count\[4\] _0156_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nor2_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1670_ clknet_4_13_0_clk _0026_ net36 VGND VGND VPWR VPWR seq_div.q_out\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1104_ osc.count\[7\] _0464_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or2_1
X_1035_ _0351_ _0361_ _0377_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__nand3_2
XFILLER_0_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0819_ _0154_ SS_FSM.count\[3\] _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1722_ clknet_4_13_0_clk pwm.pwm net36 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1653_ clknet_4_6_0_clk osc.next_count\[14\] net35 VGND VGND VPWR VPWR osc.count\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1584_ _0136_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ osc.count\[12\] _0385_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1705_ clknet_4_8_0_clk _0061_ net33 VGND VGND VPWR VPWR seq_div.dividend\[1\] sky130_fd_sc_hd__dfrtp_1
X_1636_ clknet_4_15_0_clk _0016_ net37 VGND VGND VPWR VPWR seq_div.R\[21\] sky130_fd_sc_hd__dfrtp_1
X_1567_ SS_FSM.count\[4\] _0123_ _0126_ _0127_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__o22a_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1498_ net81 _0628_ _0634_ seq_div.Q\[1\] VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__a22o_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout34 net38 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_6
XFILLER_0_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1421_ _0683_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__xnor2_1
X_1283_ _0585_ seq_div.q_out\[3\] VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__nand2_1
X_1352_ _0635_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0998_ _0344_ _0346_ _0368_ _0350_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__a31o_1
X_1619_ clknet_4_15_0_clk _0001_ net37 VGND VGND VPWR VPWR seq_div.count_div\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0921_ _0178_ _0207_ _0245_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a211o_1
X_0783_ SS_FSM.count\[4\] _0156_ SS_FSM.count\[5\] VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__o21a_2
X_0852_ _0167_ _0226_ _0211_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1404_ _0713_ _0694_ _0642_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1335_ seq_div.R\[11\] seq_div.D\[4\] VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__or2b_1
X_1266_ _0581_ mode_FSM.mode\[0\] VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__and2_2
X_1197_ clk8.count\[1\] clk8.count\[0\] clk8.count\[2\] VGND VGND VPWR VPWR _0534_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 keypad_i[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1120_ osc.count\[11\] _0476_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or2_1
X_1051_ _0375_ _0391_ _0421_ _0377_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0904_ _0206_ _0191_ _0156_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0835_ _0179_ _0155_ _0193_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__or3_2
X_1318_ _0623_ seq_div.state\[0\] VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1249_ clk8.count\[18\] _0567_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__and2_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1034_ _0388_ _0389_ _0396_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or4b_2
X_1103_ osc.count\[7\] osc.count\[6\] _0461_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0818_ SS_FSM.count\[2\] VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1721_ clknet_4_12_0_clk _0077_ net37 VGND VGND VPWR VPWR seq_div.state\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ clknet_4_3_0_clk osc.next_count\[13\] net35 VGND VGND VPWR VPWR osc.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1583_ seq_div.dividend\[3\] osc.count\[3\] _0132_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1017_ osc.count\[12\] _0385_ _0387_ osc.count\[13\] VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1704_ clknet_4_8_0_clk _0060_ net33 VGND VGND VPWR VPWR seq_div.dividend\[0\] sky130_fd_sc_hd__dfrtp_1
X_1497_ _0625_ _0707_ _0634_ net81 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a2bb2o_1
X_1635_ clknet_4_14_0_clk _0015_ net37 VGND VGND VPWR VPWR seq_div.R\[20\] sky130_fd_sc_hd__dfrtp_1
X_1566_ _0174_ _0299_ _0115_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__a21o_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout35 net38 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_6
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1351_ seq_div.D\[11\] seq_div.R\[18\] VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or2b_1
X_1420_ _0687_ _0723_ _0651_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__o21ai_1
X_1282_ _0585_ seq_div.q_out\[3\] VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1618_ clknet_4_15_0_clk _0000_ net37 VGND VGND VPWR VPWR seq_div.count_div\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0997_ kp_encoder.sync_out\[9\] _0337_ _0343_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__a211o_1
X_1549_ _0350_ _0529_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0920_ _0195_ _0292_ _0167_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a21oi_1
X_0782_ SS_FSM.count\[4\] SS_FSM.count\[5\] _0156_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__nor3_4
XFILLER_0_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0851_ _0179_ _0221_ _0225_ _0159_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__o22a_1
X_1265_ mode_FSM.mode\[1\] VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__inv_2
X_1334_ _0642_ _0643_ _0644_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__a211o_1
X_1403_ seq_div.D\[0\] VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__inv_2
X_1196_ net65 clk8.count\[0\] _0533_ VGND VGND VPWR VPWR clk8.next_count\[1\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 keypad_i[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1050_ _0375_ _0361_ _0382_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0903_ _0179_ _0165_ _0186_ _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__o31a_1
X_0834_ _0156_ _0180_ _0181_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or3_2
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1248_ _0569_ VGND VGND VPWR VPWR clk8.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_1317_ net57 _0627_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ pwm.count\[6\] _0516_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or2_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1102_ _0466_ VGND VGND VPWR VPWR osc.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_1033_ _0399_ _0400_ _0401_ _0403_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__and4b_1
XFILLER_0_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0817_ _0189_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1720_ clknet_4_13_0_clk net74 net38 VGND VGND VPWR VPWR seq_div.state\[0\] sky130_fd_sc_hd__dfrtp_4
X_1651_ clknet_4_3_0_clk osc.next_count\[12\] net35 VGND VGND VPWR VPWR osc.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _0135_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1016_ _0375_ _0379_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1703_ clknet_4_1_0_clk _0059_ net29 VGND VGND VPWR VPWR SS_FSM.count\[8\] sky130_fd_sc_hd__dfstp_1
X_1634_ clknet_4_14_0_clk _0014_ net37 VGND VGND VPWR VPWR seq_div.R\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1496_ _0085_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1565_ _0237_ _0167_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__nor2_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout36 net38 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
XFILLER_0_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1281_ seq_div.q_out\[5\] _0588_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__o21ai_1
X_1350_ _0641_ _0657_ _0658_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0996_ _0332_ _0356_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o21ai_1
X_1617_ _0153_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1479_ _0628_ _0774_ net109 VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a21o_1
X_1548_ _0113_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0850_ _0189_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or2_1
X_1402_ _0623_ seq_div.state\[0\] VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__nand2_4
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0781_ SS_FSM.count\[0\] _0155_ SS_FSM.count\[3\] SS_FSM.count\[2\] VGND VGND VPWR
+ VPWR _0156_ sky130_fd_sc_hd__or4_4
XFILLER_0_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1264_ _0274_ _0577_ _0578_ SS_FSM.sound\[1\] VGND VGND VPWR VPWR SS_FSM.next_sound\[1\]
+ sky130_fd_sc_hd__a22o_1
Xinput4 keypad_i[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_1333_ seq_div.D\[2\] seq_div.R\[9\] VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__and2b_1
X_1195_ net65 clk8.count\[0\] _0331_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0979_ net1 VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkinv_8
XFILLER_0_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0833_ _0178_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__nor2_1
X_0902_ _0179_ _0184_ SS_FSM.count\[3\] VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1247_ _0567_ _0531_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__and3b_1
X_1178_ pwm.count\[6\] _0516_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and2_1
X_1316_ _0627_ net85 VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1032_ osc.count\[14\] _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1101_ _0464_ _0417_ _0448_ _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and4b_1
XFILLER_0_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0816_ _0162_ _0183_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1650_ clknet_4_3_0_clk osc.next_count\[11\] net30 VGND VGND VPWR VPWR osc.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1581_ net128 osc.count\[2\] _0132_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1015_ _0373_ _0361_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1779_ clknet_4_0_0_clk net3 net28 VGND VGND VPWR VPWR kp_encoder.q\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1702_ clknet_4_4_0_clk _0058_ net29 VGND VGND VPWR VPWR SS_FSM.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_1633_ clknet_4_14_0_clk net92 net37 VGND VGND VPWR VPWR seq_div.R\[18\] sky130_fd_sc_hd__dfrtp_1
X_1564_ SS_FSM.count\[3\] _0115_ _0119_ _0125_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a22o_1
X_1495_ net59 _0585_ _0776_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout37 net38 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1280_ _0582_ _0594_ _0595_ _0591_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0995_ kp_encoder.sync_out\[4\] _0363_ _0332_ _0365_ kp_encoder.sync_out\[0\] VGND
+ VGND VPWR VPWR _0366_ sky130_fd_sc_hd__o32a_1
X_1616_ mode_FSM.mode\[0\] _0581_ _0151_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_1
X_1547_ seq_div.D\[15\] _0112_ _0631_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_1
X_1478_ seq_div.dividend\[15\] _0632_ _0633_ net108 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0780_ SS_FSM.count\[1\] VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__buf_4
X_1401_ _0628_ _0710_ _0711_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a21o_1
Xinput5 keypad_i[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_1194_ _0532_ VGND VGND VPWR VPWR clk8.next_count\[0\] sky130_fd_sc_hd__clkbuf_1
X_1263_ _0580_ VGND VGND VPWR VPWR SS_FSM.next_sound\[0\] sky130_fd_sc_hd__clkbuf_1
X_1332_ seq_div.D\[3\] seq_div.R\[10\] VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0978_ net21 _0344_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0901_ _0240_ SS_FSM.sound\[1\] VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__nor2_1
X_0832_ _0206_ _0191_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nor2_1
X_1315_ seq_div.count_div\[0\] _0628_ net84 VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1246_ clk8.count\[15\] clk8.count\[16\] _0560_ clk8.count\[17\] VGND VGND VPWR VPWR
+ _0568_ sky130_fd_sc_hd__a31o_1
X_1177_ _0518_ VGND VGND VPWR VPWR pwm.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap23 _0120_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1100_ osc.count\[6\] _0461_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__or2_1
X_1031_ _0375_ _0386_ _0381_ _0383_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0815_ _0154_ _0155_ SS_FSM.count\[2\] VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__or3_2
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1229_ clk8.count\[12\] _0553_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1580_ _0134_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1014_ _0374_ _0376_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1778_ clknet_4_15_0_clk net16 net38 VGND VGND VPWR VPWR kp_encoder.q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1701_ clknet_4_1_0_clk _0057_ net30 VGND VGND VPWR VPWR SS_FSM.count\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1494_ _0084_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1632_ clknet_4_14_0_clk net89 net34 VGND VGND VPWR VPWR seq_div.R\[17\] sky130_fd_sc_hd__dfrtp_1
X_1563_ _0165_ _0117_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__nand2_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout38 net17 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_6
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0994_ _0364_ kp_encoder.sync_out\[3\] kp_encoder.sync_out\[1\] VGND VGND VPWR VPWR
+ _0365_ sky130_fd_sc_hd__a21oi_1
X_1615_ _0152_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1477_ _0773_ seq_div.R\[22\] _0707_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__mux2_1
X_1546_ _0382_ _0397_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1400_ net113 _0632_ _0634_ seq_div.R\[9\] VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__a22o_1
X_1331_ seq_div.R\[9\] seq_div.D\[2\] VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or2b_1
Xinput6 keypad_i[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_1193_ clk8.count\[0\] _0531_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and2b_1
X_1262_ _0578_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__and2_1
X_0977_ _0336_ _0344_ _0346_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__nand4_2
XFILLER_0_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1529_ _0408_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0155_ _0159_ _0168_ _0273_ _0240_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__a311o_2
X_0831_ _0205_ _0165_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1314_ _0626_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1245_ clk8.count\[16\] clk8.count\[17\] _0563_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__and3_1
X_1176_ _0516_ _0331_ _0517_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap24 net25 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1030_ osc.count\[13\] _0387_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0814_ _0188_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1228_ _0555_ VGND VGND VPWR VPWR clk8.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1159_ clk_div.count\[7\] _0503_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1013_ _0378_ _0379_ _0381_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1777_ clknet_4_14_0_clk net15 net37 VGND VGND VPWR VPWR kp_encoder.q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1700_ clknet_4_1_0_clk _0056_ net29 VGND VGND VPWR VPWR SS_FSM.count\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1631_ clknet_4_11_0_clk net100 net34 VGND VGND VPWR VPWR seq_div.R\[16\] sky130_fd_sc_hd__dfrtp_1
X_1493_ seq_div.Q\[6\] seq_div.q_out\[6\] _0776_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
X_1562_ _0124_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 net17 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_6
XFILLER_0_4_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0993_ kp_encoder.sync_out\[2\] VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__inv_2
X_1614_ mode_FSM.mode\[1\] mode_FSM.mode\[0\] _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1545_ _0111_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
X_1476_ _0702_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1261_ SS_FSM.sound\[0\] _0577_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__or2_1
X_1330_ seq_div.D\[1\] seq_div.R\[8\] VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__and2b_1
Xinput7 keypad_i[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_1192_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__buf_2
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0976_ _0332_ _0333_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1459_ _0664_ _0689_ _0658_ _0661_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__or4b_1
X_1528_ _0100_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0830_ SS_FSM.count\[4\] VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1244_ net105 _0563_ _0566_ VGND VGND VPWR VPWR clk8.next_count\[16\] sky130_fd_sc_hd__o21ba_1
X_1313_ seq_div.count_div\[0\] seq_div.count_div\[1\] _0626_ VGND VGND VPWR VPWR _0627_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1175_ pwm.count\[4\] pwm.count\[3\] _0510_ pwm.count\[5\] VGND VGND VPWR VPWR _0517_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0959_ _0330_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xmax_cap25 _0157_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 keypad_i[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
X_0813_ _0163_ _0164_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1227_ _0553_ _0331_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__and3b_1
X_1158_ clk_div.count\[7\] _0503_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__or2_1
X_1089_ _0455_ _0417_ _0448_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__and4b_1
XFILLER_0_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1012_ _0382_ _0375_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1776_ clknet_4_2_0_clk net14 net17 VGND VGND VPWR VPWR kp_encoder.q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1630_ clknet_4_11_0_clk _0010_ net34 VGND VGND VPWR VPWR seq_div.R\[15\] sky130_fd_sc_hd__dfrtp_1
X_1492_ _0083_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ SS_FSM.count\[2\] _0121_ _0123_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout29 net32 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_6
X_1759_ clknet_4_2_0_clk net44 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0992_ kp_encoder.sync_out\[5\] VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__inv_2
X_1613_ kp_encoder.last_mk kp_encoder.sync_out\[13\] VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__and2b_1
X_1544_ seq_div.D\[14\] _0402_ _0631_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_1475_ _0672_ _0768_ _0679_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1191_ _0331_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and2_1
X_1260_ SS_FSM.sound\[0\] _0577_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__nand2_1
Xinput8 keypad_i[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0975_ SS_FSM.sound\[1\] _0298_ _0345_ SS_FSM.sound\[0\] VGND VGND VPWR VPWR _0346_
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1527_ seq_div.D\[8\] _0099_ _0632_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_1
X_1389_ _0666_ _0676_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__nand2_1
X_1458_ _0635_ _0658_ _0663_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1243_ clk8.count\[15\] clk8.count\[16\] _0560_ _0350_ VGND VGND VPWR VPWR _0566_
+ sky130_fd_sc_hd__a31o_1
X_1174_ pwm.count\[5\] pwm.count\[4\] _0513_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1312_ _0623_ seq_div.state\[0\] VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0958_ _0327_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0889_ _0219_ _0261_ _0262_ _0210_ _0189_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap26 net27 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput11 keypad_i[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0812_ _0179_ _0165_ _0186_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1226_ clk8.count\[9\] clk8.count\[10\] _0546_ clk8.count\[11\] VGND VGND VPWR VPWR
+ _0554_ sky130_fd_sc_hd__a31o_1
X_1157_ _0505_ VGND VGND VPWR VPWR clk_div.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_1088_ osc.count\[3\] _0452_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ net1 _0372_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__nand2_4
XFILLER_0_56_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1775_ clknet_4_2_0_clk net13 net28 VGND VGND VPWR VPWR kp_encoder.q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1209_ _0542_ VGND VGND VPWR VPWR clk8.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1560_ _0122_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1491_ net62 seq_div.q_out\[5\] _0776_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux2_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1689_ clknet_4_14_0_clk _0045_ net38 VGND VGND VPWR VPWR seq_div.D\[10\] sky130_fd_sc_hd__dfrtp_1
X_1758_ clknet_4_2_0_clk net45 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0991_ net19 _0344_ _0346_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__or3_2
X_1474_ _0628_ _0770_ _0771_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a21o_1
X_1612_ _0623_ _0132_ _0634_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__o21ai_1
X_1543_ _0110_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1190_ clk8.count\[1\] clk8.count\[0\] _0523_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__or4b_1
Xinput9 keypad_i[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0974_ _0297_ _0313_ _0326_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1457_ _0628_ _0756_ _0757_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__a21o_1
X_1526_ _0393_ _0407_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__nand2_1
X_1388_ _0697_ _0655_ _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1311_ net86 _0625_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__xnor2_1
X_1242_ _0565_ VGND VGND VPWR VPWR clk8.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
X_1173_ pwm.count\[4\] _0513_ _0515_ VGND VGND VPWR VPWR pwm.next_count\[4\] sky130_fd_sc_hd__o21ba_1
X_0957_ _0206_ _0328_ _0299_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0888_ _0162_ _0183_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1509_ _0088_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap27 _0163_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0811_ _0162_ _0183_ _0185_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__o21ba_2
Xinput12 keypad_i[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1225_ clk8.count\[11\] clk8.count\[10\] _0549_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__and3_1
X_1156_ _0503_ _0331_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__and3b_1
X_1087_ osc.count\[3\] _0452_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1774_ clknet_4_0_0_clk net12 net28 VGND VGND VPWR VPWR kp_encoder.q\[5\] sky130_fd_sc_hd__dfrtp_1
X_1208_ _0540_ _0541_ _0531_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1139_ net94 clk_div.count\[0\] _0350_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1490_ _0082_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1 kp_encoder.q\[4\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1688_ clknet_4_11_0_clk _0044_ net38 VGND VGND VPWR VPWR seq_div.D\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1757_ clknet_4_0_0_clk net41 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1611_ net73 _0149_ _0150_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0990_ _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__buf_4
X_1473_ net111 _0632_ _0634_ seq_div.R\[22\] VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__a22o_1
X_1542_ seq_div.D\[13\] _0109_ _0631_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0973_ kp_encoder.sync_out\[9\] _0337_ _0341_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a211o_2
X_1456_ net117 _0632_ _0634_ seq_div.R\[19\] VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__a22o_1
X_1387_ _0653_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__nand2_1
X_1525_ _0098_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1241_ _0563_ _0531_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__and3b_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1310_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__clkbuf_4
X_1172_ pwm.count\[4\] pwm.count\[3\] _0510_ _0350_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0956_ SS_FSM.count\[5\] _0302_ _0219_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0887_ _0179_ _0183_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__nor2_1
X_1508_ seq_div.D\[1\] _0087_ _0632_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_1
X_1439_ _0692_ _0741_ _0706_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 keypad_i[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_0810_ _0184_ _0160_ _0161_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ net110 _0549_ _0552_ VGND VGND VPWR VPWR clk8.next_count\[10\] sky130_fd_sc_hd__o21ba_1
X_1155_ clk_div.count\[6\] _0500_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or2_1
X_1086_ _0454_ VGND VGND VPWR VPWR osc.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0939_ _0189_ _0186_ _0178_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1773_ clknet_4_7_0_clk _0079_ net36 VGND VGND VPWR VPWR mode_FSM.mode\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1207_ clk8.count\[3\] clk8.count\[4\] _0534_ clk8.count\[5\] VGND VGND VPWR VPWR
+ _0541_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1138_ _0350_ net64 VGND VGND VPWR VPWR clk_div.next_count\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_0_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1069_ _0382_ _0375_ _0391_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2 kp_encoder.q\[3\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1756_ clknet_4_2_0_clk net39 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1687_ clknet_4_9_0_clk _0043_ net34 VGND VGND VPWR VPWR seq_div.D\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1610_ seq_div.count_div\[0\] seq_div.count_div\[1\] net57 _0625_ VGND VGND VPWR
+ VPWR _0150_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1472_ _0769_ seq_div.R\[21\] _0707_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__mux2_1
X_1541_ _0387_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1739_ clknet_4_4_0_clk clk8.next_count\[8\] net29 VGND VGND VPWR VPWR clk8.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0972_ _0342_ _0335_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1524_ seq_div.D\[7\] _0419_ _0632_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_1
X_1455_ _0755_ seq_div.R\[18\] _0707_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__mux2_1
X_1386_ seq_div.D\[6\] seq_div.R\[13\] VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ clk8.count\[15\] _0560_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__or2_1
X_1171_ _0513_ _0514_ VGND VGND VPWR VPWR pwm.next_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0955_ _0297_ _0313_ _0326_ _0237_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ _0247_ _0259_ _0217_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1507_ _0427_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1369_ _0677_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1438_ _0692_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 keypad_i[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
X_1223_ clk8.count\[9\] clk8.count\[10\] _0546_ _0350_ VGND VGND VPWR VPWR _0552_
+ sky130_fd_sc_hd__a31o_1
X_1154_ clk_div.count\[6\] _0500_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1085_ _0452_ _0417_ _0448_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0869_ _0154_ _0242_ _0159_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a21o_1
X_0938_ _0305_ _0309_ _0214_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1772_ clknet_4_7_0_clk _0078_ net36 VGND VGND VPWR VPWR mode_FSM.mode\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1206_ clk8.count\[4\] clk8.count\[5\] _0537_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__and3_1
X_1137_ _0492_ VGND VGND VPWR VPWR osc.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1068_ osc.count\[6\] VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 kp_encoder.q\[5\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1755_ clknet_4_2_0_clk net40 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1686_ clknet_4_11_0_clk _0042_ net34 VGND VGND VPWR VPWR seq_div.D\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1540_ _0108_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1471_ _0674_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1669_ clknet_4_13_0_clk _0025_ net36 VGND VGND VPWR VPWR seq_div.q_out\[6\] sky130_fd_sc_hd__dfrtp_1
X_1738_ clknet_4_5_0_clk clk8.next_count\[7\] net29 VGND VGND VPWR VPWR clk8.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0971_ kp_encoder.sync_out\[11\] VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1454_ _0664_ _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__xnor2_1
X_1523_ net87 _0632_ _0097_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ seq_div.R\[14\] seq_div.D\[7\] VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1170_ pwm.count\[3\] _0510_ _0331_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0954_ _0321_ _0325_ _0232_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0885_ _0252_ _0258_ _0214_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1506_ _0430_ _0712_ _0086_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__o21ai_1
X_1437_ _0638_ _0736_ _0655_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__a21oi_1
X_1299_ pwm.count\[0\] _0592_ _0610_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or4_1
X_1368_ _0678_ seq_div.R\[22\] _0668_ _0679_ _0672_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput15 keypad_i[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1222_ _0551_ VGND VGND VPWR VPWR clk8.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_1153_ _0502_ VGND VGND VPWR VPWR clk_div.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
X_1084_ osc.count\[0\] osc.count\[1\] osc.count\[2\] VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0799_ net27 _0172_ _0173_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__and3_1
X_0868_ _0206_ _0186_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__nor2_1
X_0937_ _0167_ _0306_ _0308_ _0178_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1771_ clknet_4_0_0_clk net11 net28 VGND VGND VPWR VPWR kp_encoder.q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1205_ net103 _0537_ _0539_ VGND VGND VPWR VPWR clk8.next_count\[4\] sky130_fd_sc_hd__o21a_1
X_1136_ _0331_ _0417_ _0448_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__and4_1
X_1067_ osc.count\[6\] _0373_ _0437_ _0435_ osc.count\[5\] VGND VGND VPWR VPWR _0438_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 kp_encoder.q\[10\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1754_ clknet_4_8_0_clk net48 net33 VGND VGND VPWR VPWR kp_encoder.sync_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1685_ clknet_4_11_0_clk _0041_ net34 VGND VGND VPWR VPWR seq_div.D\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1119_ osc.count\[11\] osc.count\[10\] _0473_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ _0668_ _0764_ _0669_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1668_ clknet_4_13_0_clk _0024_ net36 VGND VGND VPWR VPWR seq_div.q_out\[5\] sky130_fd_sc_hd__dfrtp_1
X_1737_ clknet_4_4_0_clk clk8.next_count\[6\] net29 VGND VGND VPWR VPWR clk8.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1599_ net125 osc.count\[11\] _0132_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0970_ _0340_ _0336_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__nand2_1
X_1453_ _0749_ _0750_ _0658_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a21o_1
X_1522_ _0382_ _0375_ _0391_ _0712_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1384_ seq_div.D\[0\] _0675_ _0695_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0953_ _0284_ _0324_ _0176_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0884_ _0167_ _0254_ _0255_ _0257_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__o31a_1
X_1367_ seq_div.D\[14\] seq_div.R\[21\] VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__and2b_1
X_1505_ net104 _0712_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__nand2_1
X_1436_ net98 _0712_ _0739_ _0625_ _0740_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o221a_1
X_1298_ seq_div.q_out\[1\] _0588_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 keypad_i[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1221_ _0549_ _0531_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__and3b_1
X_1152_ _0500_ _0331_ _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and3b_1
X_1083_ osc.count\[0\] osc.count\[2\] osc.count\[1\] VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0936_ _0165_ _0229_ _0212_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0798_ SS_FSM.count\[4\] SS_FSM.count\[5\] SS_FSM.count\[8\] VGND VGND VPWR VPWR
+ _0173_ sky130_fd_sc_hd__nor3_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0867_ _0159_ _0213_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1419_ net83 _0712_ _0725_ _0625_ _0726_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ clknet_4_2_0_clk net10 net28 VGND VGND VPWR VPWR kp_encoder.q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1204_ clk8.count\[4\] _0537_ _0350_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1135_ osc.count\[15\] _0488_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__xnor2_1
X_1066_ _0375_ _0391_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0919_ _0179_ SS_FSM.count\[2\] _0196_ _0155_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 kp_encoder.q\[13\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1753_ clknet_4_2_0_clk net53 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1684_ clknet_4_10_0_clk _0040_ net34 VGND VGND VPWR VPWR seq_div.D\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1118_ _0478_ VGND VGND VPWR VPWR osc.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
X_1049_ _0382_ _0361_ _0370_ _0351_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__o31a_2
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1736_ clknet_4_4_0_clk clk8.next_count\[5\] net29 VGND VGND VPWR VPWR clk8.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1667_ clknet_4_15_0_clk _0023_ net37 VGND VGND VPWR VPWR seq_div.q_out\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1598_ _0143_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1452_ net91 _0712_ _0717_ seq_div.R\[18\] _0753_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o221a_1
X_1383_ _0642_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1521_ _0096_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1719_ clknet_4_12_0_clk _0075_ net35 VGND VGND VPWR VPWR seq_div.dividend\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0952_ _0230_ _0323_ _0159_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__a21oi_1
X_1504_ seq_div.Q\[6\] _0628_ _0634_ net59 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0883_ _0228_ _0256_ _0159_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__o21a_1
X_1366_ seq_div.D\[15\] VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__inv_2
X_1435_ seq_div.R\[15\] _0717_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1297_ _0582_ _0611_ _0612_ _0591_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
Xinput17 n_rst VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1220_ clk8.count\[9\] _0546_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__or2_1
X_1151_ clk_div.count\[3\] clk_div.count\[4\] _0494_ clk_div.count\[5\] VGND VGND
+ VPWR VPWR _0501_ sky130_fd_sc_hd__a31o_1
X_1082_ _0451_ VGND VGND VPWR VPWR osc.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_0935_ _0179_ _0162_ _0228_ _0183_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0866_ _0154_ _0159_ _0168_ _0239_ _0240_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__a311o_1
X_0797_ SS_FSM.count\[6\] SS_FSM.count\[7\] VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1349_ _0659_ _0660_ _0640_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1418_ seq_div.R\[12\] _0717_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1134_ _0490_ VGND VGND VPWR VPWR osc.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_1203_ net90 _0534_ _0538_ VGND VGND VPWR VPWR clk8.next_count\[3\] sky130_fd_sc_hd__o21a_1
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1065_ osc.count\[4\] _0381_ _0392_ _0435_ osc.count\[5\] VGND VGND VPWR VPWR _0436_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0849_ _0219_ _0222_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__nand3_1
X_0918_ _0249_ _0250_ SS_FSM.count\[5\] _0167_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 kp_encoder.q\[7\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1752_ clknet_4_8_0_clk net49 net28 VGND VGND VPWR VPWR kp_encoder.sync_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1683_ clknet_4_10_0_clk _0039_ net34 VGND VGND VPWR VPWR seq_div.D\[4\] sky130_fd_sc_hd__dfrtp_1
X_1117_ _0476_ _0417_ _0448_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1048_ _0383_ _0381_ _0386_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__nand3_2
XFILLER_0_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1666_ clknet_4_13_0_clk _0022_ net36 VGND VGND VPWR VPWR seq_div.q_out\[3\] sky130_fd_sc_hd__dfrtp_1
X_1735_ clknet_4_4_0_clk clk8.next_count\[4\] net29 VGND VGND VPWR VPWR clk8.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1597_ net91 osc.count\[10\] _0132_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1520_ net118 _0095_ _0632_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_1
X_1451_ seq_div.R\[17\] _0707_ _0751_ _0752_ _0625_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a221o_1
X_1382_ seq_div.R\[8\] seq_div.D\[1\] VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1718_ clknet_4_6_0_clk _0074_ net35 VGND VGND VPWR VPWR seq_div.dividend\[14\] sky130_fd_sc_hd__dfrtp_1
X_1649_ clknet_4_12_0_clk osc.next_count\[10\] net35 VGND VGND VPWR VPWR osc.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0882_ _0155_ _0196_ SS_FSM.count\[2\] _0179_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a211o_1
X_0951_ _0322_ _0250_ _0167_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__o21ai_1
X_1503_ net62 _0628_ _0634_ seq_div.Q\[6\] VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1296_ _0585_ seq_div.q_out\[0\] VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1365_ _0667_ _0675_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__or3b_1
X_1434_ seq_div.R\[14\] _0707_ _0737_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a22o_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ clk_div.count\[5\] clk_div.count\[4\] _0497_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1081_ _0417_ _0448_ _0449_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__and4_1
X_0865_ SS_FSM.sound\[0\] VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0934_ _0165_ _0229_ _0212_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o21ai_1
X_0796_ SS_FSM.count\[7\] _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1417_ _0724_ seq_div.R\[11\] _0707_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1279_ _0585_ seq_div.q_out\[4\] VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__nand2_1
X_1348_ seq_div.D\[8\] seq_div.R\[15\] VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1133_ _0417_ _0448_ _0488_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__and4_1
X_1202_ _0350_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_1064_ _0373_ _0429_ _0379_ _0378_ _0406_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ _0202_ _0289_ _0178_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a21oi_1
X_0779_ SS_FSM.count\[0\] VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
X_0848_ net27 _0172_ _0173_ _0179_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 kp_encoder.q\[6\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1751_ clknet_4_5_0_clk clk8.next_count\[20\] net32 VGND VGND VPWR VPWR clk8.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_1682_ clknet_4_8_0_clk _0038_ net33 VGND VGND VPWR VPWR seq_div.D\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1116_ osc.count\[10\] _0473_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__or2_1
X_1047_ osc.count\[7\] VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1665_ clknet_4_13_0_clk _0021_ net35 VGND VGND VPWR VPWR seq_div.q_out\[2\] sky130_fd_sc_hd__dfrtp_1
X_1734_ clknet_4_4_0_clk clk8.next_count\[3\] net29 VGND VGND VPWR VPWR clk8.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1596_ _0142_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1450_ _0749_ _0750_ _0706_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a21oi_1
X_1381_ _0690_ _0691_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1717_ clknet_4_6_0_clk _0073_ net35 VGND VGND VPWR VPWR seq_div.dividend\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1648_ clknet_4_9_0_clk osc.next_count\[9\] net33 VGND VGND VPWR VPWR osc.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1579_ net126 osc.count\[1\] _0132_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0881_ _0224_ _0198_ _0165_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a21oi_1
X_0950_ _0190_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1502_ net77 _0628_ _0634_ net62 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a22o_1
X_1433_ _0735_ _0736_ _0706_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a21oi_1
X_1295_ _0585_ seq_div.q_out\[0\] VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1364_ seq_div.D\[12\] seq_div.R\[19\] VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1080_ osc.count\[0\] osc.count\[1\] VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0795_ _0169_ net25 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0933_ _0242_ _0246_ _0178_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__o21ai_1
X_0864_ _0175_ _0218_ _0233_ _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__o31a_1
X_1347_ seq_div.D\[9\] _0639_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__or2_1
X_1416_ _0687_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__xor2_1
X_1278_ _0585_ seq_div.q_out\[4\] VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1201_ clk8.count\[3\] _0534_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1132_ osc.count\[14\] _0485_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1063_ _0381_ _0392_ osc.count\[4\] VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0916_ _0195_ _0197_ _0288_ _0167_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0847_ _0179_ _0155_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 kp_encoder.q\[14\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ clknet_4_5_0_clk clk8.next_count\[19\] net32 VGND VGND VPWR VPWR clk8.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1681_ clknet_4_8_0_clk _0037_ net33 VGND VGND VPWR VPWR seq_div.D\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1046_ _0405_ _0414_ _0415_ _0416_ _0400_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o2111a_4
X_1115_ osc.count\[10\] _0473_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1733_ clknet_4_4_0_clk clk8.next_count\[2\] net29 VGND VGND VPWR VPWR clk8.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1664_ clknet_4_13_0_clk _0020_ net35 VGND VGND VPWR VPWR seq_div.q_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_1595_ net88 osc.count\[9\] _0132_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1029_ osc.count\[15\] _0398_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1380_ _0637_ _0660_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__nand2_1
X_1716_ clknet_4_12_0_clk _0072_ net35 VGND VGND VPWR VPWR seq_div.dividend\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _0133_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1647_ clknet_4_9_0_clk osc.next_count\[8\] net33 VGND VGND VPWR VPWR osc.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0880_ _0184_ SS_FSM.count\[5\] _0253_ _0198_ _0224_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__o311a_1
X_1501_ net75 _0628_ _0634_ net77 VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__a22o_1
X_1363_ _0671_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or2_1
X_1432_ _0735_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__or2_1
X_1294_ mode_FSM.mode\[1\] seq_div.q_out\[0\] VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0932_ _0274_ _0298_ _0299_ _0304_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__a22oi_4
XFILLER_0_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0794_ SS_FSM.count\[6\] VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__inv_2
X_0863_ _0175_ _0235_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1346_ seq_div.D\[10\] seq_div.R\[17\] VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__and2b_1
X_1415_ _0648_ _0719_ _0644_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a21oi_1
X_1277_ seq_div.q_out\[6\] _0588_ _0590_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1200_ _0536_ VGND VGND VPWR VPWR clk8.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_1131_ osc.count\[14\] _0485_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__nand2_1
X_1062_ _0428_ _0431_ _0432_ _0423_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0915_ _0189_ _0198_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_1
X_0846_ _0159_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1329_ _0637_ _0638_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold9 kp_encoder.q\[11\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1680_ clknet_4_10_0_clk _0036_ net34 VGND VGND VPWR VPWR seq_div.D\[1\] sky130_fd_sc_hd__dfrtp_1
X_1114_ _0475_ VGND VGND VPWR VPWR osc.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_1045_ _0399_ _0402_ osc.count\[14\] VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0829_ _0178_ _0187_ _0192_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1663_ clknet_4_6_0_clk _0019_ net35 VGND VGND VPWR VPWR seq_div.q_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_1732_ clknet_4_4_0_clk net66 net29 VGND VGND VPWR VPWR clk8.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1594_ _0141_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_1028_ osc.count\[15\] _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1715_ clknet_4_12_0_clk _0071_ net35 VGND VGND VPWR VPWR seq_div.dividend\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1646_ clknet_4_9_0_clk osc.next_count\[7\] net33 VGND VGND VPWR VPWR osc.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ net123 osc.count\[0\] _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1500_ seq_div.Q\[2\] _0628_ _0634_ net75 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__a22o_1
X_1293_ seq_div.q_out\[2\] _0588_ _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__o21ai_1
X_1362_ _0672_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__nand2_1
X_1431_ _0653_ _0731_ _0656_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1629_ clknet_4_10_0_clk _0009_ net34 VGND VGND VPWR VPWR seq_div.R\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0862_ SS_FSM.sound\[0\] _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0931_ _0189_ _0300_ _0301_ _0303_ _0228_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0793_ _0162_ _0165_ _0167_ SS_FSM.sound\[1\] VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o211a_1
X_1276_ _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1414_ _0628_ _0721_ _0722_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a21o_1
X_1345_ _0652_ _0653_ _0654_ _0655_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a311o_1
XFILLER_0_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1130_ _0487_ VGND VGND VPWR VPWR osc.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1061_ osc.count\[3\] _0420_ _0422_ osc.count\[2\] VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0845_ _0219_ _0165_ _0174_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a21o_1
X_0914_ _0214_ _0284_ _0286_ _0232_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1259_ kp_encoder.last_sk kp_encoder.sync_out\[14\] VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2b_1
X_1328_ seq_div.D\[9\] _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1044_ _0388_ _0404_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__nand2_1
X_1113_ _0473_ _0417_ _0448_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__and4b_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0828_ _0194_ _0201_ _0202_ _0159_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1731_ clknet_4_4_0_clk clk8.next_count\[0\] net29 VGND VGND VPWR VPWR clk8.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1662_ clknet_4_6_0_clk clk_div.next_count\[7\] net30 VGND VGND VPWR VPWR clk_div.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1593_ net99 osc.count\[8\] _0132_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__mux2_1
X_1027_ _0382_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold90 seq_div.dividend\[2\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1576_ _0350_ _0507_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__nor2_8
X_1714_ clknet_4_9_0_clk _0070_ net35 VGND VGND VPWR VPWR seq_div.dividend\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1645_ clknet_4_2_0_clk osc.next_count\[6\] net28 VGND VGND VPWR VPWR osc.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1430_ _0697_ _0655_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__nor2_1
X_1292_ _0582_ _0606_ _0607_ _0591_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__a31o_1
X_1361_ seq_div.D\[14\] seq_div.R\[21\] VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1559_ _0240_ _0114_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__or2_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1628_ clknet_4_10_0_clk _0008_ net34 VGND VGND VPWR VPWR seq_div.R\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0861_ SS_FSM.sound\[1\] VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_2
X_0792_ _0166_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0930_ SS_FSM.count\[5\] _0162_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1413_ seq_div.dividend\[3\] _0632_ _0634_ seq_div.R\[11\] VGND VGND VPWR VPWR _0722_
+ sky130_fd_sc_hd__a22o_1
X_1275_ _0581_ _0585_ mode_FSM.mode\[0\] VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__o21ba_2
X_1344_ seq_div.D\[6\] seq_div.R\[13\] VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1060_ osc.count\[1\] _0427_ _0430_ osc.count\[0\] VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0844_ _0160_ _0161_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__nand2_2
X_0913_ _0159_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1258_ net56 _0573_ _0576_ VGND VGND VPWR VPWR clk8.next_count\[20\] sky130_fd_sc_hd__a21oi_1
X_1189_ _0524_ _0525_ _0526_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__and4b_1
X_1327_ seq_div.R\[16\] VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1043_ _0409_ _0412_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__a21oi_1
X_1112_ osc.count\[9\] _0470_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ _0167_ _0194_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1730_ clknet_4_7_0_clk pwm.next_count\[7\] net31 VGND VGND VPWR VPWR pwm.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1661_ clknet_4_6_0_clk clk_div.next_count\[6\] net30 VGND VGND VPWR VPWR clk_div.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1592_ _0140_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1026_ _0351_ _0361_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold91 seq_div.dividend\[13\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 seq_div.D\[5\] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
X_1713_ clknet_4_9_0_clk _0069_ net38 VGND VGND VPWR VPWR seq_div.dividend\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1575_ net116 _0123_ _0131_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__o21a_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1644_ clknet_4_8_0_clk osc.next_count\[5\] net33 VGND VGND VPWR VPWR osc.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ _0373_ _0361_ _0377_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or3_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1360_ seq_div.R\[21\] seq_div.D\[14\] VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1291_ _0585_ seq_div.q_out\[1\] VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1489_ net121 seq_div.q_out\[4\] _0776_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_1
X_1558_ _0219_ net23 _0117_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__or3b_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ clknet_4_10_0_clk _0007_ net34 VGND VGND VPWR VPWR seq_div.R\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0860_ _0219_ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or2_1
X_0791_ SS_FSM.count\[4\] net27 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1412_ _0720_ seq_div.R\[10\] _0707_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux2_1
X_1343_ seq_div.D\[7\] seq_div.R\[14\] VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__and2b_1
X_1274_ _0585_ seq_div.q_out\[5\] _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0989_ _0352_ _0353_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0912_ _0179_ _0193_ _0228_ _0269_ _0209_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__o311a_1
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0843_ _0176_ _0204_ _0208_ _0215_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__o221a_1
X_1326_ seq_div.R\[14\] seq_div.D\[7\] VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or2b_1
X_1257_ net56 _0573_ _0531_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__o21ai_1
X_1188_ clk8.count\[19\] clk8.count\[18\] clk8.count\[17\] VGND VGND VPWR VPWR _0527_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1042_ osc.count\[11\] _0395_ _0411_ osc.count\[10\] VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__a22o_1
X_1111_ osc.count\[9\] osc.count\[8\] _0467_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0826_ _0195_ _0197_ _0200_ _0167_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a31o_1
X_1309_ _0623_ seq_div.state\[0\] VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1660_ clknet_4_6_0_clk clk_div.next_count\[5\] net30 VGND VGND VPWR VPWR clk_div.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1591_ net98 osc.count\[7\] _0132_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux2_1
X_1025_ osc.count\[11\] _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0809_ _0155_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold92 seq_div.dividend\[14\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 seq_div.R\[23\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 seq_div.D\[10\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1643_ clknet_4_8_0_clk osc.next_count\[4\] net33 VGND VGND VPWR VPWR osc.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_1712_ clknet_4_9_0_clk _0068_ net38 VGND VGND VPWR VPWR seq_div.dividend\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _0236_ _0175_ _0120_ _0127_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a211o_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ _0361_ _0377_ _0351_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1290_ _0585_ seq_div.q_out\[1\] VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1626_ clknet_4_10_0_clk _0006_ net34 VGND VGND VPWR VPWR seq_div.R\[11\] sky130_fd_sc_hd__dfrtp_1
X_1488_ _0081_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
X_1557_ SS_FSM.sound\[1\] _0180_ _0181_ _0269_ SS_FSM.sound\[0\] VGND VGND VPWR VPWR
+ _0120_ sky130_fd_sc_hd__o41ai_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0790_ _0163_ _0164_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__nor2_8
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1273_ _0585_ seq_div.q_out\[5\] _0582_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__o21ai_1
X_1411_ _0684_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__xnor2_1
X_1342_ seq_div.R\[12\] seq_div.D\[5\] VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0988_ _0344_ _0346_ _0358_ _0350_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a31o_1
X_1609_ seq_div.state\[0\] _0132_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0842_ _0171_ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__and2_1
X_0911_ _0211_ _0283_ _0178_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1256_ _0575_ VGND VGND VPWR VPWR clk8.next_count\[19\] sky130_fd_sc_hd__clkbuf_1
X_1325_ seq_div.R\[15\] seq_div.D\[8\] VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__or2b_1
X_1187_ clk8.count\[16\] clk8.count\[20\] clk8.count\[14\] clk8.count\[15\] VGND VGND
+ VPWR VPWR _0526_ sky130_fd_sc_hd__and4b_1
XFILLER_0_19_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1110_ _0472_ VGND VGND VPWR VPWR osc.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1041_ osc.count\[9\] _0408_ _0411_ osc.count\[10\] VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0825_ _0198_ _0199_ _0189_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1239_ clk8.count\[15\] _0560_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__and2_1
X_1308_ seq_div.state\[1\] VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1590_ _0139_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1024_ _0390_ _0392_ _0393_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0808_ _0156_ _0180_ _0181_ _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__o31a_2
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold82 seq_div.Q\[0\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 _0775_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 seq_div.dividend\[7\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1642_ clknet_4_8_0_clk osc.next_count\[3\] net33 VGND VGND VPWR VPWR osc.count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_1711_ clknet_4_9_0_clk _0067_ net38 VGND VGND VPWR VPWR seq_div.dividend\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ net112 _0123_ _0127_ _0130_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__o22a_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1007_ _0361_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__nor2_2
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1625_ clknet_4_10_0_clk _0005_ net34 VGND VGND VPWR VPWR seq_div.R\[10\] sky130_fd_sc_hd__dfrtp_1
X_1556_ _0182_ _0117_ _0119_ _0115_ _0155_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a32o_1
X_1487_ net122 seq_div.q_out\[3\] _0776_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410_ _0643_ _0714_ _0645_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1272_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1341_ seq_div.R\[13\] seq_div.D\[6\] VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0987_ _0354_ kp_encoder.sync_out\[10\] _0337_ _0343_ _0357_ VGND VGND VPWR VPWR
+ _0358_ sky130_fd_sc_hd__a311o_1
X_1608_ _0148_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
X_1539_ net115 _0107_ _0631_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0841_ SS_FSM.count\[7\] _0170_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__nand2_1
X_0910_ _0179_ _0165_ _0166_ _0186_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ _0573_ _0331_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__and3b_1
X_1186_ clk8.count\[7\] clk8.count\[6\] clk8.count\[9\] clk8.count\[8\] VGND VGND
+ VPWR VPWR _0525_ sky130_fd_sc_hd__and4b_1
X_1324_ seq_div.R\[17\] seq_div.D\[10\] VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1040_ _0382_ _0375_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0824_ _0160_ _0161_ _0155_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1307_ net61 _0586_ _0622_ _0350_ VGND VGND VPWR VPWR pwm.pwm sky130_fd_sc_hd__a211oi_1
X_1238_ _0562_ VGND VGND VPWR VPWR clk8.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_1169_ pwm.count\[3\] _0510_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1023_ _0370_ _0383_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0807_ SS_FSM.count\[0\] _0155_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold83 seq_div.Q\[4\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 clk8.count\[10\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 seq_div.dividend\[9\] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 seq_div.dividend\[8\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1572_ _0237_ _0217_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1641_ clknet_4_8_0_clk osc.next_count\[2\] net33 VGND VGND VPWR VPWR osc.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1710_ clknet_4_11_0_clk _0066_ net38 VGND VGND VPWR VPWR seq_div.dividend\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ _0352_ _0362_ _0369_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a21o_2
XFILLER_0_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1555_ _0179_ _0115_ _0118_ _0119_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__a22o_1
X_1624_ clknet_4_10_0_clk _0004_ net34 VGND VGND VPWR VPWR seq_div.R\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _0080_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1340_ _0649_ _0650_ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3b_1
X_1271_ mode_FSM.mode\[1\] mode_FSM.mode\[0\] VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0986_ _0355_ _0339_ _0356_ kp_encoder.sync_out\[1\] kp_encoder.sync_out\[0\] VGND
+ VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1469_ _0628_ _0766_ _0767_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a21o_1
X_1607_ seq_div.dividend\[15\] osc.count\[15\] _0132_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__mux2_1
X_1538_ _0385_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0840_ _0209_ _0178_ _0211_ _0213_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__a41o_1
X_1323_ seq_div.R\[18\] seq_div.D\[11\] VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or2b_1
X_1254_ clk8.count\[19\] _0570_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__or2_1
X_1185_ clk8.count\[11\] clk8.count\[10\] clk8.count\[12\] clk8.count\[13\] VGND VGND
+ VPWR VPWR _0524_ sky130_fd_sc_hd__or4b_1
XFILLER_0_46_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0969_ kp_encoder.sync_out\[9\] _0338_ _0332_ _0339_ _0337_ VGND VGND VPWR VPWR _0340_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0823_ SS_FSM.count\[0\] _0184_ SS_FSM.count\[2\] VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__or3_2
X_1306_ pwm.count\[6\] _0593_ _0586_ net67 _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__o221a_1
X_1237_ _0560_ _0531_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__and3b_1
X_1168_ _0512_ VGND VGND VPWR VPWR pwm.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_1099_ osc.count\[6\] _0461_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _0375_ _0381_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0806_ SS_FSM.count\[4\] SS_FSM.count\[5\] SS_FSM.count\[8\] VGND VGND VPWR VPWR
+ _0181_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold40 seq_div.dividend\[6\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 seq_div.Q\[3\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 seq_div.dividend\[14\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _0012_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0011_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1571_ SS_FSM.count\[6\] _0123_ _0127_ _0129_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__o22a_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ clknet_4_8_0_clk osc.next_count\[1\] net33 VGND VGND VPWR VPWR osc.count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ _0375_ _0361_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1769_ clknet_4_8_0_clk net9 net28 VGND VGND VPWR VPWR kp_encoder.q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1485_ seq_div.Q\[2\] seq_div.q_out\[2\] _0776_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1554_ SS_FSM.sound\[0\] _0114_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__and2_1
X_1623_ clknet_4_8_0_clk net69 net34 VGND VGND VPWR VPWR seq_div.R\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

