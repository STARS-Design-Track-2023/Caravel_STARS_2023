// This is the unpowered netlist.
module z23 (clk,
    interrupt_gpio_in,
    memory_wr,
    nrst,
    keypad_input,
    memory_address_out,
    memory_data_in,
    memory_data_out,
    programmable_gpio_in,
    programmable_gpio_out,
    programmable_gpio_wr,
    ss0,
    ss1,
    ss2,
    ss3,
    ss4,
    ss5,
    ss6,
    ss7);
 input clk;
 input interrupt_gpio_in;
 output memory_wr;
 input nrst;
 input [15:0] keypad_input;
 output [15:0] memory_address_out;
 input [7:0] memory_data_in;
 output [7:0] memory_data_out;
 input [7:0] programmable_gpio_in;
 output [7:0] programmable_gpio_out;
 output [7:0] programmable_gpio_wr;
 output [7:0] ss0;
 output [7:0] ss1;
 output [7:0] ss2;
 output [7:0] ss3;
 output [7:0] ss4;
 output [7:0] ss5;
 output [7:0] ss6;
 output [7:0] ss7;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire \alu.Cin ;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \cu.alu_f[1] ;
 wire \cu.alu_f[2] ;
 wire \cu.alu_f[3] ;
 wire \cu.alu_f[4] ;
 wire \cu.alu_f[5] ;
 wire \cu.alu_f[6] ;
 wire \cu.alu_f[7] ;
 wire \cu.id.alu_opcode[0] ;
 wire \cu.id.alu_opcode[1] ;
 wire \cu.id.alu_opcode[3] ;
 wire \cu.id.can_be_interrupted ;
 wire \cu.id.cb_opcode_x[0] ;
 wire \cu.id.cb_opcode_x[1] ;
 wire \cu.id.cb_opcode_y[0] ;
 wire \cu.id.cb_opcode_y[1] ;
 wire \cu.id.cb_opcode_y[2] ;
 wire \cu.id.cb_opcode_z[0] ;
 wire \cu.id.cb_opcode_z[1] ;
 wire \cu.id.cb_opcode_z[2] ;
 wire \cu.id.imm_i[10] ;
 wire \cu.id.imm_i[11] ;
 wire \cu.id.imm_i[12] ;
 wire \cu.id.imm_i[13] ;
 wire \cu.id.imm_i[14] ;
 wire \cu.id.imm_i[15] ;
 wire \cu.id.imm_i[8] ;
 wire \cu.id.imm_i[9] ;
 wire \cu.id.interrupt_requested ;
 wire \cu.id.is_halted ;
 wire \cu.id.is_interrupted ;
 wire \cu.id.opcode[0] ;
 wire \cu.id.opcode[1] ;
 wire \cu.id.opcode[2] ;
 wire \cu.id.opcode[6] ;
 wire \cu.id.opcode[7] ;
 wire \cu.id.starting_int_service ;
 wire \cu.id.state[0] ;
 wire \cu.id.state[1] ;
 wire \cu.id.state[2] ;
 wire \cu.ir.idx[0] ;
 wire \cu.ir.idx[1] ;
 wire \cu.pc.pc_o[0] ;
 wire \cu.pc.pc_o[10] ;
 wire \cu.pc.pc_o[11] ;
 wire \cu.pc.pc_o[12] ;
 wire \cu.pc.pc_o[13] ;
 wire \cu.pc.pc_o[14] ;
 wire \cu.pc.pc_o[15] ;
 wire \cu.pc.pc_o[1] ;
 wire \cu.pc.pc_o[2] ;
 wire \cu.pc.pc_o[3] ;
 wire \cu.pc.pc_o[4] ;
 wire \cu.pc.pc_o[5] ;
 wire \cu.pc.pc_o[6] ;
 wire \cu.pc.pc_o[7] ;
 wire \cu.pc.pc_o[8] ;
 wire \cu.pc.pc_o[9] ;
 wire \cu.reg_file.reg_a[0] ;
 wire \cu.reg_file.reg_a[1] ;
 wire \cu.reg_file.reg_a[2] ;
 wire \cu.reg_file.reg_a[3] ;
 wire \cu.reg_file.reg_a[4] ;
 wire \cu.reg_file.reg_a[5] ;
 wire \cu.reg_file.reg_a[6] ;
 wire \cu.reg_file.reg_a[7] ;
 wire \cu.reg_file.reg_b[0] ;
 wire \cu.reg_file.reg_b[1] ;
 wire \cu.reg_file.reg_b[2] ;
 wire \cu.reg_file.reg_b[3] ;
 wire \cu.reg_file.reg_b[4] ;
 wire \cu.reg_file.reg_b[5] ;
 wire \cu.reg_file.reg_b[6] ;
 wire \cu.reg_file.reg_b[7] ;
 wire \cu.reg_file.reg_c[0] ;
 wire \cu.reg_file.reg_c[1] ;
 wire \cu.reg_file.reg_c[2] ;
 wire \cu.reg_file.reg_c[3] ;
 wire \cu.reg_file.reg_c[4] ;
 wire \cu.reg_file.reg_c[5] ;
 wire \cu.reg_file.reg_c[6] ;
 wire \cu.reg_file.reg_c[7] ;
 wire \cu.reg_file.reg_d[0] ;
 wire \cu.reg_file.reg_d[1] ;
 wire \cu.reg_file.reg_d[2] ;
 wire \cu.reg_file.reg_d[3] ;
 wire \cu.reg_file.reg_d[4] ;
 wire \cu.reg_file.reg_d[5] ;
 wire \cu.reg_file.reg_d[6] ;
 wire \cu.reg_file.reg_d[7] ;
 wire \cu.reg_file.reg_e[0] ;
 wire \cu.reg_file.reg_e[1] ;
 wire \cu.reg_file.reg_e[2] ;
 wire \cu.reg_file.reg_e[3] ;
 wire \cu.reg_file.reg_e[4] ;
 wire \cu.reg_file.reg_e[5] ;
 wire \cu.reg_file.reg_e[6] ;
 wire \cu.reg_file.reg_e[7] ;
 wire \cu.reg_file.reg_h[0] ;
 wire \cu.reg_file.reg_h[1] ;
 wire \cu.reg_file.reg_h[2] ;
 wire \cu.reg_file.reg_h[3] ;
 wire \cu.reg_file.reg_h[4] ;
 wire \cu.reg_file.reg_h[5] ;
 wire \cu.reg_file.reg_h[6] ;
 wire \cu.reg_file.reg_h[7] ;
 wire \cu.reg_file.reg_l[0] ;
 wire \cu.reg_file.reg_l[1] ;
 wire \cu.reg_file.reg_l[2] ;
 wire \cu.reg_file.reg_l[3] ;
 wire \cu.reg_file.reg_l[4] ;
 wire \cu.reg_file.reg_l[5] ;
 wire \cu.reg_file.reg_l[6] ;
 wire \cu.reg_file.reg_l[7] ;
 wire \cu.reg_file.reg_mem[0] ;
 wire \cu.reg_file.reg_mem[10] ;
 wire \cu.reg_file.reg_mem[11] ;
 wire \cu.reg_file.reg_mem[12] ;
 wire \cu.reg_file.reg_mem[13] ;
 wire \cu.reg_file.reg_mem[14] ;
 wire \cu.reg_file.reg_mem[15] ;
 wire \cu.reg_file.reg_mem[1] ;
 wire \cu.reg_file.reg_mem[2] ;
 wire \cu.reg_file.reg_mem[3] ;
 wire \cu.reg_file.reg_mem[4] ;
 wire \cu.reg_file.reg_mem[5] ;
 wire \cu.reg_file.reg_mem[6] ;
 wire \cu.reg_file.reg_mem[7] ;
 wire \cu.reg_file.reg_mem[8] ;
 wire \cu.reg_file.reg_mem[9] ;
 wire \cu.reg_file.reg_sp[0] ;
 wire \cu.reg_file.reg_sp[10] ;
 wire \cu.reg_file.reg_sp[11] ;
 wire \cu.reg_file.reg_sp[12] ;
 wire \cu.reg_file.reg_sp[13] ;
 wire \cu.reg_file.reg_sp[14] ;
 wire \cu.reg_file.reg_sp[15] ;
 wire \cu.reg_file.reg_sp[1] ;
 wire \cu.reg_file.reg_sp[2] ;
 wire \cu.reg_file.reg_sp[3] ;
 wire \cu.reg_file.reg_sp[4] ;
 wire \cu.reg_file.reg_sp[5] ;
 wire \cu.reg_file.reg_sp[6] ;
 wire \cu.reg_file.reg_sp[7] ;
 wire \cu.reg_file.reg_sp[8] ;
 wire \cu.reg_file.reg_sp[9] ;
 wire \ih.gpio_interrupt_mask[0] ;
 wire \ih.gpio_interrupt_mask[1] ;
 wire \ih.gpio_interrupt_mask[2] ;
 wire \ih.gpio_interrupt_mask[3] ;
 wire \ih.gpio_interrupt_mask[4] ;
 wire \ih.gpio_interrupt_mask[5] ;
 wire \ih.gpio_interrupt_mask[6] ;
 wire \ih.gpio_interrupt_mask[7] ;
 wire \ih.ih.ih.prev_data[0] ;
 wire \ih.ih.ih.prev_data[10] ;
 wire \ih.ih.ih.prev_data[11] ;
 wire \ih.ih.ih.prev_data[12] ;
 wire \ih.ih.ih.prev_data[13] ;
 wire \ih.ih.ih.prev_data[14] ;
 wire \ih.ih.ih.prev_data[15] ;
 wire \ih.ih.ih.prev_data[1] ;
 wire \ih.ih.ih.prev_data[2] ;
 wire \ih.ih.ih.prev_data[3] ;
 wire \ih.ih.ih.prev_data[4] ;
 wire \ih.ih.ih.prev_data[5] ;
 wire \ih.ih.ih.prev_data[6] ;
 wire \ih.ih.ih.prev_data[7] ;
 wire \ih.ih.ih.prev_data[8] ;
 wire \ih.ih.ih.prev_data[9] ;
 wire \ih.ih.int_f.data_in ;
 wire \ih.ih.int_f.prev_data ;
 wire \ih.input_handler_enable ;
 wire \ih.interrupt_source[1] ;
 wire \ih.interrupt_source[2] ;
 wire \ih.interrupt_source[3] ;
 wire \ih.ip_ed.prev_data ;
 wire \ih.t.count[0] ;
 wire \ih.t.count[10] ;
 wire \ih.t.count[11] ;
 wire \ih.t.count[12] ;
 wire \ih.t.count[13] ;
 wire \ih.t.count[14] ;
 wire \ih.t.count[15] ;
 wire \ih.t.count[16] ;
 wire \ih.t.count[17] ;
 wire \ih.t.count[18] ;
 wire \ih.t.count[19] ;
 wire \ih.t.count[1] ;
 wire \ih.t.count[20] ;
 wire \ih.t.count[21] ;
 wire \ih.t.count[22] ;
 wire \ih.t.count[23] ;
 wire \ih.t.count[24] ;
 wire \ih.t.count[25] ;
 wire \ih.t.count[26] ;
 wire \ih.t.count[27] ;
 wire \ih.t.count[28] ;
 wire \ih.t.count[29] ;
 wire \ih.t.count[2] ;
 wire \ih.t.count[30] ;
 wire \ih.t.count[31] ;
 wire \ih.t.count[3] ;
 wire \ih.t.count[4] ;
 wire \ih.t.count[5] ;
 wire \ih.t.count[6] ;
 wire \ih.t.count[7] ;
 wire \ih.t.count[8] ;
 wire \ih.t.count[9] ;
 wire \ih.t.enable ;
 wire \ih.t.next_count[0] ;
 wire \ih.t.next_count[10] ;
 wire \ih.t.next_count[11] ;
 wire \ih.t.next_count[12] ;
 wire \ih.t.next_count[13] ;
 wire \ih.t.next_count[14] ;
 wire \ih.t.next_count[15] ;
 wire \ih.t.next_count[16] ;
 wire \ih.t.next_count[17] ;
 wire \ih.t.next_count[18] ;
 wire \ih.t.next_count[19] ;
 wire \ih.t.next_count[1] ;
 wire \ih.t.next_count[20] ;
 wire \ih.t.next_count[21] ;
 wire \ih.t.next_count[22] ;
 wire \ih.t.next_count[23] ;
 wire \ih.t.next_count[24] ;
 wire \ih.t.next_count[25] ;
 wire \ih.t.next_count[26] ;
 wire \ih.t.next_count[27] ;
 wire \ih.t.next_count[28] ;
 wire \ih.t.next_count[29] ;
 wire \ih.t.next_count[2] ;
 wire \ih.t.next_count[30] ;
 wire \ih.t.next_count[31] ;
 wire \ih.t.next_count[3] ;
 wire \ih.t.next_count[4] ;
 wire \ih.t.next_count[5] ;
 wire \ih.t.next_count[6] ;
 wire \ih.t.next_count[7] ;
 wire \ih.t.next_count[8] ;
 wire \ih.t.next_count[9] ;
 wire \ih.t.timer_max[0] ;
 wire \ih.t.timer_max[10] ;
 wire \ih.t.timer_max[11] ;
 wire \ih.t.timer_max[12] ;
 wire \ih.t.timer_max[13] ;
 wire \ih.t.timer_max[14] ;
 wire \ih.t.timer_max[15] ;
 wire \ih.t.timer_max[16] ;
 wire \ih.t.timer_max[17] ;
 wire \ih.t.timer_max[18] ;
 wire \ih.t.timer_max[19] ;
 wire \ih.t.timer_max[1] ;
 wire \ih.t.timer_max[20] ;
 wire \ih.t.timer_max[21] ;
 wire \ih.t.timer_max[22] ;
 wire \ih.t.timer_max[23] ;
 wire \ih.t.timer_max[24] ;
 wire \ih.t.timer_max[25] ;
 wire \ih.t.timer_max[26] ;
 wire \ih.t.timer_max[27] ;
 wire \ih.t.timer_max[28] ;
 wire \ih.t.timer_max[29] ;
 wire \ih.t.timer_max[2] ;
 wire \ih.t.timer_max[30] ;
 wire \ih.t.timer_max[31] ;
 wire \ih.t.timer_max[3] ;
 wire \ih.t.timer_max[4] ;
 wire \ih.t.timer_max[5] ;
 wire \ih.t.timer_max[6] ;
 wire \ih.t.timer_max[7] ;
 wire \ih.t.timer_max[8] ;
 wire \ih.t.timer_max[9] ;
 wire \mc.cc.count[0] ;
 wire \mc.cc.count[1] ;
 wire \mc.cc.count[2] ;
 wire \mc.cc.count[3] ;
 wire \mc.cc.enable ;
 wire \mc.cc.enable_edge_detector.prev_data ;
 wire \mc.cl.cmp_o ;
 wire \mc.cl.next_data[0] ;
 wire \mc.cl.next_data[10] ;
 wire \mc.cl.next_data[11] ;
 wire \mc.cl.next_data[12] ;
 wire \mc.cl.next_data[13] ;
 wire \mc.cl.next_data[14] ;
 wire \mc.cl.next_data[15] ;
 wire \mc.cl.next_data[1] ;
 wire \mc.cl.next_data[2] ;
 wire \mc.cl.next_data[3] ;
 wire \mc.cl.next_data[4] ;
 wire \mc.cl.next_data[5] ;
 wire \mc.cl.next_data[6] ;
 wire \mc.cl.next_data[7] ;
 wire \mc.cl.next_data[8] ;
 wire \mc.cl.next_data[9] ;
 wire \mc.count ;
 wire \mc.rw.next_state[0] ;
 wire \mc.rw.next_state[1] ;
 wire \mc.rw.next_state[2] ;
 wire \mc.rw.state[0] ;
 wire \mc.rw.state[1] ;
 wire \mc.rw.state[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(programmable_gpio_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(programmable_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(keypad_input[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2972__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__A_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__A_N (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A_N (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__A_N (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A (.DIODE(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__B (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__C (.DIODE(\ih.t.timer_max[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__B (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__A (.DIODE(\ih.t.timer_max[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__A (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__B (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A (.DIODE(\ih.t.timer_max[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__B (.DIODE(\ih.t.timer_max[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__B1 (.DIODE(\ih.t.timer_max[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A1 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A (.DIODE(\ih.t.timer_max[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A1 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__B1 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__A (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__A (.DIODE(\ih.t.timer_max[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__B1 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__S (.DIODE(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A1 (.DIODE(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A2 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__B1 (.DIODE(\ih.t.timer_max[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__B_N (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__C (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A2 (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A1 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__B (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A1 (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__B (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__B1 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__B1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__C1 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__A (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__D_N (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__C (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A2 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__C1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__B (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A2 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__B1_N (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A1_N (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__D1 (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__B (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__B (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__B (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__B (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__B (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__B (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__B1 (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A1 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__B1 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__B (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__B1 (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__C1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A1 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__A (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__B (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__B1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__B1 (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__B2 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__B1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__B1 (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A_N (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__D (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__B (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__C (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A1 (.DIODE(\cu.reg_file.reg_sp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__B2 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__B (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__C_N (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__B1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__B_N (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__B1 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A_N (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__B (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__B1_N (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__B2 (.DIODE(\cu.reg_file.reg_e[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__A_N (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__A (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__B (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__B2 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A1 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A1 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__B2 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__B (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A1 (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A1 (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__B1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A2 (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__C1 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__B1 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__C1 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__B2 (.DIODE(\cu.reg_file.reg_e[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A1 (.DIODE(\cu.reg_file.reg_sp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B1 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A1 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A2 (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A1 (.DIODE(\cu.pc.pc_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A2 (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B2 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__B2 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A1 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__C1 (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__C1 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__C1 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A1 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__B2 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__A1 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__D1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A1 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B1 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A1 (.DIODE(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__B1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__B_N (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__C1 (.DIODE(\cu.reg_file.reg_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__B1 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A1 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A2 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__B2 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A1 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A2 (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A1 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__B2 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__B2 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A1 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A1 (.DIODE(\cu.reg_file.reg_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__B2 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__B1 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A1 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A1 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__B2 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A1 (.DIODE(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B2 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A1 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__B2 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__C (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A0 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A1 (.DIODE(\cu.reg_file.reg_c[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__B2 (.DIODE(\cu.alu_f[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A1 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A2 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B2 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A1 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A2 (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__C1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__B1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__B2 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A1 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A1 (.DIODE(\cu.reg_file.reg_c[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__D1 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A1_N (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__C_N (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B2 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A1 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__B2 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__B2 (.DIODE(\cu.reg_file.reg_a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A1 (.DIODE(\cu.reg_file.reg_l[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__D1 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1_N (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__B2 (.DIODE(\cu.reg_file.reg_a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A1 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A1 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B1 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__C1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__B2 (.DIODE(\cu.reg_file.reg_l[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__C_N (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A1 (.DIODE(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__B2 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A1 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A1 (.DIODE(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B2 (.DIODE(\cu.reg_file.reg_a[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__D1 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A1_N (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A0 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A1 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A2 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__B2 (.DIODE(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A1 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A2 (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__B2 (.DIODE(\cu.reg_file.reg_a[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A1 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B1 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B2 (.DIODE(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__C1 (.DIODE(\cu.reg_file.reg_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A1 (.DIODE(\cu.reg_file.reg_c[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__B2 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A1 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A2 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__B2 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__B2 (.DIODE(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A1 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A2 (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__B2 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__C1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A1 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B1 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B2 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__B1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A1 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__B2 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A1 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A1 (.DIODE(\cu.reg_file.reg_c[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__B2 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A1 (.DIODE(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__B2 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(\cu.reg_file.reg_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A1_N (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__C1 (.DIODE(\cu.reg_file.reg_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__B2 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A1 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A2 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__B2 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A1 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A2 (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__C1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A1 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B1 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A2 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__B (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__B (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__B (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A1 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__B2 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A1 (.DIODE(\cu.reg_file.reg_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A1_N (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__C (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A1 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__B2 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A1 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A1 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A1 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B2 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__D (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A_N (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__B (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__B (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A1_N (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__B2 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__B2 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A1 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A1 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__B2 (.DIODE(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A1 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A1 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A1 (.DIODE(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__B2 (.DIODE(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A1 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A1 (.DIODE(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__B2 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__B2 (.DIODE(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A1 (.DIODE(\cu.reg_file.reg_a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__B2 (.DIODE(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__B2 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A1 (.DIODE(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A1 (.DIODE(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B2 (.DIODE(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A1 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A1 (.DIODE(\cu.reg_file.reg_a[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B2 (.DIODE(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A1 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A1 (.DIODE(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B2 (.DIODE(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A1 (.DIODE(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B2 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A1 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A1 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B2 (.DIODE(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A1 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A1 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__B2 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A1 (.DIODE(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B2 (.DIODE(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A1 (.DIODE(\cu.pc.pc_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A1 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A1 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A1 (.DIODE(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B2 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A1 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A1 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A1 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A1 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B_N (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B_N (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1_N (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2_N (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A_N (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__B1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A2 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A2 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B2 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A1 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A1 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__B2 (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__C1 (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B2 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__D (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A1 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B1 (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A1 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__D (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A_N (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A1 (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(_2918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__C_N (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__B1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A2 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B2 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__C1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A2 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B2 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__B (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A1_N (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B2 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A1_N (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A2_N (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A2 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__B1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A2_N (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__B1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__B (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__B2 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__B (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__B (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__B (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__B2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__B1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A2 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__B2 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A2 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__B2 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A2 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B2 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__B1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__B1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__C (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__B1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A1_N (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A3 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A3 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__B2 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__C (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__C (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__C (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__D (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__B (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__S (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A0 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A1 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__S (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__S (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A0 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__S (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__S (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A0 (.DIODE(\cu.alu_f[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A1 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__S (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A2 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__B1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__B2 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A2 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__C_N (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__A1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__B1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A1 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__B2 (.DIODE(\cu.reg_file.reg_sp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A1 (.DIODE(\cu.reg_file.reg_e[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__B2 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__C (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__A (.DIODE(\cu.pc.pc_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A1 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__B2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__B (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__C (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__B_N (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__C (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__D_N (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A1 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A2 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A1 (.DIODE(\cu.reg_file.reg_sp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(\cu.reg_file.reg_e[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__B2 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__C1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A1 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__B2 (.DIODE(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A1 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__B2 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A1 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__B2 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A1 (.DIODE(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B2 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A1 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__B2 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__B2 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A1 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B2 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A1 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__B2 (.DIODE(\cu.reg_file.reg_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__B2 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A1 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__B2 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__C1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A1 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__B2 (.DIODE(\cu.reg_file.reg_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A2 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__C1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A2 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__B1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A2 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__B2 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__B (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A1 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__B2 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A1 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__B2 (.DIODE(\cu.reg_file.reg_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A1 (.DIODE(\cu.reg_file.reg_c[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A1 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__B2 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A (.DIODE(\cu.reg_file.reg_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A1 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__B2 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A1 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B2 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(\cu.reg_file.reg_c[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__A2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A_N (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A1 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A1 (.DIODE(\cu.reg_file.reg_a[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__B2 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A1 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__B2 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A1 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__B2 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__C1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A1 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__C (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__B (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__B (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A1 (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A1 (.DIODE(\cu.reg_file.reg_a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__B2 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__A1 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__B2 (.DIODE(\cu.reg_file.reg_l[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B2 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A (.DIODE(\cu.reg_file.reg_l[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__B2 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__C1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B2 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__B (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__B (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__B (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A2 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B1_N (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A2 (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__B2 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A1 (.DIODE(\cu.reg_file.reg_c[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B2 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A1 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B2 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A1 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(\cu.reg_file.reg_c[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__B (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__B (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A1 (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A1 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__B2 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__B2 (.DIODE(\cu.reg_file.reg_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A1 (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B2 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A (.DIODE(\cu.reg_file.reg_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__B2 (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A1 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A3 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__B (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A1 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B2 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__B1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__B (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A1 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B2 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__C1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A2 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A1 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B2 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__C1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A2 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B2 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A1 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__B2 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A1 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A1 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__B2 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A1 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B2 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A1 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B (.DIODE(_1511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__B (.DIODE(_1511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A2 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__B (.DIODE(_1511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__B2 (.DIODE(_1511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A (.DIODE(\cu.pc.pc_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__B2 (.DIODE(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A1 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__B2 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__C1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A2 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A1 (.DIODE(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__B2 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A2 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A1 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A1 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__B2 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A1 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A1 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__B2 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__C1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__A2 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A1 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B2 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A2 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__B2 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A1 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B2 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__B (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__B (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A2 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__B (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__B (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A1 (.DIODE(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__B2 (.DIODE(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__B1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A1 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__B2 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A1 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A2 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A1 (.DIODE(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__B1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__B2 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__C1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A1 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A2 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B2 (.DIODE(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A1 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B2 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B (.DIODE(_1561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A2 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__C (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B (.DIODE(_1561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__B (.DIODE(_1561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A2_N (.DIODE(_1561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__B2 (.DIODE(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__B1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__B2 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A2 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A1 (.DIODE(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__B1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__C1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A2 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B2 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A1 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__B2 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A1 (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A2 (.DIODE(_1561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A2 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A (.DIODE(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A1 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__B2 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__C1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A2 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A1 (.DIODE(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__B2 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__B2 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__B2 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__B (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__B (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__B (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A2_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__B2 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__B1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A1 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__B2 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__C1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A1 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A1 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A2 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A1 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B2 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__C1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A1 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A2 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__C_N (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A2 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__B1 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A2 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__B1 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__B1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A2 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B1 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A2 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A2 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B1 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A2 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__B1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A2 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A (.DIODE(_1561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__C (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A (.DIODE(_1511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__C (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__D_N (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__C (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__C1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__C (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A2 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B1 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A1 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A2 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A0 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A1 (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A2 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__B2 (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__B (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__C (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__C (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__C (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__C (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__C (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__C (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__C (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A2 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__B1 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A0 (.DIODE(\cu.alu_f[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__B1 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B2 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A2 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A3 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A2 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A3 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A2 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__C (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__B (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A2 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A0 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A1_N (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A1 (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__C1 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A1 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A2 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A2 (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A0 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__B (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__B (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A0 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__B (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__C (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A2 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B1 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__B (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A2 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A0 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A0 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__B (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__B (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A0 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A0 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__B (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A0 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A0 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__B1 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__B (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__B (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A0 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A0 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__B (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A0 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A0 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__B (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__B (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A0 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A1 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__B1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__B (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__B (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__B1 (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A0 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__B (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A0 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A0 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__B (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A1 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A2 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__B1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__S (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A0 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__S (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__S (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A0 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__S (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A0 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A2 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__B1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__B1 (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__S (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A0 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__S (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A0 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__S (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A0 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__B1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B1_N (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__S (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A0 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__S (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__B1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A0 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A0 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__S (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A1 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A0 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A0 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A1 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A0 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A0 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A0 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A1 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A0 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A0 (.DIODE(\cu.reg_file.reg_a[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A1 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A0 (.DIODE(\cu.reg_file.reg_a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A0 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__S (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A1 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A1 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B1 (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A0 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A0 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A1 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A0 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A0 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A1 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A0 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A0 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A0 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A0 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__S (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B1 (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A0 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A0 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A1 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A0 (.DIODE(\cu.reg_file.reg_c[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A0 (.DIODE(\cu.reg_file.reg_c[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A0 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__S (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A0 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A1 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A1 (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B1 (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A0 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A0 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A1 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A0 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A0 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A0 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A0 (.DIODE(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A0 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A0 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__S (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__S (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(_2035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__B1 (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A0 (.DIODE(\cu.reg_file.reg_e[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A0 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A0 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A1 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A0 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A0 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__B1_N (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A1 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A0 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A1 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A1 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A0 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A1 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A0 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A1 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A1 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A0 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__S (.DIODE(_2066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__S (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A0 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A0 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A0 (.DIODE(\cu.reg_file.reg_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A0 (.DIODE(\cu.reg_file.reg_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A1 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A0 (.DIODE(\cu.reg_file.reg_l[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A0 (.DIODE(\cu.reg_file.reg_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__C_N (.DIODE(_2951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A0 (.DIODE(\cu.reg_file.reg_sp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__C (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A0 (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A0 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__S (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__S (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A0 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__S (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A0 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__S (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A0 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__S (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A0 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A1 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__S (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A0 (.DIODE(\ih.t.timer_max[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(_2163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A0 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__S (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__S (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A1 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__S (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__S (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__S (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__S (.DIODE(_2206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__S (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__S (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__S (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A0 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A0 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A0 (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__C (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__B (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A3 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__S0 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__S1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A0 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A1 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A2 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B2 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A1_N (.DIODE(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A1 (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__C1 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__C1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__D1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__C (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__S0 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__S1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__B2 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__C (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A1 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A1 (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__S (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__B2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__B1 (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A1 (.DIODE(\ih.t.timer_max[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B2 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A_N (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B2 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__C1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A2 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__C (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(_2372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__S (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A2 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B1 (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A1 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B2 (.DIODE(\ih.t.timer_max[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A_N (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B2 (.DIODE(\ih.t.timer_max[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__C1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__B2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A1 (.DIODE(_2391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__S (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A2 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B1 (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A1 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A_N (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__C1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A0 (.DIODE(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__S (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A2 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__B2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__B1 (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A1 (.DIODE(\ih.t.timer_max[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A_N (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__C1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A0 (.DIODE(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__S (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A2 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__B1 (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B2 (.DIODE(_2435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A1 (.DIODE(\ih.t.timer_max[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A_N (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__C1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A1 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__S (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__B1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B1 (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A_N (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__C1 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A1 (.DIODE(_2467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__B2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B1 (.DIODE(_2225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A2 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__B2 (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A_N (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__C1 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B2 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__C (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B2 (.DIODE(\ih.t.timer_max[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B2 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B2 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__B1 (.DIODE(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__B2 (.DIODE(\ih.t.timer_max[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__B1 (.DIODE(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A1 (.DIODE(\ih.t.timer_max[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__B2 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__B1 (.DIODE(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__B2 (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A2_N (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__B1 (.DIODE(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__B2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__B (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__C1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A1 (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A2 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A (.DIODE(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A1 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A2 (.DIODE(_2532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B1 (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__B1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A0 (.DIODE(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A0 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A0 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A1 (.DIODE(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A0 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A0 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A0 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A0 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A0 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A0 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A0 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A0 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A0 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A0 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A0 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A0 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A (.DIODE(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A (.DIODE(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A0 (.DIODE(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A0 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A (.DIODE(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A (.DIODE(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A0 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A0 (.DIODE(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A (.DIODE(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A (.DIODE(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A0 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A0 (.DIODE(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A (.DIODE(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A0 (.DIODE(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A (.DIODE(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A0 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A0 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A1 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A1 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A0 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A1 (.DIODE(\ih.t.timer_max[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A0 (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A1 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A1 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(\ih.t.timer_max[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A0 (.DIODE(_2163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A1 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A1 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A0 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A1 (.DIODE(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A0 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A0 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(\ih.t.timer_max[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__S (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A1 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A2 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A1 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A2 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__B1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A1 (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A2 (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A3 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A2 (.DIODE(_2532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A0 (.DIODE(_2923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A1 (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A1 (.DIODE(_2372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A1 (.DIODE(_2391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A0 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A0 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A1 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A0 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A1 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A1 (.DIODE(_2467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A0 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A1 (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A0 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A1 (.DIODE(_2372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A0 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A1 (.DIODE(_2391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A0 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A0 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A0 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A1 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A0 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1 (.DIODE(_2467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A0 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__S (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A0 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A0 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A1 (.DIODE(_2372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A0 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A1 (.DIODE(_2391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A0 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A0 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A1 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__A1 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A0 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A1 (.DIODE(_2467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A0 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__RESET_B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__RESET_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__RESET_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__RESET_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__RESET_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__SET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__RESET_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__RESET_B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__RESET_B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__RESET_B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__RESET_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__RESET_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__RESET_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__RESET_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__RESET_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__RESET_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__RESET_B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__RESET_B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__D (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__D (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__D (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__RESET_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__RESET_B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__RESET_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_85 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _2954_ (.A(\mc.rw.state[1] ),
    .Y(_2695_));
 sky130_fd_sc_hd__and3_1 _2955_ (.A(\mc.rw.state[2] ),
    .B(_2695_),
    .C(\mc.rw.state[0] ),
    .X(_2696_));
 sky130_fd_sc_hd__clkbuf_8 _2956_ (.A(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__inv_2 _2957_ (.A(\mc.rw.state[2] ),
    .Y(_2698_));
 sky130_fd_sc_hd__nor2_2 _2958_ (.A(_2695_),
    .B(\mc.rw.state[0] ),
    .Y(_2699_));
 sky130_fd_sc_hd__and3b_1 _2959_ (.A_N(\mc.rw.state[0] ),
    .B(\mc.rw.state[2] ),
    .C(_2695_),
    .X(_2700_));
 sky130_fd_sc_hd__clkbuf_4 _2960_ (.A(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__a21o_4 _2961_ (.A1(_2698_),
    .A2(_2699_),
    .B1(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__or2_1 _2962_ (.A(_2697_),
    .B(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__clkbuf_1 _2963_ (.A(_2703_),
    .X(net59));
 sky130_fd_sc_hd__and2_1 _2964_ (.A(_2695_),
    .B(\mc.rw.state[0] ),
    .X(_2704_));
 sky130_fd_sc_hd__nor2_1 _2965_ (.A(_2704_),
    .B(_2699_),
    .Y(_2705_));
 sky130_fd_sc_hd__and3_1 _2966_ (.A(_2698_),
    .B(\mc.rw.state[1] ),
    .C(\mc.rw.state[0] ),
    .X(_2706_));
 sky130_fd_sc_hd__nor2_1 _2967_ (.A(_2701_),
    .B(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__and2_2 _2968_ (.A(_2705_),
    .B(_2707_),
    .X(_2708_));
 sky130_fd_sc_hd__inv_2 _2969_ (.A(_2708_),
    .Y(\mc.cc.enable ));
 sky130_fd_sc_hd__inv_2 _2970_ (.A(net9),
    .Y(_2709_));
 sky130_fd_sc_hd__inv_2 _2971_ (.A(net4),
    .Y(_2710_));
 sky130_fd_sc_hd__inv_2 _2972_ (.A(net10),
    .Y(_2711_));
 sky130_fd_sc_hd__inv_2 _2973_ (.A(net11),
    .Y(_2712_));
 sky130_fd_sc_hd__o22a_1 _2974_ (.A1(_2711_),
    .A2(\ih.ih.ih.prev_data[2] ),
    .B1(_2712_),
    .B2(\ih.ih.ih.prev_data[3] ),
    .X(_2713_));
 sky130_fd_sc_hd__o221a_1 _2975_ (.A1(_2709_),
    .A2(\ih.ih.ih.prev_data[1] ),
    .B1(_2710_),
    .B2(net233),
    .C1(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__inv_2 _2976_ (.A(net14),
    .Y(_2715_));
 sky130_fd_sc_hd__inv_2 _2977_ (.A(net5),
    .Y(_2716_));
 sky130_fd_sc_hd__inv_2 _2978_ (.A(net12),
    .Y(_2717_));
 sky130_fd_sc_hd__inv_2 _2979_ (.A(net6),
    .Y(_2718_));
 sky130_fd_sc_hd__o22a_1 _2980_ (.A1(_2717_),
    .A2(\ih.ih.ih.prev_data[4] ),
    .B1(_2718_),
    .B2(\ih.ih.ih.prev_data[13] ),
    .X(_2719_));
 sky130_fd_sc_hd__o221a_1 _2981_ (.A1(_2715_),
    .A2(\ih.ih.ih.prev_data[6] ),
    .B1(_2716_),
    .B2(\ih.ih.ih.prev_data[12] ),
    .C1(_2719_),
    .X(_2720_));
 sky130_fd_sc_hd__inv_2 _2982_ (.A(net17),
    .Y(_2721_));
 sky130_fd_sc_hd__inv_2 _2983_ (.A(net7),
    .Y(_2722_));
 sky130_fd_sc_hd__inv_2 _2984_ (.A(net13),
    .Y(_2723_));
 sky130_fd_sc_hd__inv_2 _2985_ (.A(net3),
    .Y(_2724_));
 sky130_fd_sc_hd__o22a_1 _2986_ (.A1(_2723_),
    .A2(\ih.ih.ih.prev_data[5] ),
    .B1(_2724_),
    .B2(\ih.ih.ih.prev_data[10] ),
    .X(_2725_));
 sky130_fd_sc_hd__o221a_1 _2987_ (.A1(_2721_),
    .A2(\ih.ih.ih.prev_data[9] ),
    .B1(_2722_),
    .B2(\ih.ih.ih.prev_data[14] ),
    .C1(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__inv_2 _2988_ (.A(net2),
    .Y(_2727_));
 sky130_fd_sc_hd__inv_2 _2989_ (.A(net8),
    .Y(_2728_));
 sky130_fd_sc_hd__inv_2 _2990_ (.A(net15),
    .Y(_2729_));
 sky130_fd_sc_hd__inv_2 _2991_ (.A(net16),
    .Y(_2730_));
 sky130_fd_sc_hd__o22a_1 _2992_ (.A1(_2729_),
    .A2(\ih.ih.ih.prev_data[7] ),
    .B1(_2730_),
    .B2(\ih.ih.ih.prev_data[8] ),
    .X(_2731_));
 sky130_fd_sc_hd__o221a_1 _2993_ (.A1(_2727_),
    .A2(\ih.ih.ih.prev_data[0] ),
    .B1(_2728_),
    .B2(\ih.ih.ih.prev_data[15] ),
    .C1(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__and3_1 _2994_ (.A(_2720_),
    .B(_2726_),
    .C(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__nand2_1 _2995_ (.A(_2714_),
    .B(_2733_),
    .Y(\ih.ih.int_f.data_in ));
 sky130_fd_sc_hd__inv_2 _2996_ (.A(net69),
    .Y(_2734_));
 sky130_fd_sc_hd__and3b_1 _2997_ (.A_N(net68),
    .B(net27),
    .C(\ih.gpio_interrupt_mask[0] ),
    .X(_2735_));
 sky130_fd_sc_hd__a31o_1 _2998_ (.A1(_2734_),
    .A2(net28),
    .A3(\ih.gpio_interrupt_mask[1] ),
    .B1(_2735_),
    .X(_2736_));
 sky130_fd_sc_hd__and3b_1 _2999_ (.A_N(net70),
    .B(net29),
    .C(\ih.gpio_interrupt_mask[2] ),
    .X(_2737_));
 sky130_fd_sc_hd__and3b_1 _3000_ (.A_N(net71),
    .B(net30),
    .C(\ih.gpio_interrupt_mask[3] ),
    .X(_2738_));
 sky130_fd_sc_hd__inv_2 _3001_ (.A(net74),
    .Y(_2739_));
 sky130_fd_sc_hd__inv_2 _3002_ (.A(net73),
    .Y(_2740_));
 sky130_fd_sc_hd__and3b_1 _3003_ (.A_N(net72),
    .B(net31),
    .C(\ih.gpio_interrupt_mask[4] ),
    .X(_2741_));
 sky130_fd_sc_hd__a31o_1 _3004_ (.A1(_2740_),
    .A2(net32),
    .A3(\ih.gpio_interrupt_mask[5] ),
    .B1(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__and3b_1 _3005_ (.A_N(net75),
    .B(net34),
    .C(\ih.gpio_interrupt_mask[7] ),
    .X(_2743_));
 sky130_fd_sc_hd__a311o_1 _3006_ (.A1(_2739_),
    .A2(net33),
    .A3(\ih.gpio_interrupt_mask[6] ),
    .B1(_2742_),
    .C1(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__or4_4 _3007_ (.A(_2736_),
    .B(_2737_),
    .C(_2738_),
    .D(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__or3_1 _3008_ (.A(\ih.t.timer_max[0] ),
    .B(\ih.t.timer_max[1] ),
    .C(\ih.t.timer_max[2] ),
    .X(_2746_));
 sky130_fd_sc_hd__or2_1 _3009_ (.A(\ih.t.timer_max[3] ),
    .B(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__or2_1 _3010_ (.A(\ih.t.timer_max[4] ),
    .B(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3011_ (.A(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__or3_2 _3012_ (.A(\ih.t.timer_max[5] ),
    .B(\ih.t.timer_max[6] ),
    .C(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__or3_1 _3013_ (.A(\ih.t.timer_max[7] ),
    .B(\ih.t.timer_max[8] ),
    .C(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__or2_2 _3014_ (.A(\ih.t.timer_max[9] ),
    .B(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__or3_1 _3015_ (.A(\ih.t.timer_max[10] ),
    .B(\ih.t.timer_max[11] ),
    .C(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__or2_2 _3016_ (.A(\ih.t.timer_max[12] ),
    .B(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__or3_1 _3017_ (.A(\ih.t.timer_max[13] ),
    .B(\ih.t.timer_max[14] ),
    .C(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__or2_2 _3018_ (.A(\ih.t.timer_max[15] ),
    .B(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__or3_1 _3019_ (.A(\ih.t.timer_max[16] ),
    .B(\ih.t.timer_max[17] ),
    .C(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__or2_2 _3020_ (.A(\ih.t.timer_max[18] ),
    .B(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__or3_1 _3021_ (.A(\ih.t.timer_max[19] ),
    .B(\ih.t.timer_max[20] ),
    .C(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__or2_2 _3022_ (.A(\ih.t.timer_max[21] ),
    .B(_2759_),
    .X(_2760_));
 sky130_fd_sc_hd__or3_2 _3023_ (.A(\ih.t.timer_max[22] ),
    .B(\ih.t.timer_max[23] ),
    .C(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__or2_2 _3024_ (.A(\ih.t.timer_max[24] ),
    .B(_2761_),
    .X(_2762_));
 sky130_fd_sc_hd__or3_1 _3025_ (.A(\ih.t.timer_max[25] ),
    .B(\ih.t.timer_max[26] ),
    .C(_2762_),
    .X(_2763_));
 sky130_fd_sc_hd__or2_2 _3026_ (.A(\ih.t.timer_max[27] ),
    .B(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__or3_1 _3027_ (.A(\ih.t.timer_max[28] ),
    .B(\ih.t.timer_max[29] ),
    .C(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__nor2_1 _3028_ (.A(\ih.t.timer_max[30] ),
    .B(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__xnor2_1 _3029_ (.A(\ih.t.count[31] ),
    .B(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__xnor2_1 _3030_ (.A(\ih.t.timer_max[31] ),
    .B(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__o21ai_1 _3031_ (.A1(\ih.t.timer_max[28] ),
    .A2(_2764_),
    .B1(\ih.t.timer_max[29] ),
    .Y(_2769_));
 sky130_fd_sc_hd__and3_1 _3032_ (.A(\ih.t.count[29] ),
    .B(_2765_),
    .C(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__a21oi_1 _3033_ (.A1(_2765_),
    .A2(_2769_),
    .B1(\ih.t.count[29] ),
    .Y(_2771_));
 sky130_fd_sc_hd__xor2_1 _3034_ (.A(\ih.t.timer_max[28] ),
    .B(_2764_),
    .X(_2772_));
 sky130_fd_sc_hd__xnor2_1 _3035_ (.A(\ih.t.count[28] ),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__nand2_1 _3036_ (.A(\ih.t.timer_max[27] ),
    .B(_2763_),
    .Y(_2774_));
 sky130_fd_sc_hd__a21oi_1 _3037_ (.A1(_2764_),
    .A2(_2774_),
    .B1(\ih.t.count[27] ),
    .Y(_2775_));
 sky130_fd_sc_hd__and3_1 _3038_ (.A(\ih.t.count[27] ),
    .B(_2764_),
    .C(_2774_),
    .X(_2776_));
 sky130_fd_sc_hd__o21ai_1 _3039_ (.A1(\ih.t.timer_max[25] ),
    .A2(_2762_),
    .B1(\ih.t.timer_max[26] ),
    .Y(_2777_));
 sky130_fd_sc_hd__and3_1 _3040_ (.A(\ih.t.count[26] ),
    .B(_2763_),
    .C(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__a21oi_1 _3041_ (.A1(_2763_),
    .A2(_2777_),
    .B1(\ih.t.count[26] ),
    .Y(_2779_));
 sky130_fd_sc_hd__xor2_1 _3042_ (.A(\ih.t.timer_max[25] ),
    .B(_2762_),
    .X(_2780_));
 sky130_fd_sc_hd__xnor2_1 _3043_ (.A(\ih.t.count[25] ),
    .B(_2780_),
    .Y(_2781_));
 sky130_fd_sc_hd__nand2_1 _3044_ (.A(\ih.t.timer_max[24] ),
    .B(_2761_),
    .Y(_2782_));
 sky130_fd_sc_hd__and3_1 _3045_ (.A(\ih.t.count[24] ),
    .B(_2762_),
    .C(_2782_),
    .X(_2783_));
 sky130_fd_sc_hd__a21oi_1 _3046_ (.A1(_2762_),
    .A2(_2782_),
    .B1(\ih.t.count[24] ),
    .Y(_2784_));
 sky130_fd_sc_hd__o21ai_1 _3047_ (.A1(\ih.t.timer_max[22] ),
    .A2(_2760_),
    .B1(\ih.t.timer_max[23] ),
    .Y(_2785_));
 sky130_fd_sc_hd__and3_1 _3048_ (.A(\ih.t.count[23] ),
    .B(_2761_),
    .C(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__a21oi_1 _3049_ (.A1(_2761_),
    .A2(_2785_),
    .B1(\ih.t.count[23] ),
    .Y(_2787_));
 sky130_fd_sc_hd__xor2_1 _3050_ (.A(\ih.t.timer_max[22] ),
    .B(_2760_),
    .X(_2788_));
 sky130_fd_sc_hd__xnor2_1 _3051_ (.A(\ih.t.count[22] ),
    .B(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__nand2_1 _3052_ (.A(\ih.t.timer_max[21] ),
    .B(_2759_),
    .Y(_2790_));
 sky130_fd_sc_hd__and3_1 _3053_ (.A(\ih.t.count[21] ),
    .B(_2760_),
    .C(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__a21oi_1 _3054_ (.A1(_2760_),
    .A2(_2790_),
    .B1(\ih.t.count[21] ),
    .Y(_2792_));
 sky130_fd_sc_hd__o21ai_1 _3055_ (.A1(\ih.t.timer_max[19] ),
    .A2(_2758_),
    .B1(\ih.t.timer_max[20] ),
    .Y(_2793_));
 sky130_fd_sc_hd__a21oi_1 _3056_ (.A1(_2759_),
    .A2(_2793_),
    .B1(\ih.t.count[20] ),
    .Y(_2794_));
 sky130_fd_sc_hd__and3_1 _3057_ (.A(\ih.t.count[20] ),
    .B(_2759_),
    .C(_2793_),
    .X(_2795_));
 sky130_fd_sc_hd__xor2_1 _3058_ (.A(\ih.t.timer_max[19] ),
    .B(_2758_),
    .X(_2796_));
 sky130_fd_sc_hd__xnor2_1 _3059_ (.A(\ih.t.count[19] ),
    .B(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__nand2_1 _3060_ (.A(\ih.t.timer_max[18] ),
    .B(_2757_),
    .Y(_2798_));
 sky130_fd_sc_hd__a21oi_1 _3061_ (.A1(_2758_),
    .A2(_2798_),
    .B1(\ih.t.count[18] ),
    .Y(_2799_));
 sky130_fd_sc_hd__and3_1 _3062_ (.A(\ih.t.count[18] ),
    .B(_2758_),
    .C(_2798_),
    .X(_2800_));
 sky130_fd_sc_hd__o21ai_1 _3063_ (.A1(\ih.t.timer_max[16] ),
    .A2(_2756_),
    .B1(\ih.t.timer_max[17] ),
    .Y(_2801_));
 sky130_fd_sc_hd__a21oi_1 _3064_ (.A1(_2757_),
    .A2(_2801_),
    .B1(\ih.t.count[17] ),
    .Y(_2802_));
 sky130_fd_sc_hd__and3_1 _3065_ (.A(\ih.t.count[17] ),
    .B(_2757_),
    .C(_2801_),
    .X(_2803_));
 sky130_fd_sc_hd__xor2_1 _3066_ (.A(\ih.t.timer_max[16] ),
    .B(_2756_),
    .X(_2804_));
 sky130_fd_sc_hd__xnor2_1 _3067_ (.A(\ih.t.count[16] ),
    .B(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__nand2_1 _3068_ (.A(\ih.t.timer_max[15] ),
    .B(_2755_),
    .Y(_2806_));
 sky130_fd_sc_hd__a21oi_1 _3069_ (.A1(_2756_),
    .A2(_2806_),
    .B1(\ih.t.count[15] ),
    .Y(_2807_));
 sky130_fd_sc_hd__and3_1 _3070_ (.A(\ih.t.count[15] ),
    .B(_2756_),
    .C(_2806_),
    .X(_2808_));
 sky130_fd_sc_hd__o21ai_1 _3071_ (.A1(\ih.t.timer_max[13] ),
    .A2(_2754_),
    .B1(\ih.t.timer_max[14] ),
    .Y(_2809_));
 sky130_fd_sc_hd__and3_1 _3072_ (.A(\ih.t.count[14] ),
    .B(_2755_),
    .C(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__a21oi_1 _3073_ (.A1(_2755_),
    .A2(_2809_),
    .B1(\ih.t.count[14] ),
    .Y(_2811_));
 sky130_fd_sc_hd__xor2_1 _3074_ (.A(\ih.t.timer_max[13] ),
    .B(_2754_),
    .X(_2812_));
 sky130_fd_sc_hd__xnor2_1 _3075_ (.A(\ih.t.count[13] ),
    .B(_2812_),
    .Y(_2813_));
 sky130_fd_sc_hd__nand2_1 _3076_ (.A(\ih.t.timer_max[12] ),
    .B(_2753_),
    .Y(_2814_));
 sky130_fd_sc_hd__and3_1 _3077_ (.A(\ih.t.count[12] ),
    .B(_2754_),
    .C(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__a21oi_1 _3078_ (.A1(_2754_),
    .A2(_2814_),
    .B1(\ih.t.count[12] ),
    .Y(_2816_));
 sky130_fd_sc_hd__o21ai_1 _3079_ (.A1(\ih.t.timer_max[10] ),
    .A2(_2752_),
    .B1(\ih.t.timer_max[11] ),
    .Y(_2817_));
 sky130_fd_sc_hd__a21oi_1 _3080_ (.A1(_2753_),
    .A2(_2817_),
    .B1(\ih.t.count[11] ),
    .Y(_2818_));
 sky130_fd_sc_hd__and3_1 _3081_ (.A(\ih.t.count[11] ),
    .B(_2753_),
    .C(_2817_),
    .X(_2819_));
 sky130_fd_sc_hd__xor2_1 _3082_ (.A(\ih.t.timer_max[10] ),
    .B(_2752_),
    .X(_2820_));
 sky130_fd_sc_hd__xnor2_1 _3083_ (.A(\ih.t.count[10] ),
    .B(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__nand2_1 _3084_ (.A(\ih.t.timer_max[9] ),
    .B(_2751_),
    .Y(_2822_));
 sky130_fd_sc_hd__and3_1 _3085_ (.A(\ih.t.count[9] ),
    .B(_2752_),
    .C(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__a21oi_1 _3086_ (.A1(_2752_),
    .A2(_2822_),
    .B1(\ih.t.count[9] ),
    .Y(_2824_));
 sky130_fd_sc_hd__o21ai_1 _3087_ (.A1(\ih.t.timer_max[7] ),
    .A2(_2750_),
    .B1(\ih.t.timer_max[8] ),
    .Y(_2825_));
 sky130_fd_sc_hd__and3_1 _3088_ (.A(\ih.t.count[8] ),
    .B(_2751_),
    .C(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__a21oi_1 _3089_ (.A1(_2751_),
    .A2(_2825_),
    .B1(\ih.t.count[8] ),
    .Y(_2827_));
 sky130_fd_sc_hd__xor2_1 _3090_ (.A(\ih.t.timer_max[7] ),
    .B(_2750_),
    .X(_2828_));
 sky130_fd_sc_hd__xnor2_1 _3091_ (.A(\ih.t.count[7] ),
    .B(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__o21ai_1 _3092_ (.A1(\ih.t.timer_max[5] ),
    .A2(_2749_),
    .B1(\ih.t.timer_max[6] ),
    .Y(_2830_));
 sky130_fd_sc_hd__and3_1 _3093_ (.A(\ih.t.count[6] ),
    .B(_2750_),
    .C(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__a21oi_1 _3094_ (.A1(_2750_),
    .A2(_2830_),
    .B1(\ih.t.count[6] ),
    .Y(_2832_));
 sky130_fd_sc_hd__xor2_1 _3095_ (.A(\ih.t.timer_max[5] ),
    .B(_2749_),
    .X(_2833_));
 sky130_fd_sc_hd__xnor2_1 _3096_ (.A(\ih.t.count[5] ),
    .B(_2833_),
    .Y(_2834_));
 sky130_fd_sc_hd__nand2_1 _3097_ (.A(\ih.t.timer_max[4] ),
    .B(_2747_),
    .Y(_2835_));
 sky130_fd_sc_hd__xnor2_1 _3098_ (.A(\ih.t.timer_max[1] ),
    .B(\ih.t.count[1] ),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_1 _3099_ (.A(\ih.t.count[0] ),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(_2836_),
    .A1(\ih.t.count[0] ),
    .S(\ih.t.timer_max[0] ),
    .X(_2838_));
 sky130_fd_sc_hd__o21ai_1 _3101_ (.A1(\ih.t.timer_max[0] ),
    .A2(\ih.t.timer_max[1] ),
    .B1(\ih.t.timer_max[2] ),
    .Y(_2839_));
 sky130_fd_sc_hd__and3_1 _3102_ (.A(\ih.t.count[2] ),
    .B(_2746_),
    .C(_2839_),
    .X(_2840_));
 sky130_fd_sc_hd__a21oi_1 _3103_ (.A1(_2746_),
    .A2(_2839_),
    .B1(\ih.t.count[2] ),
    .Y(_2841_));
 sky130_fd_sc_hd__or4_1 _3104_ (.A(_2837_),
    .B(_2838_),
    .C(_2840_),
    .D(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__a31o_1 _3105_ (.A1(\ih.t.count[4] ),
    .A2(_2749_),
    .A3(_2835_),
    .B1(_2842_),
    .X(_2843_));
 sky130_fd_sc_hd__a21oi_1 _3106_ (.A1(_2749_),
    .A2(_2835_),
    .B1(\ih.t.count[4] ),
    .Y(_2844_));
 sky130_fd_sc_hd__nand2_1 _3107_ (.A(\ih.t.timer_max[3] ),
    .B(_2746_),
    .Y(_2845_));
 sky130_fd_sc_hd__nand2_1 _3108_ (.A(_2747_),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__xor2_1 _3109_ (.A(\ih.t.count[3] ),
    .B(_2846_),
    .X(_2847_));
 sky130_fd_sc_hd__or4_1 _3110_ (.A(_2834_),
    .B(_2843_),
    .C(_2844_),
    .D(_2847_),
    .X(_2848_));
 sky130_fd_sc_hd__or4_1 _3111_ (.A(_2829_),
    .B(_2831_),
    .C(_2832_),
    .D(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__or3_1 _3112_ (.A(_2826_),
    .B(_2827_),
    .C(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__or4_1 _3113_ (.A(_2821_),
    .B(_2823_),
    .C(_2824_),
    .D(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__or3_1 _3114_ (.A(_2818_),
    .B(_2819_),
    .C(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__or4_1 _3115_ (.A(_2813_),
    .B(_2815_),
    .C(_2816_),
    .D(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__or3_1 _3116_ (.A(_2810_),
    .B(_2811_),
    .C(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__or4_1 _3117_ (.A(_2805_),
    .B(_2807_),
    .C(_2808_),
    .D(_2854_),
    .X(_2855_));
 sky130_fd_sc_hd__or3_1 _3118_ (.A(_2802_),
    .B(_2803_),
    .C(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__or4_1 _3119_ (.A(_2797_),
    .B(_2799_),
    .C(_2800_),
    .D(_2856_),
    .X(_2857_));
 sky130_fd_sc_hd__or3_1 _3120_ (.A(_2794_),
    .B(_2795_),
    .C(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__or4_1 _3121_ (.A(_2789_),
    .B(_2791_),
    .C(_2792_),
    .D(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__or3_1 _3122_ (.A(_2786_),
    .B(_2787_),
    .C(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__or4_1 _3123_ (.A(_2781_),
    .B(_2783_),
    .C(_2784_),
    .D(_2860_),
    .X(_2861_));
 sky130_fd_sc_hd__or3_1 _3124_ (.A(_2778_),
    .B(_2779_),
    .C(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__or4_1 _3125_ (.A(_2773_),
    .B(_2775_),
    .C(_2776_),
    .D(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__or3_1 _3126_ (.A(_2770_),
    .B(_2771_),
    .C(_2863_),
    .X(_2864_));
 sky130_fd_sc_hd__and2_1 _3127_ (.A(\ih.t.timer_max[30] ),
    .B(_2765_),
    .X(_2865_));
 sky130_fd_sc_hd__nor2_1 _3128_ (.A(_2766_),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__nor2_1 _3129_ (.A(\ih.t.count[30] ),
    .B(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__nand2_1 _3130_ (.A(\ih.t.count[30] ),
    .B(_2866_),
    .Y(_2868_));
 sky130_fd_sc_hd__or4b_4 _3131_ (.A(_2768_),
    .B(_2864_),
    .C(_2867_),
    .D_N(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__and3b_4 _3132_ (.A_N(\ih.ih.int_f.prev_data ),
    .B(\ih.ih.int_f.data_in ),
    .C(\ih.input_handler_enable ),
    .X(_2870_));
 sky130_fd_sc_hd__inv_2 _3133_ (.A(_2870_),
    .Y(_2871_));
 sky130_fd_sc_hd__or2b_1 _3134_ (.A(_2745_),
    .B_N(_2869_),
    .X(_2872_));
 sky130_fd_sc_hd__nor3_1 _3135_ (.A(net1),
    .B(_2872_),
    .C(_2870_),
    .Y(_2873_));
 sky130_fd_sc_hd__a32o_1 _3136_ (.A1(_2745_),
    .A2(_2869_),
    .A3(_2871_),
    .B1(net140),
    .B2(net202),
    .X(_0000_));
 sky130_fd_sc_hd__and3_2 _3137_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[0] ),
    .C(\cu.id.alu_opcode[3] ),
    .X(_2874_));
 sky130_fd_sc_hd__clkbuf_4 _3138_ (.A(\cu.id.opcode[6] ),
    .X(_2875_));
 sky130_fd_sc_hd__clkbuf_4 _3139_ (.A(\cu.id.opcode[7] ),
    .X(_2876_));
 sky130_fd_sc_hd__nand2b_4 _3140_ (.A_N(_2875_),
    .B(_2876_),
    .Y(_2877_));
 sky130_fd_sc_hd__nand3b_4 _3141_ (.A_N(\cu.id.opcode[0] ),
    .B(\cu.id.opcode[2] ),
    .C(\cu.id.opcode[1] ),
    .Y(_2878_));
 sky130_fd_sc_hd__nand2_1 _3142_ (.A(_2875_),
    .B(_2876_),
    .Y(_2879_));
 sky130_fd_sc_hd__or2_2 _3143_ (.A(_2878_),
    .B(_2879_),
    .X(_2880_));
 sky130_fd_sc_hd__and2_1 _3144_ (.A(_2877_),
    .B(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__nor2_1 _3145_ (.A(_2874_),
    .B(_2881_),
    .Y(_2882_));
 sky130_fd_sc_hd__inv_2 _3146_ (.A(\cu.id.alu_opcode[1] ),
    .Y(_2883_));
 sky130_fd_sc_hd__clkbuf_4 _3147_ (.A(\cu.id.alu_opcode[3] ),
    .X(_2884_));
 sky130_fd_sc_hd__and2_2 _3148_ (.A(\cu.id.alu_opcode[0] ),
    .B(\cu.id.opcode[0] ),
    .X(_2885_));
 sky130_fd_sc_hd__and4bb_1 _3149_ (.A_N(\cu.id.opcode[6] ),
    .B_N(\cu.id.opcode[7] ),
    .C(\cu.id.opcode[2] ),
    .D(\cu.id.opcode[1] ),
    .X(_2886_));
 sky130_fd_sc_hd__and4_2 _3150_ (.A(_2883_),
    .B(_2884_),
    .C(_2885_),
    .D(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__nor2_2 _3151_ (.A(_2875_),
    .B(_2876_),
    .Y(_2888_));
 sky130_fd_sc_hd__and3_1 _3152_ (.A(\cu.id.opcode[0] ),
    .B(\cu.id.opcode[2] ),
    .C(\cu.id.opcode[1] ),
    .X(_2889_));
 sky130_fd_sc_hd__and2b_1 _3153_ (.A_N(\cu.id.alu_opcode[3] ),
    .B(\cu.id.alu_opcode[1] ),
    .X(_2890_));
 sky130_fd_sc_hd__and3_1 _3154_ (.A(_2888_),
    .B(_2889_),
    .C(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__clkbuf_4 _3155_ (.A(\cu.id.alu_opcode[0] ),
    .X(_2892_));
 sky130_fd_sc_hd__clkbuf_4 _3156_ (.A(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__buf_4 _3157_ (.A(\cu.id.opcode[0] ),
    .X(_2894_));
 sky130_fd_sc_hd__nor4b_1 _3158_ (.A(\cu.id.opcode[2] ),
    .B(\cu.id.opcode[6] ),
    .C(\cu.id.opcode[7] ),
    .D_N(\cu.id.opcode[1] ),
    .Y(_2895_));
 sky130_fd_sc_hd__nand2_4 _3159_ (.A(_2894_),
    .B(net243),
    .Y(_2896_));
 sky130_fd_sc_hd__inv_2 _3160_ (.A(_2894_),
    .Y(_2897_));
 sky130_fd_sc_hd__nand2_1 _3161_ (.A(_2893_),
    .B(_2897_),
    .Y(_2898_));
 sky130_fd_sc_hd__buf_2 _3162_ (.A(\cu.id.opcode[2] ),
    .X(_2899_));
 sky130_fd_sc_hd__buf_2 _3163_ (.A(\cu.id.opcode[1] ),
    .X(_2900_));
 sky130_fd_sc_hd__or4b_4 _3164_ (.A(_2899_),
    .B(_2875_),
    .C(_2876_),
    .D_N(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__buf_4 _3165_ (.A(\cu.id.alu_opcode[1] ),
    .X(_2902_));
 sky130_fd_sc_hd__or3b_2 _3166_ (.A(_2901_),
    .B(_2902_),
    .C_N(_2884_),
    .X(_2903_));
 sky130_fd_sc_hd__or2_2 _3167_ (.A(_2898_),
    .B(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__o21ai_1 _3168_ (.A1(_2893_),
    .A2(_2896_),
    .B1(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__or3_1 _3169_ (.A(_2887_),
    .B(_2891_),
    .C(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__and3b_1 _3170_ (.A_N(\cu.id.alu_opcode[0] ),
    .B(\cu.id.alu_opcode[3] ),
    .C(\cu.id.alu_opcode[1] ),
    .X(_2907_));
 sky130_fd_sc_hd__and2b_2 _3171_ (.A_N(\cu.id.opcode[7] ),
    .B(\cu.id.opcode[6] ),
    .X(_2908_));
 sky130_fd_sc_hd__or2_1 _3172_ (.A(\cu.id.opcode[6] ),
    .B(\cu.id.opcode[7] ),
    .X(_2909_));
 sky130_fd_sc_hd__or2b_1 _3173_ (.A(_2900_),
    .B_N(_2899_),
    .X(_2910_));
 sky130_fd_sc_hd__or2_1 _3174_ (.A(_2909_),
    .B(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__clkbuf_4 _3175_ (.A(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__or2_2 _3176_ (.A(_2909_),
    .B(_2878_),
    .X(_2913_));
 sky130_fd_sc_hd__nand2_2 _3177_ (.A(_2912_),
    .B(_2913_),
    .Y(_2914_));
 sky130_fd_sc_hd__nor2_1 _3178_ (.A(_2908_),
    .B(_2914_),
    .Y(_2915_));
 sky130_fd_sc_hd__or4bb_4 _3179_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[3] ),
    .C_N(\cu.id.opcode[0] ),
    .D_N(\cu.id.alu_opcode[0] ),
    .X(_2916_));
 sky130_fd_sc_hd__and4b_2 _3180_ (.A_N(_2899_),
    .B(_2900_),
    .C(_2875_),
    .D(_2876_),
    .X(_2917_));
 sky130_fd_sc_hd__nand2b_4 _3181_ (.A_N(_2916_),
    .B(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__and3b_1 _3182_ (.A_N(\cu.id.cb_opcode_z[0] ),
    .B(\cu.id.cb_opcode_z[1] ),
    .C(\cu.id.cb_opcode_z[2] ),
    .X(_2919_));
 sky130_fd_sc_hd__buf_4 _3183_ (.A(\cu.id.cb_opcode_x[1] ),
    .X(_2920_));
 sky130_fd_sc_hd__inv_2 _3184_ (.A(\cu.id.cb_opcode_x[0] ),
    .Y(_2921_));
 sky130_fd_sc_hd__nor2_1 _3185_ (.A(_2920_),
    .B(_2921_),
    .Y(_2922_));
 sky130_fd_sc_hd__clkbuf_4 _3186_ (.A(_2894_),
    .X(_2923_));
 sky130_fd_sc_hd__or3b_2 _3187_ (.A(_2901_),
    .B(_2923_),
    .C_N(_2874_),
    .X(_2924_));
 sky130_fd_sc_hd__nand2_4 _3188_ (.A(_2892_),
    .B(_2894_),
    .Y(_2925_));
 sky130_fd_sc_hd__nor2_1 _3189_ (.A(_2925_),
    .B(_2901_),
    .Y(_2926_));
 sky130_fd_sc_hd__nor2_1 _3190_ (.A(_2902_),
    .B(\cu.id.alu_opcode[3] ),
    .Y(_2927_));
 sky130_fd_sc_hd__and3_1 _3191_ (.A(_2888_),
    .B(_2889_),
    .C(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__nor2_1 _3192_ (.A(_2926_),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__o311a_1 _3193_ (.A1(_2918_),
    .A2(_2919_),
    .A3(_2922_),
    .B1(_2924_),
    .C1(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__or4_1 _3194_ (.A(\cu.id.opcode[2] ),
    .B(\cu.id.opcode[1] ),
    .C(\cu.id.opcode[6] ),
    .D(\cu.id.opcode[7] ),
    .X(_2931_));
 sky130_fd_sc_hd__buf_2 _3195_ (.A(_2931_),
    .X(_2932_));
 sky130_fd_sc_hd__nor2_2 _3196_ (.A(_2899_),
    .B(_2900_),
    .Y(_2933_));
 sky130_fd_sc_hd__nor2_2 _3197_ (.A(\cu.id.alu_opcode[0] ),
    .B(\cu.id.opcode[0] ),
    .Y(_2934_));
 sky130_fd_sc_hd__nand4_4 _3198_ (.A(_2888_),
    .B(_2890_),
    .C(_2933_),
    .D(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__clkbuf_4 _3199_ (.A(_2884_),
    .X(_2936_));
 sky130_fd_sc_hd__or3_2 _3200_ (.A(_2936_),
    .B(_2901_),
    .C(_2898_),
    .X(_2937_));
 sky130_fd_sc_hd__or2b_1 _3201_ (.A(\cu.id.alu_opcode[0] ),
    .B_N(_2894_),
    .X(_2938_));
 sky130_fd_sc_hd__or4bb_4 _3202_ (.A(_2899_),
    .B(\cu.id.opcode[1] ),
    .C_N(_2875_),
    .D_N(_2876_),
    .X(_2939_));
 sky130_fd_sc_hd__nor2_2 _3203_ (.A(_2938_),
    .B(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__and4bb_2 _3204_ (.A_N(\cu.id.opcode[2] ),
    .B_N(\cu.id.opcode[1] ),
    .C(_2875_),
    .D(_2876_),
    .X(_2941_));
 sky130_fd_sc_hd__and4_1 _3205_ (.A(_2902_),
    .B(_2936_),
    .C(_2885_),
    .D(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__nor2_1 _3206_ (.A(_2940_),
    .B(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__o2111a_1 _3207_ (.A1(_2897_),
    .A2(_2932_),
    .B1(_2935_),
    .C1(_2937_),
    .D1(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__o211ai_1 _3208_ (.A1(_2907_),
    .A2(_2915_),
    .B1(_2930_),
    .C1(_2944_),
    .Y(_2945_));
 sky130_fd_sc_hd__inv_2 _3209_ (.A(\cu.id.state[2] ),
    .Y(_2946_));
 sky130_fd_sc_hd__nand2_2 _3210_ (.A(\cu.id.state[1] ),
    .B(\cu.id.state[0] ),
    .Y(_2947_));
 sky130_fd_sc_hd__nor2_8 _3211_ (.A(_2946_),
    .B(_2947_),
    .Y(_2948_));
 sky130_fd_sc_hd__inv_2 _3212_ (.A(\cu.id.starting_int_service ),
    .Y(_2949_));
 sky130_fd_sc_hd__buf_4 _3213_ (.A(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__o311a_4 _3214_ (.A1(_2882_),
    .A2(_2906_),
    .A3(_2945_),
    .B1(_2948_),
    .C1(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__or2_2 _3215_ (.A(_2938_),
    .B(_2932_),
    .X(_2952_));
 sky130_fd_sc_hd__nand2_2 _3216_ (.A(_2896_),
    .B(_2952_),
    .Y(_2953_));
 sky130_fd_sc_hd__clkbuf_4 _3217_ (.A(\cu.id.starting_int_service ),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_4 _3218_ (.A(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_4 _3219_ (.A(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_4 _3220_ (.A(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__o21ai_1 _3221_ (.A1(_2925_),
    .A2(_2932_),
    .B1(_2904_),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _3222_ (.A(_2892_),
    .Y(_0298_));
 sky130_fd_sc_hd__and2_1 _3223_ (.A(_2902_),
    .B(_2884_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _3224_ (.A(_0298_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2b_4 _3225_ (.A_N(_2876_),
    .B(_2875_),
    .Y(_0301_));
 sky130_fd_sc_hd__nor2_1 _3226_ (.A(_0300_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__and3b_1 _3227_ (.A_N(_2916_),
    .B(_2917_),
    .C(_2919_),
    .X(_0303_));
 sky130_fd_sc_hd__nand3_2 _3228_ (.A(_2936_),
    .B(_2885_),
    .C(_2941_),
    .Y(_0304_));
 sky130_fd_sc_hd__or4bb_1 _3229_ (.A(_2902_),
    .B(_2884_),
    .C_N(_2875_),
    .D_N(_2876_),
    .X(_0305_));
 sky130_fd_sc_hd__or4bb_1 _3230_ (.A(_2892_),
    .B(_2899_),
    .C_N(_2900_),
    .D_N(_2923_),
    .X(_0306_));
 sky130_fd_sc_hd__o2bb2a_2 _3231_ (.A1_N(_2897_),
    .A2_N(_2917_),
    .B1(_0305_),
    .B2(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__o21ai_2 _3232_ (.A1(_2902_),
    .A2(_0304_),
    .B1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__and4b_1 _3233_ (.A_N(\cu.id.opcode[1] ),
    .B(\cu.id.opcode[6] ),
    .C(\cu.id.opcode[7] ),
    .D(\cu.id.opcode[2] ),
    .X(_0309_));
 sky130_fd_sc_hd__and3_1 _3234_ (.A(_2923_),
    .B(_2874_),
    .C(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__and3_1 _3235_ (.A(_2885_),
    .B(_2927_),
    .C(_0309_),
    .X(_0311_));
 sky130_fd_sc_hd__a21oi_4 _3236_ (.A1(_2894_),
    .A2(_2916_),
    .B1(_2939_),
    .Y(_0312_));
 sky130_fd_sc_hd__or2_2 _3237_ (.A(_2892_),
    .B(\cu.id.opcode[0] ),
    .X(_0313_));
 sky130_fd_sc_hd__or3_1 _3238_ (.A(_2910_),
    .B(_0313_),
    .C(_0305_),
    .X(_0314_));
 sky130_fd_sc_hd__or4b_4 _3239_ (.A(_0310_),
    .B(_0311_),
    .C(_0312_),
    .D_N(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__nor2_1 _3240_ (.A(_0308_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _3241_ (.A(_2943_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nor2_1 _3242_ (.A(_2938_),
    .B(_2931_),
    .Y(_0318_));
 sky130_fd_sc_hd__o211a_1 _3243_ (.A1(_2892_),
    .A2(_2884_),
    .B1(net151),
    .C1(_2897_),
    .X(_0319_));
 sky130_fd_sc_hd__and3b_2 _3244_ (.A_N(_2884_),
    .B(net151),
    .C(_2934_),
    .X(_0320_));
 sky130_fd_sc_hd__or4b_4 _3245_ (.A(_0318_),
    .B(_0319_),
    .C(_0320_),
    .D_N(_2913_),
    .X(_0321_));
 sky130_fd_sc_hd__nand3_2 _3246_ (.A(_2896_),
    .B(_2911_),
    .C(_2935_),
    .Y(_0322_));
 sky130_fd_sc_hd__and3b_1 _3247_ (.A_N(_2878_),
    .B(_2907_),
    .C(_2908_),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_2 _3248_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[3] ),
    .Y(_0324_));
 sky130_fd_sc_hd__or2_1 _3249_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[3] ),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_1 _3250_ (.A(_2899_),
    .B(_2900_),
    .Y(_0326_));
 sky130_fd_sc_hd__a2111o_1 _3251_ (.A1(_0324_),
    .A2(_0325_),
    .B1(_2897_),
    .C1(_2909_),
    .D1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__or4b_2 _3252_ (.A(_2887_),
    .B(_2891_),
    .C(_0323_),
    .D_N(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__nor2_1 _3253_ (.A(_2925_),
    .B(_2932_),
    .Y(_0329_));
 sky130_fd_sc_hd__or2b_1 _3254_ (.A(_2894_),
    .B_N(_2884_),
    .X(_0330_));
 sky130_fd_sc_hd__or4bb_1 _3255_ (.A(\cu.id.opcode[0] ),
    .B(\cu.id.alu_opcode[3] ),
    .C_N(\cu.id.alu_opcode[1] ),
    .D_N(_2892_),
    .X(_0331_));
 sky130_fd_sc_hd__a21oi_1 _3256_ (.A1(_0330_),
    .A2(_0331_),
    .B1(_2932_),
    .Y(_0332_));
 sky130_fd_sc_hd__and4_1 _3257_ (.A(_2888_),
    .B(_2927_),
    .C(_2933_),
    .D(_2934_),
    .X(_0333_));
 sky130_fd_sc_hd__or3_1 _3258_ (.A(_0329_),
    .B(_0332_),
    .C(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__nor4_1 _3259_ (.A(_0321_),
    .B(_0322_),
    .C(_0328_),
    .D(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__buf_2 _3260_ (.A(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__o31a_1 _3261_ (.A1(_0302_),
    .A2(_0303_),
    .A3(_0317_),
    .B1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _3262_ (.A(_2907_),
    .B(_2914_),
    .X(_0338_));
 sky130_fd_sc_hd__or4_2 _3263_ (.A(_0296_),
    .B(_0297_),
    .C(_0337_),
    .D(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__buf_4 _3264_ (.A(\cu.id.cb_opcode_z[1] ),
    .X(_0340_));
 sky130_fd_sc_hd__buf_4 _3265_ (.A(\cu.id.cb_opcode_z[2] ),
    .X(_0341_));
 sky130_fd_sc_hd__and3_1 _3266_ (.A(_2885_),
    .B(_2927_),
    .C(_2917_),
    .X(_0342_));
 sky130_fd_sc_hd__buf_4 _3267_ (.A(\cu.id.cb_opcode_z[0] ),
    .X(_0343_));
 sky130_fd_sc_hd__nand3_1 _3268_ (.A(_0343_),
    .B(\cu.id.cb_opcode_z[1] ),
    .C(\cu.id.cb_opcode_z[2] ),
    .Y(_0344_));
 sky130_fd_sc_hd__o211a_1 _3269_ (.A1(_0340_),
    .A2(_0341_),
    .B1(_0342_),
    .C1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _3270_ (.A(_2874_),
    .B(_2927_),
    .X(_0346_));
 sky130_fd_sc_hd__o21ai_1 _3271_ (.A1(_0301_),
    .A2(_0346_),
    .B1(_0316_),
    .Y(_0347_));
 sky130_fd_sc_hd__o31a_1 _3272_ (.A1(_2942_),
    .A2(_0345_),
    .A3(_0347_),
    .B1(_0336_),
    .X(_0348_));
 sky130_fd_sc_hd__nor2_1 _3273_ (.A(_2874_),
    .B(_2927_),
    .Y(_0349_));
 sky130_fd_sc_hd__clkbuf_4 _3274_ (.A(_0296_),
    .X(_0350_));
 sky130_fd_sc_hd__a221o_1 _3275_ (.A1(_0299_),
    .A2(_2953_),
    .B1(_0349_),
    .B2(_2914_),
    .C1(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_2 _3276_ (.A(_0348_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _3277_ (.A(_2892_),
    .B(_0324_),
    .Y(_0353_));
 sky130_fd_sc_hd__or2_1 _3278_ (.A(_2883_),
    .B(_2936_),
    .X(_0354_));
 sky130_fd_sc_hd__a21bo_1 _3279_ (.A1(_0340_),
    .A2(_0341_),
    .B1_N(_0343_),
    .X(_0355_));
 sky130_fd_sc_hd__a2bb2o_1 _3280_ (.A1_N(_2918_),
    .A2_N(_0355_),
    .B1(_2883_),
    .B2(_2940_),
    .X(_0356_));
 sky130_fd_sc_hd__a2111o_1 _3281_ (.A1(_0354_),
    .A2(_2953_),
    .B1(_0297_),
    .C1(_0356_),
    .D1(_2942_),
    .X(_0357_));
 sky130_fd_sc_hd__o21ba_1 _3282_ (.A1(_2915_),
    .A2(_0353_),
    .B1_N(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_4 _3283_ (.A(_2902_),
    .X(_0359_));
 sky130_fd_sc_hd__inv_2 _3284_ (.A(_0340_),
    .Y(_0360_));
 sky130_fd_sc_hd__clkbuf_4 _3285_ (.A(_0342_),
    .X(_0361_));
 sky130_fd_sc_hd__and4_1 _3286_ (.A(_2888_),
    .B(_2890_),
    .C(_2933_),
    .D(_2934_),
    .X(_0362_));
 sky130_fd_sc_hd__a2111oi_1 _3287_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0362_),
    .C1(_0297_),
    .D1(_0296_),
    .Y(_0363_));
 sky130_fd_sc_hd__xnor2_4 _3288_ (.A(_2902_),
    .B(_2884_),
    .Y(_0364_));
 sky130_fd_sc_hd__o21bai_1 _3289_ (.A1(_2940_),
    .A2(_2953_),
    .B1_N(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__o2111a_1 _3290_ (.A1(_0359_),
    .A2(_2915_),
    .B1(_0316_),
    .C1(_0363_),
    .D1(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__o21a_1 _3291_ (.A1(_0350_),
    .A2(_0358_),
    .B1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__o211a_4 _3292_ (.A1(_2953_),
    .A2(_0339_),
    .B1(_0352_),
    .C1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _3293_ (.A(_2951_),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__buf_2 _3294_ (.A(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_2 _3295_ (.A(_2950_),
    .B(_0361_),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_2 _3296_ (.A(\cu.id.cb_opcode_x[1] ),
    .Y(_0372_));
 sky130_fd_sc_hd__buf_4 _3297_ (.A(\cu.id.cb_opcode_y[2] ),
    .X(_0373_));
 sky130_fd_sc_hd__buf_4 _3298_ (.A(\cu.id.cb_opcode_y[1] ),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _3299_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__and3_1 _3300_ (.A(_0372_),
    .B(_2921_),
    .C(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__nor2_1 _3301_ (.A(_0371_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__and2b_1 _3302_ (.A_N(_2892_),
    .B(_2894_),
    .X(_0378_));
 sky130_fd_sc_hd__and2_2 _3303_ (.A(_0378_),
    .B(_0309_),
    .X(_0379_));
 sky130_fd_sc_hd__or3_1 _3304_ (.A(_0296_),
    .B(_2891_),
    .C(_0318_),
    .X(_0380_));
 sky130_fd_sc_hd__a211o_1 _3305_ (.A1(_0361_),
    .A2(_0376_),
    .B1(_2926_),
    .C1(_2928_),
    .X(_0381_));
 sky130_fd_sc_hd__o21bai_4 _3306_ (.A1(_2903_),
    .A2(_0313_),
    .B1_N(_0329_),
    .Y(_0382_));
 sky130_fd_sc_hd__or4_1 _3307_ (.A(_2905_),
    .B(_0380_),
    .C(_0381_),
    .D(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or3_2 _3308_ (.A(_0317_),
    .B(_0379_),
    .C(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _3309_ (.A(_0359_),
    .B(_2893_),
    .Y(_0385_));
 sky130_fd_sc_hd__nand2_2 _3310_ (.A(_2877_),
    .B(_2880_),
    .Y(_0386_));
 sky130_fd_sc_hd__buf_4 _3311_ (.A(\cu.id.cb_opcode_x[0] ),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _3312_ (.A(\cu.id.cb_opcode_x[1] ),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__or3_1 _3313_ (.A(_0374_),
    .B(\cu.id.cb_opcode_x[1] ),
    .C(\cu.id.cb_opcode_x[0] ),
    .X(_0389_));
 sky130_fd_sc_hd__a21oi_1 _3314_ (.A1(_0388_),
    .A2(_0389_),
    .B1(_2918_),
    .Y(_0390_));
 sky130_fd_sc_hd__a311o_1 _3315_ (.A1(_2936_),
    .A2(_0385_),
    .A3(_0386_),
    .B1(_2928_),
    .C1(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__o21ai_2 _3316_ (.A1(_2887_),
    .A2(_0391_),
    .B1(_2950_),
    .Y(_0392_));
 sky130_fd_sc_hd__or2b_1 _3317_ (.A(_0384_),
    .B_N(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _3318_ (.A(_0377_),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__buf_2 _3319_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _3320_ (.A(_0373_),
    .B(_0374_),
    .X(_0396_));
 sky130_fd_sc_hd__a211o_1 _3321_ (.A1(_0375_),
    .A2(_0396_),
    .B1(\cu.id.cb_opcode_x[1] ),
    .C1(_0387_),
    .X(_0397_));
 sky130_fd_sc_hd__a311o_1 _3322_ (.A1(_0361_),
    .A2(_0388_),
    .A3(_0397_),
    .B1(_2891_),
    .C1(_2887_),
    .X(_0398_));
 sky130_fd_sc_hd__a31o_2 _3323_ (.A1(_2893_),
    .A2(_0386_),
    .A3(_0324_),
    .B1(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_2 _3324_ (.A(_2950_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__or2_2 _3325_ (.A(_0395_),
    .B(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__a21bo_1 _3326_ (.A1(_2899_),
    .A2(_2900_),
    .B1_N(_2894_),
    .X(_0402_));
 sky130_fd_sc_hd__a21o_1 _3327_ (.A1(_2878_),
    .A2(_0402_),
    .B1(_2877_),
    .X(_0403_));
 sky130_fd_sc_hd__or3_1 _3328_ (.A(_2925_),
    .B(_2890_),
    .C(_2932_),
    .X(_0404_));
 sky130_fd_sc_hd__a21o_2 _3329_ (.A1(_0403_),
    .A2(_0404_),
    .B1(\cu.id.starting_int_service ),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _3330_ (.A(_2889_),
    .B(_2933_),
    .X(_0406_));
 sky130_fd_sc_hd__o2bb2a_2 _3331_ (.A1_N(_0299_),
    .A2_N(_0329_),
    .B1(_0406_),
    .B2(_2877_),
    .X(_0407_));
 sky130_fd_sc_hd__o22a_1 _3332_ (.A1(_2877_),
    .A2(_2878_),
    .B1(_2932_),
    .B2(_2925_),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_2 _3333_ (.A(\cu.id.starting_int_service ),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__or3_1 _3334_ (.A(_2925_),
    .B(_2932_),
    .C(_0364_),
    .X(_0410_));
 sky130_fd_sc_hd__a21o_1 _3335_ (.A1(_2900_),
    .A2(_2878_),
    .B1(_2877_),
    .X(_0411_));
 sky130_fd_sc_hd__a21o_2 _3336_ (.A1(_0410_),
    .A2(_0411_),
    .B1(\cu.id.starting_int_service ),
    .X(_0412_));
 sky130_fd_sc_hd__and4bb_4 _3337_ (.A_N(_0405_),
    .B_N(_0407_),
    .C(_0409_),
    .D(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__or3b_4 _3338_ (.A(_0293_),
    .B(_0407_),
    .C_N(_0408_),
    .X(_0414_));
 sky130_fd_sc_hd__and3b_4 _3339_ (.A_N(_0414_),
    .B(_0405_),
    .C(_0412_),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _3340_ (.A1(\cu.reg_file.reg_sp[0] ),
    .A2(_0413_),
    .B1(_0415_),
    .B2(\cu.reg_file.reg_d[0] ),
    .X(_0416_));
 sky130_fd_sc_hd__or2_4 _3341_ (.A(_0412_),
    .B(_0405_),
    .X(_0417_));
 sky130_fd_sc_hd__nor3b_4 _3342_ (.A(_0407_),
    .B(_0417_),
    .C_N(_0409_),
    .Y(_0418_));
 sky130_fd_sc_hd__nor3b_4 _3343_ (.A(_0412_),
    .B(_0414_),
    .C_N(_0405_),
    .Y(_0419_));
 sky130_fd_sc_hd__a22o_1 _3344_ (.A1(\cu.reg_file.reg_mem[0] ),
    .A2(_0418_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_4 _3345_ (.A(_0409_),
    .B(_0407_),
    .Y(_0421_));
 sky130_fd_sc_hd__a21oi_4 _3346_ (.A1(_0414_),
    .A2(_0421_),
    .B1(_0417_),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_2 _3347_ (.A(_0417_),
    .Y(_0423_));
 sky130_fd_sc_hd__a21o_1 _3348_ (.A1(_0408_),
    .A2(_0407_),
    .B1(_0293_),
    .X(_0424_));
 sky130_fd_sc_hd__or2b_2 _3349_ (.A(_0405_),
    .B_N(_0412_),
    .X(_0425_));
 sky130_fd_sc_hd__nor2_4 _3350_ (.A(_0425_),
    .B(_0421_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21o_2 _3351_ (.A1(_0423_),
    .A2(_0424_),
    .B1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__and4b_1 _3352_ (.A_N(_0412_),
    .B(_0405_),
    .C(_0409_),
    .D(_0407_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_4 _3353_ (.A(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__o21bai_4 _3354_ (.A1(_0425_),
    .A2(_0414_),
    .B1_N(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__a22o_1 _3355_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[0] ),
    .X(_0431_));
 sky130_fd_sc_hd__and3b_4 _3356_ (.A_N(_0412_),
    .B(_0405_),
    .C(_0424_),
    .X(_0432_));
 sky130_fd_sc_hd__and3_2 _3357_ (.A(_0412_),
    .B(_0405_),
    .C(_0424_),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _3358_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(_0432_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[0] ),
    .X(_0434_));
 sky130_fd_sc_hd__nor3_1 _3359_ (.A(_2940_),
    .B(_2942_),
    .C(_0379_),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _3360_ (.A(_2908_),
    .B(_0342_),
    .Y(_0436_));
 sky130_fd_sc_hd__and4bb_2 _3361_ (.A_N(_0308_),
    .B_N(_0315_),
    .C(_0435_),
    .D(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__a21oi_1 _3362_ (.A1(_2880_),
    .A2(_0437_),
    .B1(_0323_),
    .Y(_0438_));
 sky130_fd_sc_hd__or3_1 _3363_ (.A(net151),
    .B(_2914_),
    .C(_0318_),
    .X(_0439_));
 sky130_fd_sc_hd__or4_4 _3364_ (.A(_0293_),
    .B(_0362_),
    .C(_0438_),
    .D(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__a2111o_1 _3365_ (.A1(\cu.reg_file.reg_l[0] ),
    .A2(_0422_),
    .B1(_0431_),
    .C1(_0434_),
    .D1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__inv_2 _3366_ (.A(_0321_),
    .Y(_0442_));
 sky130_fd_sc_hd__or2_1 _3367_ (.A(_0328_),
    .B(_0334_),
    .X(_0443_));
 sky130_fd_sc_hd__a21o_1 _3368_ (.A1(_0442_),
    .A2(_0437_),
    .B1(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__a221o_1 _3369_ (.A1(\cu.id.cb_opcode_y[0] ),
    .A2(_0361_),
    .B1(_0444_),
    .B2(_0343_),
    .C1(_0322_),
    .X(_0445_));
 sky130_fd_sc_hd__a21bo_1 _3370_ (.A1(_2949_),
    .A2(_0445_),
    .B1_N(_0440_),
    .X(_0446_));
 sky130_fd_sc_hd__o31a_4 _3371_ (.A1(_0416_),
    .A2(_0420_),
    .A3(_0441_),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__a2111oi_1 _3372_ (.A1(_2925_),
    .A2(_0313_),
    .B1(_0325_),
    .C1(_2910_),
    .D1(_2879_),
    .Y(_0448_));
 sky130_fd_sc_hd__a32o_2 _3373_ (.A1(_2894_),
    .A2(_2874_),
    .A3(_0309_),
    .B1(_2941_),
    .B2(_0378_),
    .X(_0449_));
 sky130_fd_sc_hd__or3_1 _3374_ (.A(_0312_),
    .B(net242),
    .C(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_1 _3375_ (.A(_2878_),
    .B(_0301_),
    .Y(_0451_));
 sky130_fd_sc_hd__and3_1 _3376_ (.A(_2884_),
    .B(_2885_),
    .C(_2941_),
    .X(_0452_));
 sky130_fd_sc_hd__nor2_1 _3377_ (.A(_0452_),
    .B(_0303_),
    .Y(_0453_));
 sky130_fd_sc_hd__or4b_2 _3378_ (.A(_0379_),
    .B(_0450_),
    .C(_0451_),
    .D_N(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__or3_1 _3379_ (.A(_0298_),
    .B(_2923_),
    .C(_2901_),
    .X(_0455_));
 sky130_fd_sc_hd__o21ai_1 _3380_ (.A1(_0300_),
    .A2(_2911_),
    .B1(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__or4b_2 _3381_ (.A(\cu.id.starting_int_service ),
    .B(_0382_),
    .C(_0456_),
    .D_N(_2896_),
    .X(_0457_));
 sky130_fd_sc_hd__a21oi_4 _3382_ (.A1(net148),
    .A2(_0454_),
    .B1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__or3_1 _3383_ (.A(_2889_),
    .B(_0301_),
    .C(_2933_),
    .X(_0459_));
 sky130_fd_sc_hd__or3b_2 _3384_ (.A(_0345_),
    .B(_0450_),
    .C_N(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__o221a_1 _3385_ (.A1(_2896_),
    .A2(_0324_),
    .B1(_2912_),
    .B2(_0346_),
    .C1(_2949_),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(_0455_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21o_1 _3387_ (.A1(_0336_),
    .A2(_0460_),
    .B1(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_2 _3388_ (.A(_0458_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__and3_1 _3389_ (.A(_2892_),
    .B(_2897_),
    .C(net151),
    .X(_0465_));
 sky130_fd_sc_hd__a21oi_1 _3390_ (.A1(_0300_),
    .A2(_0353_),
    .B1(_2912_),
    .Y(_0466_));
 sky130_fd_sc_hd__a311o_1 _3391_ (.A1(_2923_),
    .A2(_0354_),
    .A3(net151),
    .B1(_0382_),
    .C1(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__nor3_2 _3392_ (.A(_0465_),
    .B(net149),
    .C(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nor2_4 _3393_ (.A(_0312_),
    .B(_0449_),
    .Y(_0469_));
 sky130_fd_sc_hd__nand2_1 _3394_ (.A(_0378_),
    .B(_0309_),
    .Y(_0470_));
 sky130_fd_sc_hd__a21o_1 _3395_ (.A1(_2878_),
    .A2(_0402_),
    .B1(_0301_),
    .X(_0471_));
 sky130_fd_sc_hd__o221a_1 _3396_ (.A1(_2918_),
    .A2(_0355_),
    .B1(_0470_),
    .B2(_2902_),
    .C1(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__a41o_4 _3397_ (.A1(net149),
    .A2(_0469_),
    .A3(_0453_),
    .A4(_0472_),
    .B1(_0293_),
    .X(_0473_));
 sky130_fd_sc_hd__a21o_1 _3398_ (.A1(_2900_),
    .A2(_2878_),
    .B1(_0301_),
    .X(_0474_));
 sky130_fd_sc_hd__o221a_1 _3399_ (.A1(\cu.id.cb_opcode_z[1] ),
    .A2(_2918_),
    .B1(_0364_),
    .B2(_0470_),
    .C1(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__or4b_1 _3400_ (.A(_0452_),
    .B(_0303_),
    .C(_0450_),
    .D_N(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__a21o_1 _3401_ (.A1(_2902_),
    .A2(_0300_),
    .B1(_2912_),
    .X(_0477_));
 sky130_fd_sc_hd__o2111ai_2 _3402_ (.A1(_2896_),
    .A2(_0364_),
    .B1(_0477_),
    .C1(_2935_),
    .D1(_2949_),
    .Y(_0478_));
 sky130_fd_sc_hd__a2111o_2 _3403_ (.A1(net241),
    .A2(_0476_),
    .B1(_0478_),
    .C1(_0382_),
    .D1(_0465_),
    .X(_0479_));
 sky130_fd_sc_hd__nor3_2 _3404_ (.A(net147),
    .B(_0473_),
    .C(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a2111oi_1 _3405_ (.A1(net149),
    .A2(_0476_),
    .B1(_0478_),
    .C1(_0382_),
    .D1(_0465_),
    .Y(_0481_));
 sky130_fd_sc_hd__nor3_4 _3406_ (.A(_0468_),
    .B(_0473_),
    .C(net146),
    .Y(_0482_));
 sky130_fd_sc_hd__a21o_1 _3407_ (.A1(net149),
    .A2(_0454_),
    .B1(_0457_),
    .X(_0483_));
 sky130_fd_sc_hd__nor2_1 _3408_ (.A(_0483_),
    .B(_0463_),
    .Y(_0484_));
 sky130_fd_sc_hd__a22o_2 _3409_ (.A1(_0464_),
    .A2(_0480_),
    .B1(_0482_),
    .B2(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__a21oi_4 _3410_ (.A1(net148),
    .A2(_0460_),
    .B1(_0462_),
    .Y(_0486_));
 sky130_fd_sc_hd__nor2_2 _3411_ (.A(_0483_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__o2111a_4 _3412_ (.A1(net147),
    .A2(_0473_),
    .B1(_0479_),
    .C1(_0486_),
    .D1(_0483_),
    .X(_0488_));
 sky130_fd_sc_hd__a21o_2 _3413_ (.A1(_0480_),
    .A2(_0487_),
    .B1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__o211a_1 _3414_ (.A1(_0464_),
    .A2(_0487_),
    .B1(_0482_),
    .C1(\cu.reg_file.reg_l[0] ),
    .X(_0490_));
 sky130_fd_sc_hd__a221o_1 _3415_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_0485_),
    .B1(_0489_),
    .B2(\cu.reg_file.reg_e[0] ),
    .C1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o2111a_4 _3416_ (.A1(net147),
    .A2(_0473_),
    .B1(net146),
    .C1(_0463_),
    .D1(_0458_),
    .X(_0492_));
 sky130_fd_sc_hd__nor2_1 _3417_ (.A(_0458_),
    .B(_0486_),
    .Y(_0493_));
 sky130_fd_sc_hd__and2_2 _3418_ (.A(_0482_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__o2111a_4 _3419_ (.A1(net147),
    .A2(_0473_),
    .B1(_0479_),
    .C1(_0463_),
    .D1(_0458_),
    .X(_0495_));
 sky130_fd_sc_hd__a32o_1 _3420_ (.A1(\cu.reg_file.reg_sp[0] ),
    .A2(_0480_),
    .A3(_0493_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0496_));
 sky130_fd_sc_hd__a221o_1 _3421_ (.A1(\cu.reg_file.reg_d[0] ),
    .A2(_0492_),
    .B1(_0494_),
    .B2(\cu.reg_file.reg_mem[0] ),
    .C1(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__o2111a_2 _3422_ (.A1(net147),
    .A2(_0473_),
    .B1(net239),
    .C1(_0486_),
    .D1(_0483_),
    .X(_0498_));
 sky130_fd_sc_hd__o2111a_4 _3423_ (.A1(net147),
    .A2(_0473_),
    .B1(net146),
    .C1(_0486_),
    .D1(_0458_),
    .X(_0499_));
 sky130_fd_sc_hd__or2_1 _3424_ (.A(\cu.id.starting_int_service ),
    .B(net150),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_4 _3425_ (.A(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__o2111a_4 _3426_ (.A1(net147),
    .A2(_0473_),
    .B1(_0479_),
    .C1(_0486_),
    .D1(_0458_),
    .X(_0502_));
 sky130_fd_sc_hd__a31o_1 _3427_ (.A1(_2913_),
    .A2(_2952_),
    .A3(_0307_),
    .B1(_0293_),
    .X(_0503_));
 sky130_fd_sc_hd__a21bo_2 _3428_ (.A1(_2948_),
    .A2(_0501_),
    .B1_N(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__a221o_1 _3429_ (.A1(\cu.pc.pc_o[0] ),
    .A2(_0501_),
    .B1(_0502_),
    .B2(\cu.reg_file.reg_b[0] ),
    .C1(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__a221o_1 _3430_ (.A1(\alu.Cin ),
    .A2(_0498_),
    .B1(_0499_),
    .B2(\cu.reg_file.reg_a[0] ),
    .C1(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__inv_2 _3431_ (.A(_0504_),
    .Y(_0507_));
 sky130_fd_sc_hd__a21o_1 _3432_ (.A1(_0343_),
    .A2(_2949_),
    .B1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__o31ai_2 _3433_ (.A1(_0491_),
    .A2(_0497_),
    .A3(_0506_),
    .B1(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__xnor2_2 _3434_ (.A(_0447_),
    .B(net143),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _3435_ (.A(\alu.Cin ),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__nor2_2 _3436_ (.A(_0395_),
    .B(_0400_),
    .Y(_0512_));
 sky130_fd_sc_hd__a21o_1 _3437_ (.A1(\alu.Cin ),
    .A2(_0512_),
    .B1(_0510_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _3438_ (.A(_0384_),
    .B(_0392_),
    .Y(_0514_));
 sky130_fd_sc_hd__or2b_1 _3439_ (.A(_0514_),
    .B_N(_0400_),
    .X(_0515_));
 sky130_fd_sc_hd__buf_8 _3440_ (.A(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_2 _3441_ (.A(_0395_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__o211a_1 _3442_ (.A1(_0401_),
    .A2(_0511_),
    .B1(_0513_),
    .C1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__or2_1 _3443_ (.A(_0384_),
    .B(_0392_),
    .X(_0519_));
 sky130_fd_sc_hd__nand2_1 _3444_ (.A(_2886_),
    .B(_0378_),
    .Y(_0520_));
 sky130_fd_sc_hd__nor2_1 _3445_ (.A(_2936_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _3446_ (.A(_0373_),
    .B(\cu.id.cb_opcode_y[0] ),
    .Y(_0522_));
 sky130_fd_sc_hd__or2_1 _3447_ (.A(_0373_),
    .B(\cu.id.cb_opcode_y[0] ),
    .X(_0523_));
 sky130_fd_sc_hd__a311o_1 _3448_ (.A1(_0372_),
    .A2(_0522_),
    .A3(_0523_),
    .B1(_0387_),
    .C1(_2918_),
    .X(_0524_));
 sky130_fd_sc_hd__a21oi_1 _3449_ (.A1(_0359_),
    .A2(_0386_),
    .B1(_2887_),
    .Y(_0525_));
 sky130_fd_sc_hd__o221a_1 _3450_ (.A1(_2925_),
    .A2(_2901_),
    .B1(_2912_),
    .B2(_2897_),
    .C1(_2935_),
    .X(_0526_));
 sky130_fd_sc_hd__and4b_1 _3451_ (.A_N(_0521_),
    .B(_0524_),
    .C(_0525_),
    .D(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _3452_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__or2_1 _3453_ (.A(_0400_),
    .B(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__or2_1 _3454_ (.A(_0519_),
    .B(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__buf_2 _3455_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__inv_2 _3456_ (.A(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__o211a_1 _3457_ (.A1(_0464_),
    .A2(_0487_),
    .B1(_0482_),
    .C1(\cu.reg_file.reg_l[1] ),
    .X(_0533_));
 sky130_fd_sc_hd__and2_1 _3458_ (.A(\cu.pc.pc_o[1] ),
    .B(_0501_),
    .X(_0534_));
 sky130_fd_sc_hd__a221o_1 _3459_ (.A1(\cu.reg_file.reg_e[1] ),
    .A2(_0488_),
    .B1(_0502_),
    .B2(\cu.reg_file.reg_b[1] ),
    .C1(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_4 _3460_ (.A(_0504_),
    .X(_0536_));
 sky130_fd_sc_hd__a2111o_1 _3461_ (.A1(\cu.reg_file.reg_c[1] ),
    .A2(_0485_),
    .B1(_0533_),
    .C1(_0535_),
    .D1(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__a22o_1 _3462_ (.A1(\cu.reg_file.reg_d[1] ),
    .A2(_0492_),
    .B1(_0498_),
    .B2(\cu.alu_f[1] ),
    .X(_0538_));
 sky130_fd_sc_hd__and2_2 _3463_ (.A(_0480_),
    .B(_0493_),
    .X(_0539_));
 sky130_fd_sc_hd__and2_1 _3464_ (.A(\cu.reg_file.reg_a[1] ),
    .B(_0499_),
    .X(_0540_));
 sky130_fd_sc_hd__and3_1 _3465_ (.A(\cu.reg_file.reg_e[1] ),
    .B(_0480_),
    .C(_0487_),
    .X(_0541_));
 sky130_fd_sc_hd__a32o_1 _3466_ (.A1(\cu.reg_file.reg_mem[1] ),
    .A2(_0482_),
    .A3(_0493_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_h[1] ),
    .X(_0542_));
 sky130_fd_sc_hd__a2111o_1 _3467_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_0539_),
    .B1(_0540_),
    .C1(_0541_),
    .D1(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__o21ai_1 _3468_ (.A1(_0294_),
    .A2(_0360_),
    .B1(_0536_),
    .Y(_0544_));
 sky130_fd_sc_hd__o31a_4 _3469_ (.A1(_0537_),
    .A2(_0538_),
    .A3(_0543_),
    .B1(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__or2_2 _3470_ (.A(_0296_),
    .B(_0528_),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_2 _3471_ (.A(_0399_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__or2_1 _3472_ (.A(_0371_),
    .B(_0376_),
    .X(_0548_));
 sky130_fd_sc_hd__nor2_1 _3473_ (.A(_0548_),
    .B(_0393_),
    .Y(_0549_));
 sky130_fd_sc_hd__and2b_1 _3474_ (.A_N(_0392_),
    .B(_0384_),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_1 _3475_ (.A(_0399_),
    .B(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__nor2_1 _3476_ (.A(_0528_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__or2b_1 _3477_ (.A(_0400_),
    .B_N(_0528_),
    .X(_0553_));
 sky130_fd_sc_hd__nor2_1 _3478_ (.A(_0514_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__and2_1 _3479_ (.A(_0400_),
    .B(_0546_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _3480_ (.A(_0550_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_2 _3481_ (.A(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__a2111o_4 _3482_ (.A1(_0547_),
    .A2(_0549_),
    .B1(_0552_),
    .C1(_0554_),
    .D1(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__o211a_1 _3483_ (.A1(_0464_),
    .A2(_0487_),
    .B1(_0482_),
    .C1(\cu.reg_file.reg_l[7] ),
    .X(_0559_));
 sky130_fd_sc_hd__a221o_1 _3484_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_0485_),
    .B1(_0489_),
    .B2(\cu.reg_file.reg_e[7] ),
    .C1(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a22o_1 _3485_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(_0502_),
    .B1(_0492_),
    .B2(\cu.reg_file.reg_d[7] ),
    .X(_0561_));
 sky130_fd_sc_hd__a221o_1 _3486_ (.A1(\cu.reg_file.reg_h[7] ),
    .A2(_0495_),
    .B1(_0539_),
    .B2(\cu.reg_file.reg_sp[7] ),
    .C1(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__a221o_1 _3487_ (.A1(\cu.pc.pc_o[7] ),
    .A2(_0501_),
    .B1(_0498_),
    .B2(\cu.alu_f[7] ),
    .C1(_0504_),
    .X(_0563_));
 sky130_fd_sc_hd__a221o_1 _3488_ (.A1(\cu.reg_file.reg_a[7] ),
    .A2(_0499_),
    .B1(_0494_),
    .B2(\cu.reg_file.reg_mem[7] ),
    .C1(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__o21ai_1 _3489_ (.A1(_0294_),
    .A2(_0372_),
    .B1(_0536_),
    .Y(_0565_));
 sky130_fd_sc_hd__o31a_4 _3490_ (.A1(_0560_),
    .A2(_0562_),
    .A3(_0564_),
    .B1(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__and3_1 _3491_ (.A(_0566_),
    .B(_0547_),
    .C(_0550_),
    .X(_0567_));
 sky130_fd_sc_hd__a221o_1 _3492_ (.A1(net143),
    .A2(_0532_),
    .B1(_0545_),
    .B2(_0558_),
    .C1(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__or2_1 _3493_ (.A(_0519_),
    .B(_0553_),
    .X(_0569_));
 sky130_fd_sc_hd__buf_2 _3494_ (.A(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__and2b_1 _3495_ (.A_N(_0570_),
    .B(_0510_),
    .X(_0571_));
 sky130_fd_sc_hd__inv_2 _3496_ (.A(\alu.Cin ),
    .Y(_0572_));
 sky130_fd_sc_hd__or2_1 _3497_ (.A(_0514_),
    .B(_0529_),
    .X(_0573_));
 sky130_fd_sc_hd__inv_2 _3498_ (.A(net143),
    .Y(_0574_));
 sky130_fd_sc_hd__o31ai_2 _3499_ (.A1(_0416_),
    .A2(_0420_),
    .A3(_0441_),
    .B1(_0446_),
    .Y(_0575_));
 sky130_fd_sc_hd__clkbuf_4 _3500_ (.A(_0440_),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _3501_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[2] ),
    .X(_0577_));
 sky130_fd_sc_hd__a22o_1 _3502_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(_0432_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[2] ),
    .X(_0578_));
 sky130_fd_sc_hd__a221o_1 _3503_ (.A1(\cu.reg_file.reg_sp[2] ),
    .A2(_0413_),
    .B1(_0415_),
    .B2(\cu.reg_file.reg_d[2] ),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__a22o_1 _3504_ (.A1(\cu.reg_file.reg_mem[2] ),
    .A2(_0418_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[2] ),
    .X(_0580_));
 sky130_fd_sc_hd__a2111o_1 _3505_ (.A1(\cu.reg_file.reg_l[2] ),
    .A2(_0422_),
    .B1(_0577_),
    .C1(_0579_),
    .D1(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__a21o_1 _3506_ (.A1(_0341_),
    .A2(_0443_),
    .B1(_0336_),
    .X(_0582_));
 sky130_fd_sc_hd__or4_4 _3507_ (.A(_0321_),
    .B(_0322_),
    .C(_0328_),
    .D(_0334_),
    .X(_0583_));
 sky130_fd_sc_hd__a221o_1 _3508_ (.A1(\cu.id.cb_opcode_y[2] ),
    .A2(_0361_),
    .B1(_0437_),
    .B2(_0341_),
    .C1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__nand2_1 _3509_ (.A(_0582_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__o21ai_1 _3510_ (.A1(_0294_),
    .A2(_0585_),
    .B1(_0576_),
    .Y(_0586_));
 sky130_fd_sc_hd__o21ai_2 _3511_ (.A1(_0576_),
    .A2(_0581_),
    .B1(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__buf_2 _3512_ (.A(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__a22o_1 _3513_ (.A1(\cu.reg_file.reg_c[1] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[1] ),
    .X(_0589_));
 sky130_fd_sc_hd__a22o_1 _3514_ (.A1(\cu.reg_file.reg_mem[1] ),
    .A2(_0418_),
    .B1(_0415_),
    .B2(\cu.reg_file.reg_d[1] ),
    .X(_0590_));
 sky130_fd_sc_hd__a221o_1 _3515_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_0413_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[1] ),
    .C1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__a22o_1 _3516_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_0432_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[1] ),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_1 _3517_ (.A1(\cu.reg_file.reg_l[1] ),
    .A2(_0422_),
    .B1(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__a21o_1 _3518_ (.A1(_0340_),
    .A2(_0443_),
    .B1(_0336_),
    .X(_0594_));
 sky130_fd_sc_hd__a221o_1 _3519_ (.A1(\cu.id.cb_opcode_y[1] ),
    .A2(_0361_),
    .B1(_0437_),
    .B2(_0340_),
    .C1(_0583_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _3520_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__o21ai_1 _3521_ (.A1(_0293_),
    .A2(_0596_),
    .B1(_0440_),
    .Y(_0597_));
 sky130_fd_sc_hd__o41a_4 _3522_ (.A1(_0440_),
    .A2(_0589_),
    .A3(_0591_),
    .A4(_0593_),
    .B1(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__buf_2 _3523_ (.A(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__inv_2 _3524_ (.A(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__and3_1 _3525_ (.A(_0575_),
    .B(_0588_),
    .C(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__or2b_2 _3526_ (.A(_0519_),
    .B_N(_0555_),
    .X(_0602_));
 sky130_fd_sc_hd__nor2_2 _3527_ (.A(_0548_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(_0447_),
    .A1(_0601_),
    .S(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__or2_1 _3529_ (.A(_0399_),
    .B(_0546_),
    .X(_0605_));
 sky130_fd_sc_hd__nor2_2 _3530_ (.A(_0519_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__or2_2 _3531_ (.A(_0603_),
    .B(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__o21ai_1 _3532_ (.A1(_0574_),
    .A2(_0604_),
    .B1(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__or3_1 _3533_ (.A(_0548_),
    .B(_0393_),
    .C(_0529_),
    .X(_0609_));
 sky130_fd_sc_hd__buf_2 _3534_ (.A(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_4 _3535_ (.A(_0377_),
    .B(_0602_),
    .Y(_0611_));
 sky130_fd_sc_hd__nand2_1 _3536_ (.A(_0447_),
    .B(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__a211o_1 _3537_ (.A1(_0610_),
    .A2(_0612_),
    .B1(net143),
    .C1(_0601_),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_1 _3538_ (.A(_0549_),
    .B(_0555_),
    .Y(_0614_));
 sky130_fd_sc_hd__o2111a_1 _3539_ (.A1(_0572_),
    .A2(_0573_),
    .B1(_0608_),
    .C1(_0613_),
    .D1(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__or4b_1 _3540_ (.A(_0518_),
    .B(_0568_),
    .C(_0571_),
    .D_N(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_4 _3541_ (.A(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_4 _3542_ (.A(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__buf_4 _3543_ (.A(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__nor2_1 _3544_ (.A(_0377_),
    .B(_0393_),
    .Y(_0620_));
 sky130_fd_sc_hd__o21a_1 _3545_ (.A1(_0464_),
    .A2(_0487_),
    .B1(_0482_),
    .X(_0621_));
 sky130_fd_sc_hd__a22o_1 _3546_ (.A1(\cu.reg_file.reg_e[6] ),
    .A2(_0489_),
    .B1(_0621_),
    .B2(\cu.reg_file.reg_l[6] ),
    .X(_0622_));
 sky130_fd_sc_hd__a21o_1 _3547_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_0485_),
    .B1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_4 _3548_ (.A(_0539_),
    .X(_0624_));
 sky130_fd_sc_hd__clkbuf_4 _3549_ (.A(_0498_),
    .X(_0625_));
 sky130_fd_sc_hd__a22o_1 _3550_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_0492_),
    .B1(_0625_),
    .B2(\cu.alu_f[6] ),
    .X(_0626_));
 sky130_fd_sc_hd__a221o_1 _3551_ (.A1(\cu.reg_file.reg_h[6] ),
    .A2(_0495_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[6] ),
    .C1(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_4 _3552_ (.A(_0494_),
    .X(_0628_));
 sky130_fd_sc_hd__a221o_1 _3553_ (.A1(\cu.pc.pc_o[6] ),
    .A2(_0501_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[6] ),
    .C1(_0536_),
    .X(_0629_));
 sky130_fd_sc_hd__a221o_1 _3554_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(_0502_),
    .B1(_0499_),
    .B2(\cu.reg_file.reg_a[6] ),
    .C1(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__o21ai_1 _3555_ (.A1(_0295_),
    .A2(_2921_),
    .B1(_0536_),
    .Y(_0631_));
 sky130_fd_sc_hd__o31a_4 _3556_ (.A1(_0623_),
    .A2(_0627_),
    .A3(_0630_),
    .B1(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__nand2_1 _3557_ (.A(_0442_),
    .B(_0437_),
    .Y(_0633_));
 sky130_fd_sc_hd__o21ba_1 _3558_ (.A1(_0322_),
    .A2(_0633_),
    .B1_N(_0443_),
    .X(_0634_));
 sky130_fd_sc_hd__or3_1 _3559_ (.A(_0295_),
    .B(_2921_),
    .C(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_4 _3560_ (.A(_0413_),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_1 _3561_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_0415_),
    .B1(_0432_),
    .B2(\cu.reg_file.reg_b[6] ),
    .X(_0637_));
 sky130_fd_sc_hd__a221o_1 _3562_ (.A1(\cu.reg_file.reg_sp[6] ),
    .A2(_0636_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[6] ),
    .C1(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__a22o_1 _3563_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[6] ),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_8 _3564_ (.A(_0418_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _3565_ (.A1(\cu.reg_file.reg_mem[6] ),
    .A2(_0640_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[6] ),
    .X(_0641_));
 sky130_fd_sc_hd__a2111o_1 _3566_ (.A1(\cu.reg_file.reg_l[6] ),
    .A2(_0422_),
    .B1(_0639_),
    .C1(_0641_),
    .D1(_0576_),
    .X(_0642_));
 sky130_fd_sc_hd__o2bb2a_2 _3567_ (.A1_N(_0576_),
    .A2_N(_0635_),
    .B1(_0638_),
    .B2(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__xnor2_2 _3568_ (.A(_0632_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__inv_2 _3569_ (.A(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__or3b_1 _3570_ (.A(_0295_),
    .B(_0634_),
    .C_N(_0373_),
    .X(_0646_));
 sky130_fd_sc_hd__a22o_1 _3571_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_0415_),
    .B1(_0432_),
    .B2(\cu.reg_file.reg_b[5] ),
    .X(_0647_));
 sky130_fd_sc_hd__a221o_1 _3572_ (.A1(\cu.reg_file.reg_sp[5] ),
    .A2(_0636_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[5] ),
    .C1(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__a22o_1 _3573_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[5] ),
    .X(_0649_));
 sky130_fd_sc_hd__a22o_1 _3574_ (.A1(\cu.reg_file.reg_mem[5] ),
    .A2(_0640_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[5] ),
    .X(_0650_));
 sky130_fd_sc_hd__a2111o_1 _3575_ (.A1(\cu.reg_file.reg_l[5] ),
    .A2(_0422_),
    .B1(_0649_),
    .C1(_0650_),
    .D1(_0576_),
    .X(_0651_));
 sky130_fd_sc_hd__o2bb2a_4 _3576_ (.A1_N(_0576_),
    .A2_N(_0646_),
    .B1(_0648_),
    .B2(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__buf_8 _3577_ (.A(_0507_),
    .X(_0653_));
 sky130_fd_sc_hd__or2_1 _3578_ (.A(\ih.interrupt_source[3] ),
    .B(\ih.interrupt_source[1] ),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(\cu.id.cb_opcode_y[2] ),
    .A1(_0654_),
    .S(_0294_),
    .X(_0655_));
 sky130_fd_sc_hd__and2_1 _3580_ (.A(\cu.pc.pc_o[5] ),
    .B(_0501_),
    .X(_0656_));
 sky130_fd_sc_hd__a221o_1 _3581_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_0492_),
    .B1(_0625_),
    .B2(\cu.alu_f[5] ),
    .C1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__a22o_1 _3582_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(_0502_),
    .B1(_0499_),
    .B2(\cu.reg_file.reg_a[5] ),
    .X(_0658_));
 sky130_fd_sc_hd__a221o_1 _3583_ (.A1(\cu.reg_file.reg_sp[5] ),
    .A2(_0539_),
    .B1(_0494_),
    .B2(\cu.reg_file.reg_mem[5] ),
    .C1(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__a221o_1 _3584_ (.A1(\cu.reg_file.reg_e[5] ),
    .A2(_0489_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_h[5] ),
    .C1(_0536_),
    .X(_0660_));
 sky130_fd_sc_hd__a22o_1 _3585_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_0485_),
    .B1(_0621_),
    .B2(\cu.reg_file.reg_l[5] ),
    .X(_0661_));
 sky130_fd_sc_hd__or3_2 _3586_ (.A(_0659_),
    .B(_0660_),
    .C(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__o22a_4 _3587_ (.A1(_0653_),
    .A2(_0655_),
    .B1(_0657_),
    .B2(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__xnor2_4 _3588_ (.A(_0652_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__or3b_1 _3589_ (.A(_0294_),
    .B(_0634_),
    .C_N(_0374_),
    .X(_0665_));
 sky130_fd_sc_hd__a22o_1 _3590_ (.A1(\cu.reg_file.reg_d[4] ),
    .A2(_0415_),
    .B1(_0432_),
    .B2(\cu.reg_file.reg_b[4] ),
    .X(_0666_));
 sky130_fd_sc_hd__a221o_1 _3591_ (.A1(\cu.reg_file.reg_sp[4] ),
    .A2(_0413_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[4] ),
    .C1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_1 _3592_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[4] ),
    .X(_0668_));
 sky130_fd_sc_hd__a22o_1 _3593_ (.A1(\cu.reg_file.reg_mem[4] ),
    .A2(_0418_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[4] ),
    .X(_0669_));
 sky130_fd_sc_hd__a2111o_1 _3594_ (.A1(\cu.reg_file.reg_l[4] ),
    .A2(_0422_),
    .B1(_0668_),
    .C1(_0669_),
    .D1(_0576_),
    .X(_0670_));
 sky130_fd_sc_hd__o2bb2a_1 _3595_ (.A1_N(_0576_),
    .A2_N(_0665_),
    .B1(_0667_),
    .B2(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__or2_1 _3596_ (.A(\ih.interrupt_source[3] ),
    .B(\ih.interrupt_source[2] ),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(_0374_),
    .A1(_0672_),
    .S(_0294_),
    .X(_0673_));
 sky130_fd_sc_hd__a22o_1 _3598_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_0485_),
    .B1(_0489_),
    .B2(\cu.reg_file.reg_e[4] ),
    .X(_0674_));
 sky130_fd_sc_hd__a21o_1 _3599_ (.A1(\cu.reg_file.reg_l[4] ),
    .A2(_0621_),
    .B1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__a22o_1 _3600_ (.A1(\cu.reg_file.reg_h[4] ),
    .A2(_0495_),
    .B1(_0498_),
    .B2(\cu.alu_f[4] ),
    .X(_0676_));
 sky130_fd_sc_hd__a221o_1 _3601_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(_0502_),
    .B1(_0494_),
    .B2(\cu.reg_file.reg_mem[4] ),
    .C1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__a221o_1 _3602_ (.A1(\cu.pc.pc_o[4] ),
    .A2(_0501_),
    .B1(_0499_),
    .B2(\cu.reg_file.reg_a[4] ),
    .C1(_0504_),
    .X(_0678_));
 sky130_fd_sc_hd__a221o_1 _3603_ (.A1(\cu.reg_file.reg_sp[4] ),
    .A2(_0539_),
    .B1(_0492_),
    .B2(\cu.reg_file.reg_d[4] ),
    .C1(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__or2_1 _3604_ (.A(_0677_),
    .B(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__o22a_2 _3605_ (.A1(_0653_),
    .A2(_0673_),
    .B1(_0675_),
    .B2(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__and2b_1 _3606_ (.A_N(_0671_),
    .B(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__and2b_1 _3607_ (.A_N(_0681_),
    .B(_0671_),
    .X(_0683_));
 sky130_fd_sc_hd__nor2_2 _3608_ (.A(_0682_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__nor2_1 _3609_ (.A(_0664_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__o211a_1 _3610_ (.A1(_0464_),
    .A2(_0487_),
    .B1(_0482_),
    .C1(\cu.reg_file.reg_l[3] ),
    .X(_0686_));
 sky130_fd_sc_hd__a221o_1 _3611_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_0485_),
    .B1(_0489_),
    .B2(\cu.reg_file.reg_e[3] ),
    .C1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__a22o_1 _3612_ (.A1(\cu.reg_file.reg_h[3] ),
    .A2(_0495_),
    .B1(_0499_),
    .B2(\cu.reg_file.reg_a[3] ),
    .X(_0688_));
 sky130_fd_sc_hd__a221o_1 _3613_ (.A1(\cu.alu_f[3] ),
    .A2(_0498_),
    .B1(_0494_),
    .B2(\cu.reg_file.reg_mem[3] ),
    .C1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__a221o_1 _3614_ (.A1(\cu.pc.pc_o[3] ),
    .A2(_0501_),
    .B1(_0502_),
    .B2(\cu.reg_file.reg_b[3] ),
    .C1(_0536_),
    .X(_0690_));
 sky130_fd_sc_hd__a221o_1 _3615_ (.A1(\cu.reg_file.reg_sp[3] ),
    .A2(_0539_),
    .B1(_0492_),
    .B2(\cu.reg_file.reg_d[3] ),
    .C1(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__inv_2 _3616_ (.A(\cu.id.cb_opcode_y[0] ),
    .Y(_0692_));
 sky130_fd_sc_hd__o21ai_1 _3617_ (.A1(_0294_),
    .A2(_0692_),
    .B1(_0536_),
    .Y(_0693_));
 sky130_fd_sc_hd__o31a_4 _3618_ (.A1(_0687_),
    .A2(_0689_),
    .A3(_0691_),
    .B1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__or3_1 _3619_ (.A(_0294_),
    .B(_0692_),
    .C(_0634_),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _3620_ (.A1(\cu.reg_file.reg_d[3] ),
    .A2(_0415_),
    .B1(_0432_),
    .B2(\cu.reg_file.reg_b[3] ),
    .X(_0696_));
 sky130_fd_sc_hd__a221o_1 _3621_ (.A1(\cu.reg_file.reg_sp[3] ),
    .A2(_0413_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[3] ),
    .C1(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__a22o_1 _3622_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[3] ),
    .X(_0698_));
 sky130_fd_sc_hd__a22o_1 _3623_ (.A1(\cu.reg_file.reg_mem[3] ),
    .A2(_0418_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[3] ),
    .X(_0699_));
 sky130_fd_sc_hd__a2111o_1 _3624_ (.A1(\cu.reg_file.reg_l[3] ),
    .A2(_0422_),
    .B1(_0698_),
    .C1(_0699_),
    .D1(_0440_),
    .X(_0700_));
 sky130_fd_sc_hd__o2bb2a_2 _3625_ (.A1_N(_0576_),
    .A2_N(_0695_),
    .B1(_0697_),
    .B2(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nor2_1 _3626_ (.A(_0694_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__o211a_1 _3627_ (.A1(_0464_),
    .A2(_0487_),
    .B1(_0482_),
    .C1(\cu.reg_file.reg_l[2] ),
    .X(_0703_));
 sky130_fd_sc_hd__a221o_1 _3628_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_0485_),
    .B1(_0489_),
    .B2(\cu.reg_file.reg_e[2] ),
    .C1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__a22o_1 _3629_ (.A1(\cu.reg_file.reg_h[2] ),
    .A2(_0495_),
    .B1(_0499_),
    .B2(\cu.reg_file.reg_a[2] ),
    .X(_0705_));
 sky130_fd_sc_hd__a221o_1 _3630_ (.A1(\cu.alu_f[2] ),
    .A2(_0498_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[2] ),
    .C1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__a221o_1 _3631_ (.A1(\cu.pc.pc_o[2] ),
    .A2(_0501_),
    .B1(_0502_),
    .B2(\cu.reg_file.reg_b[2] ),
    .C1(_0536_),
    .X(_0707_));
 sky130_fd_sc_hd__a221o_1 _3632_ (.A1(\cu.reg_file.reg_sp[2] ),
    .A2(_0624_),
    .B1(_0492_),
    .B2(\cu.reg_file.reg_d[2] ),
    .C1(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__a21o_1 _3633_ (.A1(_2950_),
    .A2(_0341_),
    .B1(_0507_),
    .X(_0709_));
 sky130_fd_sc_hd__o31ai_4 _3634_ (.A1(_0704_),
    .A2(_0706_),
    .A3(_0708_),
    .B1(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _3635_ (.A(_0587_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__xnor2_4 _3636_ (.A(_0545_),
    .B(_0598_),
    .Y(_0712_));
 sky130_fd_sc_hd__or2_1 _3637_ (.A(_0575_),
    .B(net143),
    .X(_0713_));
 sky130_fd_sc_hd__a2bb2o_1 _3638_ (.A1_N(_0712_),
    .A2_N(_0713_),
    .B1(_0545_),
    .B2(_0599_),
    .X(_0714_));
 sky130_fd_sc_hd__nor2_1 _3639_ (.A(_0587_),
    .B(_0710_),
    .Y(_0715_));
 sky130_fd_sc_hd__a21oi_2 _3640_ (.A1(_0711_),
    .A2(_0714_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nand2_1 _3641_ (.A(_0694_),
    .B(_0701_),
    .Y(_0717_));
 sky130_fd_sc_hd__o21ai_2 _3642_ (.A1(_0702_),
    .A2(_0716_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__nor2_1 _3643_ (.A(_0652_),
    .B(_0663_),
    .Y(_0719_));
 sky130_fd_sc_hd__and2_1 _3644_ (.A(_0671_),
    .B(_0681_),
    .X(_0720_));
 sky130_fd_sc_hd__and2b_1 _3645_ (.A_N(_0719_),
    .B(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__a221o_1 _3646_ (.A1(_0652_),
    .A2(_0663_),
    .B1(_0685_),
    .B2(_0718_),
    .C1(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__or3_1 _3647_ (.A(_0293_),
    .B(_0372_),
    .C(_0634_),
    .X(_0723_));
 sky130_fd_sc_hd__a22o_1 _3648_ (.A1(\cu.reg_file.reg_d[7] ),
    .A2(_0415_),
    .B1(_0432_),
    .B2(\cu.reg_file.reg_b[7] ),
    .X(_0724_));
 sky130_fd_sc_hd__a221o_1 _3649_ (.A1(\cu.reg_file.reg_sp[7] ),
    .A2(_0413_),
    .B1(_0419_),
    .B2(\cu.reg_file.reg_h[7] ),
    .C1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__a22o_1 _3650_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_e[7] ),
    .X(_0726_));
 sky130_fd_sc_hd__a22o_1 _3651_ (.A1(\cu.reg_file.reg_mem[7] ),
    .A2(_0418_),
    .B1(_0433_),
    .B2(\cu.reg_file.reg_a[7] ),
    .X(_0727_));
 sky130_fd_sc_hd__a2111o_1 _3652_ (.A1(\cu.reg_file.reg_l[7] ),
    .A2(_0422_),
    .B1(_0726_),
    .C1(_0727_),
    .D1(_0440_),
    .X(_0728_));
 sky130_fd_sc_hd__o2bb2a_2 _3653_ (.A1_N(_0576_),
    .A2_N(_0723_),
    .B1(_0725_),
    .B2(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__and2_1 _3654_ (.A(_0566_),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__nor2_1 _3655_ (.A(_0566_),
    .B(_0729_),
    .Y(_0731_));
 sky130_fd_sc_hd__or2_1 _3656_ (.A(_0730_),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__buf_2 _3657_ (.A(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__inv_2 _3658_ (.A(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__and2_1 _3659_ (.A(_0632_),
    .B(_0643_),
    .X(_0735_));
 sky130_fd_sc_hd__and2b_1 _3660_ (.A_N(_0731_),
    .B(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__a311o_1 _3661_ (.A1(_0645_),
    .A2(_0722_),
    .A3(_0734_),
    .B1(_0736_),
    .C1(_0730_),
    .X(_0737_));
 sky130_fd_sc_hd__and3_1 _3662_ (.A(_2950_),
    .B(_2913_),
    .C(_0536_),
    .X(_0738_));
 sky130_fd_sc_hd__clkbuf_8 _3663_ (.A(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__buf_4 _3664_ (.A(_0501_),
    .X(_0740_));
 sky130_fd_sc_hd__and2_2 _3665_ (.A(_0464_),
    .B(_0482_),
    .X(_0741_));
 sky130_fd_sc_hd__a22o_1 _3666_ (.A1(\cu.reg_file.reg_d[0] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0742_));
 sky130_fd_sc_hd__and2_2 _3667_ (.A(_0464_),
    .B(_0480_),
    .X(_0743_));
 sky130_fd_sc_hd__a22o_1 _3668_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[8] ),
    .X(_0744_));
 sky130_fd_sc_hd__a211o_1 _3669_ (.A1(\cu.pc.pc_o[8] ),
    .A2(_0740_),
    .B1(_0742_),
    .C1(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__a221o_1 _3670_ (.A1(\cu.reg_file.reg_a[0] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[8] ),
    .C1(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__a22oi_4 _3671_ (.A1(\cu.id.imm_i[8] ),
    .A2(_0739_),
    .B1(_0746_),
    .B2(_0653_),
    .Y(_0747_));
 sky130_fd_sc_hd__nor2_4 _3672_ (.A(_0417_),
    .B(_0421_),
    .Y(_0748_));
 sky130_fd_sc_hd__a22o_1 _3673_ (.A1(\cu.reg_file.reg_sp[8] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _3674_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[0] ),
    .X(_0750_));
 sky130_fd_sc_hd__a211oi_4 _3675_ (.A1(\cu.reg_file.reg_mem[8] ),
    .A2(_0640_),
    .B1(_0749_),
    .C1(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__xor2_4 _3676_ (.A(_0747_),
    .B(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__xor2_1 _3677_ (.A(_0737_),
    .B(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__xnor2_1 _3678_ (.A(_0645_),
    .B(_0722_),
    .Y(_0754_));
 sky130_fd_sc_hd__inv_2 _3679_ (.A(_0684_),
    .Y(_0755_));
 sky130_fd_sc_hd__a21oi_1 _3680_ (.A1(_0718_),
    .A2(_0755_),
    .B1(_0720_),
    .Y(_0756_));
 sky130_fd_sc_hd__xnor2_1 _3681_ (.A(_0664_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__nor2_1 _3682_ (.A(_0511_),
    .B(_0712_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand2b_2 _3683_ (.A_N(_0715_),
    .B(_0711_),
    .Y(_0759_));
 sky130_fd_sc_hd__xnor2_1 _3684_ (.A(_0714_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _3685_ (.A(_0758_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__xor2_1 _3686_ (.A(_0694_),
    .B(_0701_),
    .X(_0762_));
 sky130_fd_sc_hd__inv_2 _3687_ (.A(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__xnor2_1 _3688_ (.A(_0716_),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__nor2_1 _3689_ (.A(_0761_),
    .B(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__xnor2_1 _3690_ (.A(_0718_),
    .B(_0684_),
    .Y(_0766_));
 sky130_fd_sc_hd__nand2_1 _3691_ (.A(_0765_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__or3_1 _3692_ (.A(_0754_),
    .B(_0757_),
    .C(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__a21o_1 _3693_ (.A1(_0645_),
    .A2(_0722_),
    .B1(_0735_),
    .X(_0769_));
 sky130_fd_sc_hd__xnor2_2 _3694_ (.A(_0769_),
    .B(_0734_),
    .Y(_0770_));
 sky130_fd_sc_hd__or3b_1 _3695_ (.A(_0768_),
    .B(_0770_),
    .C_N(_0753_),
    .X(_0771_));
 sky130_fd_sc_hd__and2_1 _3696_ (.A(_0512_),
    .B(_0528_),
    .X(_0772_));
 sky130_fd_sc_hd__clkbuf_4 _3697_ (.A(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__or2_2 _3698_ (.A(_0514_),
    .B(_0605_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _3699_ (.A(_0620_),
    .B(_0547_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_4 _3700_ (.A(_0774_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_2 _3701_ (.A(_0512_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__a21o_1 _3702_ (.A1(_0771_),
    .A2(_0773_),
    .B1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__nand2_2 _3703_ (.A(_0512_),
    .B(_0528_),
    .Y(_0779_));
 sky130_fd_sc_hd__nor4_1 _3704_ (.A(_0768_),
    .B(_0770_),
    .C(_0753_),
    .D(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand2_1 _3705_ (.A(_0447_),
    .B(net143),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_1 _3706_ (.A(_0545_),
    .B(_0600_),
    .Y(_0782_));
 sky130_fd_sc_hd__a21bo_1 _3707_ (.A1(_0781_),
    .A2(_0712_),
    .B1_N(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__and2b_1 _3708_ (.A_N(_0710_),
    .B(_0587_),
    .X(_0784_));
 sky130_fd_sc_hd__and2b_1 _3709_ (.A_N(_0762_),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__and2b_1 _3710_ (.A_N(_0701_),
    .B(_0694_),
    .X(_0786_));
 sky130_fd_sc_hd__a311o_2 _3711_ (.A1(_0759_),
    .A2(_0763_),
    .A3(_0783_),
    .B1(_0785_),
    .C1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_1 _3712_ (.A(_0644_),
    .B(_0733_),
    .X(_0788_));
 sky130_fd_sc_hd__nand4_1 _3713_ (.A(_0664_),
    .B(_0684_),
    .C(_0787_),
    .D(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__and2b_1 _3714_ (.A_N(_0643_),
    .B(_0632_),
    .X(_0790_));
 sky130_fd_sc_hd__inv_2 _3715_ (.A(_0566_),
    .Y(_0791_));
 sky130_fd_sc_hd__o2bb2a_1 _3716_ (.A1_N(_0733_),
    .A2_N(_0790_),
    .B1(_0729_),
    .B2(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__and2b_1 _3717_ (.A_N(_0652_),
    .B(_0663_),
    .X(_0793_));
 sky130_fd_sc_hd__a21o_1 _3718_ (.A1(_0664_),
    .A2(_0682_),
    .B1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__nand2_1 _3719_ (.A(_0788_),
    .B(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__a31o_1 _3720_ (.A1(_0789_),
    .A2(_0792_),
    .A3(_0795_),
    .B1(_0752_),
    .X(_0796_));
 sky130_fd_sc_hd__nand4_1 _3721_ (.A(_0752_),
    .B(_0789_),
    .C(_0792_),
    .D(_0795_),
    .Y(_0797_));
 sky130_fd_sc_hd__and2_1 _3722_ (.A(_0796_),
    .B(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__a31o_1 _3723_ (.A1(_0664_),
    .A2(_0684_),
    .A3(_0787_),
    .B1(_0794_),
    .X(_0799_));
 sky130_fd_sc_hd__a21oi_1 _3724_ (.A1(_0644_),
    .A2(_0799_),
    .B1(_0790_),
    .Y(_0800_));
 sky130_fd_sc_hd__xnor2_2 _3725_ (.A(_0733_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__xnor2_1 _3726_ (.A(_0645_),
    .B(_0799_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21oi_1 _3727_ (.A1(_0684_),
    .A2(_0787_),
    .B1(_0682_),
    .Y(_0803_));
 sky130_fd_sc_hd__xnor2_1 _3728_ (.A(_0664_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__xnor2_1 _3729_ (.A(_0755_),
    .B(_0787_),
    .Y(_0805_));
 sky130_fd_sc_hd__xor2_1 _3730_ (.A(_0759_),
    .B(_0783_),
    .X(_0806_));
 sky130_fd_sc_hd__or3b_1 _3731_ (.A(_0572_),
    .B(_0510_),
    .C_N(_0712_),
    .X(_0807_));
 sky130_fd_sc_hd__or2_1 _3732_ (.A(_0806_),
    .B(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__a21oi_1 _3733_ (.A1(_0759_),
    .A2(_0783_),
    .B1(_0784_),
    .Y(_0809_));
 sky130_fd_sc_hd__xnor2_1 _3734_ (.A(_0763_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__or3_2 _3735_ (.A(_0805_),
    .B(_0808_),
    .C(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__or3_2 _3736_ (.A(_0802_),
    .B(_0804_),
    .C(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__or3_1 _3737_ (.A(_0801_),
    .B(_0812_),
    .C(_0798_),
    .X(_0813_));
 sky130_fd_sc_hd__o21ai_1 _3738_ (.A1(_0801_),
    .A2(_0812_),
    .B1(_0798_),
    .Y(_0814_));
 sky130_fd_sc_hd__nand2_1 _3739_ (.A(_0813_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__nor2_1 _3740_ (.A(_0401_),
    .B(_0528_),
    .Y(_0816_));
 sky130_fd_sc_hd__buf_2 _3741_ (.A(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__a22o_1 _3742_ (.A1(_0776_),
    .A2(_0798_),
    .B1(_0815_),
    .B2(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__a211o_1 _3743_ (.A1(_0753_),
    .A2(_0778_),
    .B1(_0780_),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__nand2_1 _3744_ (.A(_0605_),
    .B(_0553_),
    .Y(_0820_));
 sky130_fd_sc_hd__nand2_1 _3745_ (.A(_0614_),
    .B(_0573_),
    .Y(_0821_));
 sky130_fd_sc_hd__a21o_2 _3746_ (.A1(_0550_),
    .A2(_0820_),
    .B1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__a22o_1 _3747_ (.A1(_0574_),
    .A2(_0558_),
    .B1(_0822_),
    .B2(_0566_),
    .X(_0823_));
 sky130_fd_sc_hd__and3_2 _3748_ (.A(_0384_),
    .B(_0392_),
    .C(_0400_),
    .X(_0824_));
 sky130_fd_sc_hd__a22o_1 _3749_ (.A1(\cu.reg_file.reg_d[7] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[7] ),
    .X(_0825_));
 sky130_fd_sc_hd__a22o_1 _3750_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[15] ),
    .X(_0826_));
 sky130_fd_sc_hd__a211o_1 _3751_ (.A1(\cu.pc.pc_o[15] ),
    .A2(_0740_),
    .B1(_0825_),
    .C1(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__a221o_1 _3752_ (.A1(\cu.reg_file.reg_a[7] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[15] ),
    .C1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__a22oi_4 _3753_ (.A1(\cu.id.imm_i[15] ),
    .A2(_0739_),
    .B1(_0828_),
    .B2(_0653_),
    .Y(_0829_));
 sky130_fd_sc_hd__a22o_1 _3754_ (.A1(\cu.reg_file.reg_sp[15] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[7] ),
    .X(_0830_));
 sky130_fd_sc_hd__a22o_1 _3755_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[7] ),
    .X(_0831_));
 sky130_fd_sc_hd__a211oi_4 _3756_ (.A1(\cu.reg_file.reg_mem[15] ),
    .A2(_0640_),
    .B1(_0830_),
    .C1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__xnor2_4 _3757_ (.A(_0829_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__a22o_1 _3758_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[6] ),
    .X(_0834_));
 sky130_fd_sc_hd__a22o_1 _3759_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[14] ),
    .X(_0835_));
 sky130_fd_sc_hd__a211o_1 _3760_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_0740_),
    .B1(_0834_),
    .C1(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__a221o_1 _3761_ (.A1(\cu.reg_file.reg_a[6] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[14] ),
    .C1(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__a22oi_4 _3762_ (.A1(\cu.id.imm_i[14] ),
    .A2(_0739_),
    .B1(_0837_),
    .B2(_0653_),
    .Y(_0838_));
 sky130_fd_sc_hd__a22o_1 _3763_ (.A1(\cu.reg_file.reg_sp[14] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[6] ),
    .X(_0839_));
 sky130_fd_sc_hd__a22o_1 _3764_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[6] ),
    .X(_0840_));
 sky130_fd_sc_hd__a211oi_2 _3765_ (.A1(\cu.reg_file.reg_mem[14] ),
    .A2(_0640_),
    .B1(_0839_),
    .C1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__and2b_1 _3766_ (.A_N(_0838_),
    .B(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__or2b_1 _3767_ (.A(_0841_),
    .B_N(_0838_),
    .X(_0843_));
 sky130_fd_sc_hd__and2b_1 _3768_ (.A_N(_0842_),
    .B(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__inv_2 _3769_ (.A(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__a22o_1 _3770_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[5] ),
    .X(_0846_));
 sky130_fd_sc_hd__a22o_1 _3771_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[13] ),
    .X(_0847_));
 sky130_fd_sc_hd__a211o_1 _3772_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_0740_),
    .B1(_0846_),
    .C1(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__a221o_1 _3773_ (.A1(\cu.reg_file.reg_a[5] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[13] ),
    .C1(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__a22oi_4 _3774_ (.A1(\cu.id.imm_i[13] ),
    .A2(_0739_),
    .B1(_0849_),
    .B2(_0653_),
    .Y(_0850_));
 sky130_fd_sc_hd__a22o_1 _3775_ (.A1(\cu.reg_file.reg_sp[13] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[5] ),
    .X(_0851_));
 sky130_fd_sc_hd__a22o_1 _3776_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[5] ),
    .X(_0852_));
 sky130_fd_sc_hd__a211oi_2 _3777_ (.A1(\cu.reg_file.reg_mem[13] ),
    .A2(_0640_),
    .B1(_0851_),
    .C1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__or2b_1 _3778_ (.A(_0850_),
    .B_N(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__or2b_1 _3779_ (.A(_0853_),
    .B_N(_0850_),
    .X(_0855_));
 sky130_fd_sc_hd__nand2_2 _3780_ (.A(_0854_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a22o_1 _3781_ (.A1(\cu.reg_file.reg_d[4] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[4] ),
    .X(_0857_));
 sky130_fd_sc_hd__a22o_1 _3782_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[12] ),
    .X(_0858_));
 sky130_fd_sc_hd__a211o_1 _3783_ (.A1(\cu.pc.pc_o[12] ),
    .A2(_0740_),
    .B1(_0857_),
    .C1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__a221o_1 _3784_ (.A1(\cu.reg_file.reg_a[4] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[12] ),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a22oi_4 _3785_ (.A1(\cu.id.imm_i[12] ),
    .A2(_0739_),
    .B1(_0860_),
    .B2(_0653_),
    .Y(_0861_));
 sky130_fd_sc_hd__a22o_1 _3786_ (.A1(\cu.reg_file.reg_sp[12] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[4] ),
    .X(_0862_));
 sky130_fd_sc_hd__a22o_1 _3787_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[4] ),
    .X(_0863_));
 sky130_fd_sc_hd__a211oi_2 _3788_ (.A1(\cu.reg_file.reg_mem[12] ),
    .A2(_0640_),
    .B1(_0862_),
    .C1(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__xnor2_1 _3789_ (.A(_0861_),
    .B(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__inv_2 _3790_ (.A(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__a22o_1 _3791_ (.A1(\cu.reg_file.reg_b[3] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[11] ),
    .X(_0867_));
 sky130_fd_sc_hd__a221o_1 _3792_ (.A1(\cu.reg_file.reg_d[3] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[3] ),
    .C1(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__a21o_1 _3793_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_0740_),
    .B1(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__a221o_1 _3794_ (.A1(\cu.reg_file.reg_a[3] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[11] ),
    .C1(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__a22oi_4 _3795_ (.A1(\cu.id.imm_i[11] ),
    .A2(_0739_),
    .B1(_0870_),
    .B2(_0653_),
    .Y(_0871_));
 sky130_fd_sc_hd__a22o_1 _3796_ (.A1(\cu.reg_file.reg_sp[11] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[3] ),
    .X(_0872_));
 sky130_fd_sc_hd__a22o_1 _3797_ (.A1(\cu.reg_file.reg_b[3] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[3] ),
    .X(_0873_));
 sky130_fd_sc_hd__a211oi_2 _3798_ (.A1(\cu.reg_file.reg_mem[11] ),
    .A2(_0640_),
    .B1(_0872_),
    .C1(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__and2b_1 _3799_ (.A_N(_0871_),
    .B(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__and2b_1 _3800_ (.A_N(_0874_),
    .B(_0871_),
    .X(_0876_));
 sky130_fd_sc_hd__or2_1 _3801_ (.A(_0875_),
    .B(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _3802_ (.A1(\cu.reg_file.reg_d[2] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[2] ),
    .X(_0878_));
 sky130_fd_sc_hd__a22o_1 _3803_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[10] ),
    .X(_0879_));
 sky130_fd_sc_hd__a211o_1 _3804_ (.A1(\cu.pc.pc_o[10] ),
    .A2(_0740_),
    .B1(_0878_),
    .C1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__a221o_1 _3805_ (.A1(\cu.reg_file.reg_a[2] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[10] ),
    .C1(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__a22o_2 _3806_ (.A1(\cu.id.imm_i[10] ),
    .A2(_0739_),
    .B1(_0881_),
    .B2(_0653_),
    .X(_0882_));
 sky130_fd_sc_hd__a22o_1 _3807_ (.A1(\cu.reg_file.reg_sp[10] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[2] ),
    .X(_0883_));
 sky130_fd_sc_hd__a22o_1 _3808_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[2] ),
    .X(_0884_));
 sky130_fd_sc_hd__a211oi_4 _3809_ (.A1(\cu.reg_file.reg_mem[10] ),
    .A2(_0640_),
    .B1(_0883_),
    .C1(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__xor2_1 _3810_ (.A(_0882_),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__inv_2 _3811_ (.A(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__a22o_1 _3812_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_0743_),
    .B1(_0624_),
    .B2(\cu.reg_file.reg_sp[9] ),
    .X(_0888_));
 sky130_fd_sc_hd__a221o_1 _3813_ (.A1(\cu.reg_file.reg_d[1] ),
    .A2(_0488_),
    .B1(_0741_),
    .B2(\cu.reg_file.reg_h[1] ),
    .C1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__a21o_1 _3814_ (.A1(\cu.pc.pc_o[9] ),
    .A2(_0740_),
    .B1(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__a221o_1 _3815_ (.A1(\cu.reg_file.reg_a[1] ),
    .A2(_0625_),
    .B1(_0628_),
    .B2(\cu.reg_file.reg_mem[9] ),
    .C1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__a22oi_4 _3816_ (.A1(\cu.id.imm_i[9] ),
    .A2(_0739_),
    .B1(_0891_),
    .B2(_0653_),
    .Y(_0892_));
 sky130_fd_sc_hd__a22o_1 _3817_ (.A1(\cu.reg_file.reg_sp[9] ),
    .A2(_0636_),
    .B1(_0748_),
    .B2(\cu.reg_file.reg_h[1] ),
    .X(_0893_));
 sky130_fd_sc_hd__a22o_1 _3818_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_0426_),
    .B1(_0429_),
    .B2(\cu.reg_file.reg_d[1] ),
    .X(_0894_));
 sky130_fd_sc_hd__a211oi_4 _3819_ (.A1(\cu.reg_file.reg_mem[9] ),
    .A2(_0640_),
    .B1(_0893_),
    .C1(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2b_1 _3820_ (.A(_0892_),
    .B_N(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__or2b_1 _3821_ (.A(_0895_),
    .B_N(_0892_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_2 _3822_ (.A(_0896_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__nor2_1 _3823_ (.A(_0747_),
    .B(_0751_),
    .Y(_0899_));
 sky130_fd_sc_hd__a2bb2o_1 _3824_ (.A1_N(_0892_),
    .A2_N(_0895_),
    .B1(_0898_),
    .B2(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__a31o_1 _3825_ (.A1(_0737_),
    .A2(_0752_),
    .A3(_0898_),
    .B1(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__inv_2 _3826_ (.A(_0882_),
    .Y(_0902_));
 sky130_fd_sc_hd__nor2_1 _3827_ (.A(_0902_),
    .B(_0885_),
    .Y(_0903_));
 sky130_fd_sc_hd__a21o_1 _3828_ (.A1(_0887_),
    .A2(_0901_),
    .B1(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__nor2_1 _3829_ (.A(_0871_),
    .B(_0874_),
    .Y(_0905_));
 sky130_fd_sc_hd__a21o_1 _3830_ (.A1(_0877_),
    .A2(_0904_),
    .B1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__nor2_1 _3831_ (.A(_0861_),
    .B(_0864_),
    .Y(_0907_));
 sky130_fd_sc_hd__a21o_1 _3832_ (.A1(_0866_),
    .A2(_0906_),
    .B1(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__nor2_1 _3833_ (.A(_0850_),
    .B(_0853_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21o_1 _3834_ (.A1(_0856_),
    .A2(_0908_),
    .B1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__nor2_1 _3835_ (.A(_0838_),
    .B(_0841_),
    .Y(_0911_));
 sky130_fd_sc_hd__a21oi_1 _3836_ (.A1(_0845_),
    .A2(_0910_),
    .B1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__or2_1 _3837_ (.A(_0829_),
    .B(_0832_),
    .X(_0913_));
 sky130_fd_sc_hd__o21a_1 _3838_ (.A1(_0833_),
    .A2(_0912_),
    .B1(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__nand2_1 _3839_ (.A(_0777_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__and2_2 _3840_ (.A(_0774_),
    .B(_0775_),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _3841_ (.A(_0401_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__buf_2 _3842_ (.A(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__inv_2 _3843_ (.A(_0832_),
    .Y(_0919_));
 sky130_fd_sc_hd__or2b_1 _3844_ (.A(_0747_),
    .B_N(_0751_),
    .X(_0920_));
 sky130_fd_sc_hd__and2b_1 _3845_ (.A_N(_0895_),
    .B(_0892_),
    .X(_0921_));
 sky130_fd_sc_hd__a31o_1 _3846_ (.A1(_0920_),
    .A2(_0896_),
    .A3(_0796_),
    .B1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__or2_1 _3847_ (.A(_0887_),
    .B(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__a21boi_1 _3848_ (.A1(_0882_),
    .A2(_0885_),
    .B1_N(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__o21ba_1 _3849_ (.A1(_0876_),
    .A2(_0924_),
    .B1_N(_0875_),
    .X(_0925_));
 sky130_fd_sc_hd__or2b_1 _3850_ (.A(_0861_),
    .B_N(_0864_),
    .X(_0926_));
 sky130_fd_sc_hd__o21a_1 _3851_ (.A1(_0866_),
    .A2(_0925_),
    .B1(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__and2b_1 _3852_ (.A_N(_0853_),
    .B(_0850_),
    .X(_0928_));
 sky130_fd_sc_hd__a21oi_2 _3853_ (.A1(_0854_),
    .A2(_0927_),
    .B1(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__o21ai_2 _3854_ (.A1(_0842_),
    .A2(_0929_),
    .B1(_0843_),
    .Y(_0930_));
 sky130_fd_sc_hd__o21a_1 _3855_ (.A1(_0829_),
    .A2(_0919_),
    .B1(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__a21o_1 _3856_ (.A1(_0829_),
    .A2(_0919_),
    .B1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__xnor2_1 _3857_ (.A(_0865_),
    .B(_0925_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_0920_),
    .B(_0796_),
    .Y(_0934_));
 sky130_fd_sc_hd__xor2_2 _3859_ (.A(_0898_),
    .B(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__or2b_1 _3860_ (.A(_0813_),
    .B_N(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__nand2_1 _3861_ (.A(_0887_),
    .B(_0922_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _3862_ (.A(_0923_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__and2b_1 _3863_ (.A_N(_0936_),
    .B(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__xnor2_1 _3864_ (.A(_0877_),
    .B(_0924_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand2_1 _3865_ (.A(_0939_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__nor2_1 _3866_ (.A(_0933_),
    .B(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__xnor2_2 _3867_ (.A(_0856_),
    .B(_0927_),
    .Y(_0943_));
 sky130_fd_sc_hd__xnor2_1 _3868_ (.A(_0844_),
    .B(_0929_),
    .Y(_0944_));
 sky130_fd_sc_hd__and3_1 _3869_ (.A(_0942_),
    .B(_0943_),
    .C(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__xor2_2 _3870_ (.A(_0833_),
    .B(_0930_),
    .X(_0946_));
 sky130_fd_sc_hd__and3_1 _3871_ (.A(_0817_),
    .B(_0945_),
    .C(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__xor2_1 _3872_ (.A(_0833_),
    .B(_0912_),
    .X(_0948_));
 sky130_fd_sc_hd__xnor2_1 _3873_ (.A(_0845_),
    .B(_0910_),
    .Y(_0949_));
 sky130_fd_sc_hd__xnor2_1 _3874_ (.A(_0856_),
    .B(_0908_),
    .Y(_0950_));
 sky130_fd_sc_hd__xnor2_1 _3875_ (.A(_0877_),
    .B(_0904_),
    .Y(_0951_));
 sky130_fd_sc_hd__xnor2_1 _3876_ (.A(_0887_),
    .B(_0901_),
    .Y(_0952_));
 sky130_fd_sc_hd__a21oi_1 _3877_ (.A1(_0737_),
    .A2(_0752_),
    .B1(_0899_),
    .Y(_0953_));
 sky130_fd_sc_hd__xnor2_1 _3878_ (.A(_0898_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__or2b_1 _3879_ (.A(_0771_),
    .B_N(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__or3_1 _3880_ (.A(_0951_),
    .B(_0952_),
    .C(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__xnor2_1 _3881_ (.A(_0866_),
    .B(_0906_),
    .Y(_0957_));
 sky130_fd_sc_hd__or3_1 _3882_ (.A(_0950_),
    .B(_0956_),
    .C(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__nor2_1 _3883_ (.A(_0949_),
    .B(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__nand2_1 _3884_ (.A(_0948_),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__o2bb2a_1 _3885_ (.A1_N(_0914_),
    .A2_N(_0960_),
    .B1(_0773_),
    .B2(_0777_),
    .X(_0961_));
 sky130_fd_sc_hd__a311o_1 _3886_ (.A1(_0918_),
    .A2(_0779_),
    .A3(_0932_),
    .B1(_0947_),
    .C1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__and3_1 _3887_ (.A(_0824_),
    .B(_0915_),
    .C(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__a211o_1 _3888_ (.A1(_0620_),
    .A2(_0819_),
    .B1(_0823_),
    .C1(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__nor2_1 _3889_ (.A(_2897_),
    .B(_0324_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _3890_ (.A(_2917_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__o221a_1 _3891_ (.A1(_2883_),
    .A2(_0304_),
    .B1(_0966_),
    .B2(_2893_),
    .C1(_0301_),
    .X(_0967_));
 sky130_fd_sc_hd__or2_2 _3892_ (.A(_0379_),
    .B(net150),
    .X(_0968_));
 sky130_fd_sc_hd__a211oi_1 _3893_ (.A1(_2893_),
    .A2(_0386_),
    .B1(_0308_),
    .C1(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__a21oi_1 _3894_ (.A1(_0967_),
    .A2(_0969_),
    .B1(_0328_),
    .Y(_0970_));
 sky130_fd_sc_hd__o22a_1 _3895_ (.A1(_2893_),
    .A2(_2896_),
    .B1(_2912_),
    .B2(_2923_),
    .X(_0971_));
 sky130_fd_sc_hd__nand2_1 _3896_ (.A(_2935_),
    .B(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__and2_1 _3897_ (.A(_2885_),
    .B(_2886_),
    .X(_0973_));
 sky130_fd_sc_hd__inv_2 _3898_ (.A(_0520_),
    .Y(_0974_));
 sky130_fd_sc_hd__a221o_1 _3899_ (.A1(_0359_),
    .A2(_0973_),
    .B1(_0364_),
    .B2(_0974_),
    .C1(_0296_),
    .X(_0975_));
 sky130_fd_sc_hd__or4_4 _3900_ (.A(_0321_),
    .B(_0970_),
    .C(_0972_),
    .D(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__nor2_1 _3901_ (.A(_0361_),
    .B(_0332_),
    .Y(_0977_));
 sky130_fd_sc_hd__a22oi_1 _3902_ (.A1(_2886_),
    .A2(_0965_),
    .B1(_0521_),
    .B2(_0359_),
    .Y(_0978_));
 sky130_fd_sc_hd__and4b_1 _3903_ (.A_N(_0308_),
    .B(_0525_),
    .C(_0977_),
    .D(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__and4b_2 _3904_ (.A_N(_0449_),
    .B(_0971_),
    .C(_0979_),
    .D(_2935_),
    .X(_0980_));
 sky130_fd_sc_hd__nor2_1 _3905_ (.A(_0350_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__nand2_1 _3906_ (.A(_0976_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__inv_2 _3907_ (.A(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_2918_),
    .B(_0966_),
    .Y(_0984_));
 sky130_fd_sc_hd__nor4_1 _3909_ (.A(_0310_),
    .B(_0328_),
    .C(_0740_),
    .D(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__nand2_4 _3910_ (.A(_0526_),
    .B(net145),
    .Y(_0986_));
 sky130_fd_sc_hd__nor3_1 _3911_ (.A(_0973_),
    .B(_0329_),
    .C(_0379_),
    .Y(_0987_));
 sky130_fd_sc_hd__o21a_1 _3912_ (.A1(_2936_),
    .A2(_2881_),
    .B1(_0469_),
    .X(_0988_));
 sky130_fd_sc_hd__a41o_2 _3913_ (.A1(_0966_),
    .A2(_0971_),
    .A3(_0987_),
    .A4(_0988_),
    .B1(_0296_),
    .X(_0989_));
 sky130_fd_sc_hd__a2111o_1 _3914_ (.A1(_2936_),
    .A2(_0386_),
    .B1(_0312_),
    .C1(_0323_),
    .D1(_0984_),
    .X(_0990_));
 sky130_fd_sc_hd__or2_1 _3915_ (.A(_0295_),
    .B(_0968_),
    .X(_0991_));
 sky130_fd_sc_hd__buf_2 _3916_ (.A(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_4 _3917_ (.A(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__or4_2 _3918_ (.A(_0449_),
    .B(_0972_),
    .C(_0990_),
    .D(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__nand3b_1 _3919_ (.A_N(_0986_),
    .B(_0989_),
    .C(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__inv_2 _3920_ (.A(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__or2_1 _3921_ (.A(_0989_),
    .B(_0994_),
    .X(_0997_));
 sky130_fd_sc_hd__nor2_1 _3922_ (.A(_0986_),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__inv_2 _3923_ (.A(_0980_),
    .Y(_0999_));
 sky130_fd_sc_hd__nor2_1 _3924_ (.A(_0976_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__nand2_1 _3925_ (.A(_0998_),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__nand2_1 _3926_ (.A(_0981_),
    .B(_0998_),
    .Y(_1002_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_1001_),
    .B(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__or2b_1 _3928_ (.A(_0994_),
    .B_N(_0989_),
    .X(_1004_));
 sky130_fd_sc_hd__or3_1 _3929_ (.A(_0976_),
    .B(_0980_),
    .C(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__o21ai_1 _3930_ (.A1(_0999_),
    .A2(_0997_),
    .B1(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__inv_2 _3931_ (.A(_0976_),
    .Y(_1007_));
 sky130_fd_sc_hd__and2b_1 _3932_ (.A_N(_1004_),
    .B(_0986_),
    .X(_1008_));
 sky130_fd_sc_hd__nor2_1 _3933_ (.A(_0998_),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__or3_1 _3934_ (.A(_1007_),
    .B(_0981_),
    .C(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__a21bo_1 _3935_ (.A1(_0986_),
    .A2(_1006_),
    .B1_N(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_2 _3936_ (.A(_0296_),
    .B(_2918_),
    .Y(_1012_));
 sky130_fd_sc_hd__and3_1 _3937_ (.A(_0372_),
    .B(_2921_),
    .C(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__o21a_1 _3938_ (.A1(\alu.Cin ),
    .A2(_1013_),
    .B1(_1012_),
    .X(_1014_));
 sky130_fd_sc_hd__a2111o_1 _3939_ (.A1(_0983_),
    .A2(_0996_),
    .B1(_1003_),
    .C1(_1011_),
    .D1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__and3_1 _3940_ (.A(_0976_),
    .B(_0981_),
    .C(_1008_),
    .X(_1016_));
 sky130_fd_sc_hd__and2b_1 _3941_ (.A_N(_1013_),
    .B(_1014_),
    .X(_1017_));
 sky130_fd_sc_hd__nand2_1 _3942_ (.A(_1000_),
    .B(_1008_),
    .Y(_1018_));
 sky130_fd_sc_hd__or2_2 _3943_ (.A(_0971_),
    .B(_0986_),
    .X(_1019_));
 sky130_fd_sc_hd__nand3_1 _3944_ (.A(_0531_),
    .B(_1018_),
    .C(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__nor3b_1 _3945_ (.A(_0982_),
    .B(_0997_),
    .C_N(_0986_),
    .Y(_1021_));
 sky130_fd_sc_hd__or4_1 _3946_ (.A(_1012_),
    .B(_0996_),
    .C(_1016_),
    .D(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__o41a_2 _3947_ (.A1(_1003_),
    .A2(_1011_),
    .A3(_1020_),
    .A4(_1022_),
    .B1(_2948_),
    .X(_1023_));
 sky130_fd_sc_hd__nor2_1 _3948_ (.A(_0572_),
    .B(_1020_),
    .Y(_1024_));
 sky130_fd_sc_hd__o2bb2a_1 _3949_ (.A1_N(_1023_),
    .A2_N(_1024_),
    .B1(\alu.Cin ),
    .B2(_1021_),
    .X(_1025_));
 sky130_fd_sc_hd__a2111o_1 _3950_ (.A1(_0964_),
    .A2(_1015_),
    .B1(_1016_),
    .C1(_1017_),
    .D1(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__nand2_4 _3951_ (.A(_2951_),
    .B(_0368_),
    .Y(_1027_));
 sky130_fd_sc_hd__o21a_1 _3952_ (.A1(\alu.Cin ),
    .A2(_1023_),
    .B1(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__a22o_1 _3953_ (.A1(_0370_),
    .A2(_0619_),
    .B1(_1026_),
    .B2(_1028_),
    .X(_0007_));
 sky130_fd_sc_hd__xor2_1 _3954_ (.A(_0712_),
    .B(_0713_),
    .X(_1029_));
 sky130_fd_sc_hd__inv_2 _3955_ (.A(_0511_),
    .Y(_1030_));
 sky130_fd_sc_hd__o21ai_1 _3956_ (.A1(_1030_),
    .A2(_1029_),
    .B1(_0773_),
    .Y(_1031_));
 sky130_fd_sc_hd__or2_4 _3957_ (.A(_0401_),
    .B(_0528_),
    .X(_1032_));
 sky130_fd_sc_hd__or2_1 _3958_ (.A(_1032_),
    .B(_0807_),
    .X(_1033_));
 sky130_fd_sc_hd__o211ai_1 _3959_ (.A1(_0758_),
    .A2(_1031_),
    .B1(_1033_),
    .C1(_0918_),
    .Y(_1034_));
 sky130_fd_sc_hd__or2_1 _3960_ (.A(_0781_),
    .B(_0712_),
    .X(_1035_));
 sky130_fd_sc_hd__a21oi_1 _3961_ (.A1(_0781_),
    .A2(_0712_),
    .B1(_0773_),
    .Y(_1036_));
 sky130_fd_sc_hd__o311a_1 _3962_ (.A1(_0572_),
    .A2(_0510_),
    .A3(_0401_),
    .B1(_1035_),
    .C1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__o22a_1 _3963_ (.A1(_0918_),
    .A2(_1029_),
    .B1(_1034_),
    .B2(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__nor2_1 _3964_ (.A(_0570_),
    .B(_0712_),
    .Y(_1039_));
 sky130_fd_sc_hd__inv_2 _3965_ (.A(_0710_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand2_1 _3966_ (.A(_0447_),
    .B(_0588_),
    .Y(_1041_));
 sky130_fd_sc_hd__nor2_1 _3967_ (.A(_0599_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__o22a_1 _3968_ (.A1(_0599_),
    .A2(_0603_),
    .B1(_0606_),
    .B2(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__inv_2 _3969_ (.A(_0611_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_1 _3970_ (.A(_0603_),
    .B(_0606_),
    .Y(_1045_));
 sky130_fd_sc_hd__o221ai_1 _3971_ (.A1(_0600_),
    .A2(_1044_),
    .B1(_1042_),
    .B2(_0610_),
    .C1(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__nor2_1 _3972_ (.A(_0531_),
    .B(_0545_),
    .Y(_1047_));
 sky130_fd_sc_hd__a221o_1 _3973_ (.A1(_0574_),
    .A2(_0822_),
    .B1(_1046_),
    .B2(_0545_),
    .C1(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__a211o_1 _3974_ (.A1(_0558_),
    .A2(_1040_),
    .B1(_1043_),
    .C1(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__a211o_4 _3975_ (.A1(_0517_),
    .A2(_1038_),
    .B1(_1039_),
    .C1(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__clkbuf_4 _3976_ (.A(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_8 _3977_ (.A(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__inv_2 _3978_ (.A(_1021_),
    .Y(_1053_));
 sky130_fd_sc_hd__o2111a_1 _3979_ (.A1(_0372_),
    .A2(_0371_),
    .B1(_0774_),
    .C1(_1019_),
    .D1(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nor2_1 _3980_ (.A(_0395_),
    .B(_1019_),
    .Y(_1055_));
 sky130_fd_sc_hd__o2bb2a_1 _3981_ (.A1_N(_1023_),
    .A2_N(_1054_),
    .B1(_1055_),
    .B2(\cu.alu_f[1] ),
    .X(_1056_));
 sky130_fd_sc_hd__o21ai_1 _3982_ (.A1(_0298_),
    .A2(_1001_),
    .B1(_1002_),
    .Y(_1057_));
 sky130_fd_sc_hd__o221a_1 _3983_ (.A1(\cu.alu_f[1] ),
    .A2(_1023_),
    .B1(_1056_),
    .B2(_1057_),
    .C1(_1027_),
    .X(_1058_));
 sky130_fd_sc_hd__a21o_1 _3984_ (.A1(_0370_),
    .A2(_1052_),
    .B1(_1058_),
    .X(_0008_));
 sky130_fd_sc_hd__inv_2 _3985_ (.A(_0603_),
    .Y(_1059_));
 sky130_fd_sc_hd__clkbuf_4 _3986_ (.A(_0575_),
    .X(_1060_));
 sky130_fd_sc_hd__and3_1 _3987_ (.A(_1060_),
    .B(_0588_),
    .C(_0599_),
    .X(_1061_));
 sky130_fd_sc_hd__o2bb2a_1 _3988_ (.A1_N(_0588_),
    .A2_N(_1059_),
    .B1(_0606_),
    .B2(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__a221o_1 _3989_ (.A1(_0558_),
    .A2(_0694_),
    .B1(_0822_),
    .B2(_0545_),
    .C1(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__a21oi_1 _3990_ (.A1(_0761_),
    .A2(_0772_),
    .B1(_0777_),
    .Y(_1064_));
 sky130_fd_sc_hd__o21bai_1 _3991_ (.A1(_0758_),
    .A2(_0760_),
    .B1_N(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__a21oi_1 _3992_ (.A1(_0816_),
    .A2(_0807_),
    .B1(_0776_),
    .Y(_1066_));
 sky130_fd_sc_hd__mux2_1 _3993_ (.A0(_1033_),
    .A1(_1066_),
    .S(_0806_),
    .X(_1067_));
 sky130_fd_sc_hd__a2bb2o_1 _3994_ (.A1_N(_0918_),
    .A2_N(_0760_),
    .B1(_1065_),
    .B2(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__nor2_1 _3995_ (.A(_0620_),
    .B(_0824_),
    .Y(_1069_));
 sky130_fd_sc_hd__o22a_1 _3996_ (.A1(_0570_),
    .A2(_0759_),
    .B1(_1068_),
    .B2(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__o221a_1 _3997_ (.A1(_0588_),
    .A2(_1044_),
    .B1(_1061_),
    .B2(_0610_),
    .C1(_1045_),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _3998_ (.A0(_0531_),
    .A1(_1071_),
    .S(_1040_),
    .X(_1072_));
 sky130_fd_sc_hd__nand3b_4 _3999_ (.A_N(_1063_),
    .B(_1070_),
    .C(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__buf_4 _4000_ (.A(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_8 _4001_ (.A(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__and3b_1 _4002_ (.A_N(_0761_),
    .B(_0764_),
    .C(_0772_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_1 _4003_ (.A(_0764_),
    .B(_1064_),
    .Y(_1077_));
 sky130_fd_sc_hd__nor2_1 _4004_ (.A(_0808_),
    .B(_0810_),
    .Y(_1078_));
 sky130_fd_sc_hd__a21o_1 _4005_ (.A1(_0817_),
    .A2(_0808_),
    .B1(_0776_),
    .X(_1079_));
 sky130_fd_sc_hd__a22o_1 _4006_ (.A1(_0817_),
    .A2(_1078_),
    .B1(_1079_),
    .B2(_0810_),
    .X(_1080_));
 sky130_fd_sc_hd__o31a_1 _4007_ (.A1(_1076_),
    .A2(_1077_),
    .A3(_1080_),
    .B1(_0517_),
    .X(_1081_));
 sky130_fd_sc_hd__nor2_1 _4008_ (.A(_0570_),
    .B(_0763_),
    .Y(_1082_));
 sky130_fd_sc_hd__nor2_1 _4009_ (.A(_0600_),
    .B(_1041_),
    .Y(_1083_));
 sky130_fd_sc_hd__nor2_1 _4010_ (.A(_0531_),
    .B(_0694_),
    .Y(_1084_));
 sky130_fd_sc_hd__a221o_1 _4011_ (.A1(_0606_),
    .A2(_0701_),
    .B1(_1083_),
    .B2(_0603_),
    .C1(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__a2bb2o_1 _4012_ (.A1_N(_0610_),
    .A2_N(_1083_),
    .B1(_0701_),
    .B2(_0611_),
    .X(_1086_));
 sky130_fd_sc_hd__o21a_1 _4013_ (.A1(_0607_),
    .A2(_1086_),
    .B1(_0694_),
    .X(_1087_));
 sky130_fd_sc_hd__a221o_1 _4014_ (.A1(_0558_),
    .A2(_0681_),
    .B1(_0822_),
    .B2(_1040_),
    .C1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__or4_4 _4015_ (.A(_1081_),
    .B(_1082_),
    .C(_1085_),
    .D(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__xnor2_1 _4016_ (.A(_1073_),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(_0770_),
    .B(_0773_),
    .Y(_1091_));
 sky130_fd_sc_hd__o2bb2a_1 _4018_ (.A1_N(_0776_),
    .A2_N(_0801_),
    .B1(_1091_),
    .B2(_0768_),
    .X(_1092_));
 sky130_fd_sc_hd__nor2_1 _4019_ (.A(_0801_),
    .B(_0812_),
    .Y(_1093_));
 sky130_fd_sc_hd__and2_1 _4020_ (.A(_0801_),
    .B(_0812_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _4021_ (.A(_1093_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _4022_ (.A(_0768_),
    .B(_0772_),
    .Y(_1096_));
 sky130_fd_sc_hd__and2_1 _4023_ (.A(_0918_),
    .B(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__o22a_1 _4024_ (.A1(_1032_),
    .A2(_1095_),
    .B1(_1097_),
    .B2(_0770_),
    .X(_1098_));
 sky130_fd_sc_hd__a21oi_1 _4025_ (.A1(_1092_),
    .A2(_1098_),
    .B1(_1069_),
    .Y(_1099_));
 sky130_fd_sc_hd__or2_1 _4026_ (.A(_1060_),
    .B(_0588_),
    .X(_1100_));
 sky130_fd_sc_hd__inv_2 _4027_ (.A(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__a21oi_1 _4028_ (.A1(_0599_),
    .A2(_1101_),
    .B1(_0610_),
    .Y(_1102_));
 sky130_fd_sc_hd__a211o_1 _4029_ (.A1(_0611_),
    .A2(_0729_),
    .B1(_0607_),
    .C1(_0552_),
    .X(_1103_));
 sky130_fd_sc_hd__a32o_1 _4030_ (.A1(_0599_),
    .A2(_0603_),
    .A3(_1101_),
    .B1(_0729_),
    .B2(_0606_),
    .X(_1104_));
 sky130_fd_sc_hd__o22a_1 _4031_ (.A1(_1102_),
    .A2(_1103_),
    .B1(_1104_),
    .B2(_0566_),
    .X(_1105_));
 sky130_fd_sc_hd__o2bb2a_1 _4032_ (.A1_N(\alu.Cin ),
    .A2_N(_0554_),
    .B1(_0556_),
    .B2(_0509_),
    .X(_1106_));
 sky130_fd_sc_hd__o2bb2a_1 _4033_ (.A1_N(_0822_),
    .A2_N(_0632_),
    .B1(_0566_),
    .B2(_0531_),
    .X(_1107_));
 sky130_fd_sc_hd__o211a_1 _4034_ (.A1(_0570_),
    .A2(_0733_),
    .B1(_1106_),
    .C1(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__or3b_1 _4035_ (.A(_1099_),
    .B(_1105_),
    .C_N(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__buf_4 _4036_ (.A(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__nand2_1 _4037_ (.A(_0611_),
    .B(_0643_),
    .Y(_1111_));
 sky130_fd_sc_hd__or2_1 _4038_ (.A(_0588_),
    .B(_0610_),
    .X(_1112_));
 sky130_fd_sc_hd__nand2_1 _4039_ (.A(_1060_),
    .B(_0599_),
    .Y(_1113_));
 sky130_fd_sc_hd__o2bb2a_1 _4040_ (.A1_N(_0610_),
    .A2_N(_1111_),
    .B1(_1112_),
    .B2(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__o21a_1 _4041_ (.A1(_0607_),
    .A2(_1114_),
    .B1(_0632_),
    .X(_1115_));
 sky130_fd_sc_hd__a2bb2o_1 _4042_ (.A1_N(_0531_),
    .A2_N(_0632_),
    .B1(_0566_),
    .B2(_0558_),
    .X(_1116_));
 sky130_fd_sc_hd__or2_1 _4043_ (.A(_0588_),
    .B(_1059_),
    .X(_1117_));
 sky130_fd_sc_hd__nor2_1 _4044_ (.A(_1113_),
    .B(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__a221o_1 _4045_ (.A1(_0606_),
    .A2(_0643_),
    .B1(_0663_),
    .B2(_0822_),
    .C1(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__or2_1 _4046_ (.A(_0757_),
    .B(_0767_),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_1 _4047_ (.A(_0804_),
    .B(_0811_),
    .Y(_1121_));
 sky130_fd_sc_hd__o21ai_1 _4048_ (.A1(_1032_),
    .A2(_1121_),
    .B1(_0916_),
    .Y(_1122_));
 sky130_fd_sc_hd__o2bb2a_1 _4049_ (.A1_N(_0802_),
    .A2_N(_1122_),
    .B1(_0812_),
    .B2(_1032_),
    .X(_1123_));
 sky130_fd_sc_hd__o221a_1 _4050_ (.A1(_1120_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_0754_),
    .C1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__o22a_1 _4051_ (.A1(_0570_),
    .A2(_0644_),
    .B1(_1124_),
    .B2(_1069_),
    .X(_1125_));
 sky130_fd_sc_hd__or4b_4 _4052_ (.A(_1115_),
    .B(_1116_),
    .C(_1119_),
    .D_N(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_1 _4053_ (.A(_1110_),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__and2_1 _4054_ (.A(_1110_),
    .B(_1126_),
    .X(_1128_));
 sky130_fd_sc_hd__nor2_1 _4055_ (.A(_1127_),
    .B(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__and2_1 _4056_ (.A(_0804_),
    .B(_0811_),
    .X(_1130_));
 sky130_fd_sc_hd__o21a_1 _4057_ (.A1(_1121_),
    .A2(_1130_),
    .B1(_0817_),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _4058_ (.A(_0757_),
    .B(_0767_),
    .Y(_1132_));
 sky130_fd_sc_hd__a2bb2o_1 _4059_ (.A1_N(_0917_),
    .A2_N(_0757_),
    .B1(_0804_),
    .B2(_0776_),
    .X(_1133_));
 sky130_fd_sc_hd__a31o_1 _4060_ (.A1(_1120_),
    .A2(_0773_),
    .A3(_1132_),
    .B1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__o21a_1 _4061_ (.A1(_1131_),
    .A2(_1134_),
    .B1(_0517_),
    .X(_1135_));
 sky130_fd_sc_hd__nor2_1 _4062_ (.A(_0599_),
    .B(_1100_),
    .Y(_1136_));
 sky130_fd_sc_hd__nand2_1 _4063_ (.A(_0603_),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__a21oi_1 _4064_ (.A1(_0719_),
    .A2(_1137_),
    .B1(_1045_),
    .Y(_1138_));
 sky130_fd_sc_hd__a2bb2o_1 _4065_ (.A1_N(_0610_),
    .A2_N(_1136_),
    .B1(_0652_),
    .B2(_0611_),
    .X(_1139_));
 sky130_fd_sc_hd__a2bb2o_1 _4066_ (.A1_N(_0531_),
    .A2_N(_0663_),
    .B1(_0681_),
    .B2(_0822_),
    .X(_1140_));
 sky130_fd_sc_hd__a221o_1 _4067_ (.A1(_0558_),
    .A2(_0632_),
    .B1(_0663_),
    .B2(_1139_),
    .C1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__nor2_1 _4068_ (.A(_0570_),
    .B(_0664_),
    .Y(_1142_));
 sky130_fd_sc_hd__or4_1 _4069_ (.A(_1135_),
    .B(_1138_),
    .C(_1141_),
    .D(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__buf_4 _4070_ (.A(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__or2_1 _4071_ (.A(_0765_),
    .B(_0766_),
    .X(_1145_));
 sky130_fd_sc_hd__o21ai_1 _4072_ (.A1(_0808_),
    .A2(_0810_),
    .B1(_0805_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _4073_ (.A(_0811_),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__a221o_1 _4074_ (.A1(_0776_),
    .A2(_0805_),
    .B1(_1147_),
    .B2(_0817_),
    .C1(_0777_),
    .X(_1148_));
 sky130_fd_sc_hd__a31o_1 _4075_ (.A1(_0767_),
    .A2(_0773_),
    .A3(_1145_),
    .B1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__o211a_1 _4076_ (.A1(_0918_),
    .A2(_0766_),
    .B1(_1149_),
    .C1(_0517_),
    .X(_1150_));
 sky130_fd_sc_hd__nor2_1 _4077_ (.A(_0570_),
    .B(_0684_),
    .Y(_1151_));
 sky130_fd_sc_hd__a22o_1 _4078_ (.A1(_0558_),
    .A2(_0663_),
    .B1(_0822_),
    .B2(_0694_),
    .X(_1152_));
 sky130_fd_sc_hd__nand2_1 _4079_ (.A(_1060_),
    .B(_0600_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_1 _4080_ (.A(_0611_),
    .B(_0671_),
    .Y(_1154_));
 sky130_fd_sc_hd__a2bb2o_1 _4081_ (.A1_N(_1153_),
    .A2_N(_1112_),
    .B1(_1154_),
    .B2(_0610_),
    .X(_1155_));
 sky130_fd_sc_hd__nor2_1 _4082_ (.A(_1153_),
    .B(_1117_),
    .Y(_1156_));
 sky130_fd_sc_hd__a211oi_1 _4083_ (.A1(_0606_),
    .A2(_0671_),
    .B1(_0681_),
    .C1(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__a32o_1 _4084_ (.A1(_1045_),
    .A2(_0681_),
    .A3(_1155_),
    .B1(_1157_),
    .B2(_0531_),
    .X(_1158_));
 sky130_fd_sc_hd__or4b_1 _4085_ (.A(_1150_),
    .B(_1151_),
    .C(_1152_),
    .D_N(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__buf_4 _4086_ (.A(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__xor2_1 _4087_ (.A(_1144_),
    .B(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__xor2_1 _4088_ (.A(_0617_),
    .B(_1050_),
    .X(_1162_));
 sky130_fd_sc_hd__xnor2_1 _4089_ (.A(_1161_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__xnor2_1 _4090_ (.A(_1129_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__inv_2 _4091_ (.A(_0820_),
    .Y(_1165_));
 sky130_fd_sc_hd__o211ai_1 _4092_ (.A1(_0519_),
    .A2(_1165_),
    .B1(_0614_),
    .C1(_0551_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _4093_ (.A(_1090_),
    .B(_1164_),
    .Y(_1167_));
 sky130_fd_sc_hd__o221a_1 _4094_ (.A1(_1090_),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0611_),
    .C1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__xnor2_1 _4095_ (.A(_0566_),
    .B(_1110_),
    .Y(_1169_));
 sky130_fd_sc_hd__xor2_1 _4096_ (.A(_0546_),
    .B(_0733_),
    .X(_1170_));
 sky130_fd_sc_hd__xor2_1 _4097_ (.A(_0945_),
    .B(_0946_),
    .X(_1171_));
 sky130_fd_sc_hd__o221a_1 _4098_ (.A1(_0916_),
    .A2(_0946_),
    .B1(_1171_),
    .B2(_1032_),
    .C1(_0918_),
    .X(_1172_));
 sky130_fd_sc_hd__o21a_1 _4099_ (.A1(_0948_),
    .A2(_0959_),
    .B1(_0773_),
    .X(_1173_));
 sky130_fd_sc_hd__nand2_1 _4100_ (.A(_0960_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__a2bb2o_2 _4101_ (.A1_N(_0918_),
    .A2_N(_0948_),
    .B1(_1172_),
    .B2(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__xnor2_1 _4102_ (.A(_0829_),
    .B(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__o21ai_1 _4103_ (.A1(_0547_),
    .A2(_0833_),
    .B1(_0824_),
    .Y(_1177_));
 sky130_fd_sc_hd__a211o_1 _4104_ (.A1(_0547_),
    .A2(_0833_),
    .B1(_1176_),
    .C1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__o31ai_1 _4105_ (.A1(_0395_),
    .A2(_1169_),
    .A3(_1170_),
    .B1(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__o21a_1 _4106_ (.A1(\cu.alu_f[2] ),
    .A2(_1013_),
    .B1(_1012_),
    .X(_1180_));
 sky130_fd_sc_hd__a21oi_1 _4107_ (.A1(_1018_),
    .A2(_1019_),
    .B1(_0395_),
    .Y(_1181_));
 sky130_fd_sc_hd__or4b_2 _4108_ (.A(_0996_),
    .B(_1003_),
    .C(_1181_),
    .D_N(_1010_),
    .X(_1182_));
 sky130_fd_sc_hd__o221a_1 _4109_ (.A1(_1168_),
    .A2(_1179_),
    .B1(_1180_),
    .B2(_1182_),
    .C1(_1023_),
    .X(_1183_));
 sky130_fd_sc_hd__o21ai_2 _4110_ (.A1(_1013_),
    .A2(_1182_),
    .B1(_1023_),
    .Y(_1184_));
 sky130_fd_sc_hd__a21o_1 _4111_ (.A1(\cu.alu_f[2] ),
    .A2(_1184_),
    .B1(_0370_),
    .X(_1185_));
 sky130_fd_sc_hd__o22a_1 _4112_ (.A1(_1027_),
    .A2(_1075_),
    .B1(_1183_),
    .B2(_1185_),
    .X(_0009_));
 sky130_fd_sc_hd__or2_2 _4113_ (.A(_2946_),
    .B(_2947_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_4 _4114_ (.A(_1089_),
    .X(_1187_));
 sky130_fd_sc_hd__buf_4 _4115_ (.A(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__a22o_1 _4116_ (.A1(net209),
    .A2(_1186_),
    .B1(_0370_),
    .B2(_1188_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_4 _4117_ (.A(_1160_),
    .X(_1189_));
 sky130_fd_sc_hd__buf_4 _4118_ (.A(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__a22o_1 _4119_ (.A1(net212),
    .A2(_1186_),
    .B1(_0370_),
    .B2(_1190_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_4 _4120_ (.A(_1144_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_8 _4121_ (.A(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__a22o_1 _4122_ (.A1(net208),
    .A2(_1186_),
    .B1(_0370_),
    .B2(_1192_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_4 _4123_ (.A(_1126_),
    .X(_1193_));
 sky130_fd_sc_hd__buf_4 _4124_ (.A(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__a21oi_1 _4125_ (.A1(_0942_),
    .A2(_0943_),
    .B1(_0944_),
    .Y(_1195_));
 sky130_fd_sc_hd__nor2_1 _4126_ (.A(_0945_),
    .B(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__o221a_1 _4127_ (.A1(_0916_),
    .A2(_0944_),
    .B1(_1196_),
    .B2(_1032_),
    .C1(_0918_),
    .X(_1197_));
 sky130_fd_sc_hd__a21o_1 _4128_ (.A1(_0949_),
    .A2(_0958_),
    .B1(_0779_),
    .X(_1198_));
 sky130_fd_sc_hd__or2_1 _4129_ (.A(_0959_),
    .B(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__a22o_1 _4130_ (.A1(_0777_),
    .A2(_0949_),
    .B1(_1197_),
    .B2(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__nand2_1 _4131_ (.A(_0942_),
    .B(_0943_),
    .Y(_1201_));
 sky130_fd_sc_hd__or2_1 _4132_ (.A(_0942_),
    .B(_0943_),
    .X(_1202_));
 sky130_fd_sc_hd__a21o_1 _4133_ (.A1(_1201_),
    .A2(_1202_),
    .B1(_1032_),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_1 _4134_ (.A(_0956_),
    .B(_0957_),
    .Y(_1204_));
 sky130_fd_sc_hd__or2_1 _4135_ (.A(_1204_),
    .B(_0779_),
    .X(_1205_));
 sky130_fd_sc_hd__and2_1 _4136_ (.A(_0918_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__nand3_1 _4137_ (.A(_0950_),
    .B(_1204_),
    .C(_0773_),
    .Y(_1207_));
 sky130_fd_sc_hd__o221a_1 _4138_ (.A1(_0916_),
    .A2(_0943_),
    .B1(_1206_),
    .B2(_0950_),
    .C1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__a21oi_4 _4139_ (.A1(_1203_),
    .A2(_1208_),
    .B1(_0516_),
    .Y(_1209_));
 sky130_fd_sc_hd__a21o_1 _4140_ (.A1(_0817_),
    .A2(_0941_),
    .B1(_0776_),
    .X(_1210_));
 sky130_fd_sc_hd__a22oi_1 _4141_ (.A1(_0817_),
    .A2(_0942_),
    .B1(_1210_),
    .B2(_0933_),
    .Y(_1211_));
 sky130_fd_sc_hd__o221a_1 _4142_ (.A1(_0956_),
    .A2(_1205_),
    .B1(_1206_),
    .B2(_0957_),
    .C1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__nor2_4 _4143_ (.A(_0516_),
    .B(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__nor2_1 _4144_ (.A(_0952_),
    .B(_0955_),
    .Y(_1214_));
 sky130_fd_sc_hd__or2_1 _4145_ (.A(_1214_),
    .B(_0779_),
    .X(_1215_));
 sky130_fd_sc_hd__and2_1 _4146_ (.A(_0917_),
    .B(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__nor2_1 _4147_ (.A(_0951_),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__or2_1 _4148_ (.A(_0939_),
    .B(_0940_),
    .X(_1218_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(_0941_),
    .B(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__a2bb2o_1 _4150_ (.A1_N(_0916_),
    .A2_N(_0940_),
    .B1(_1219_),
    .B2(_0817_),
    .X(_1220_));
 sky130_fd_sc_hd__a31o_1 _4151_ (.A1(_0951_),
    .A2(_1214_),
    .A3(_0773_),
    .B1(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__o21a_4 _4152_ (.A1(_1217_),
    .A2(_1221_),
    .B1(_0824_),
    .X(_1222_));
 sky130_fd_sc_hd__a21oi_1 _4153_ (.A1(_0816_),
    .A2(_0936_),
    .B1(_0776_),
    .Y(_1223_));
 sky130_fd_sc_hd__o2bb2a_1 _4154_ (.A1_N(_0817_),
    .A2_N(_0939_),
    .B1(_1223_),
    .B2(_0938_),
    .X(_1224_));
 sky130_fd_sc_hd__o221a_1 _4155_ (.A1(_0955_),
    .A2(_1215_),
    .B1(_1216_),
    .B2(_0952_),
    .C1(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__nor2_4 _4156_ (.A(_0516_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__xnor2_1 _4157_ (.A(_0935_),
    .B(_0813_),
    .Y(_1227_));
 sky130_fd_sc_hd__o32a_1 _4158_ (.A1(_0771_),
    .A2(_0954_),
    .A3(_0779_),
    .B1(_0935_),
    .B2(_0916_),
    .X(_1228_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(_0954_),
    .B(_0778_),
    .Y(_1229_));
 sky130_fd_sc_hd__o211a_2 _4160_ (.A1(_1032_),
    .A2(_1227_),
    .B1(_1228_),
    .C1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__or4b_1 _4161_ (.A(_0516_),
    .B(_0819_),
    .C(_1226_),
    .D_N(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__nor4_1 _4162_ (.A(_1209_),
    .B(_1213_),
    .C(_1222_),
    .D(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__buf_4 _4163_ (.A(_2920_),
    .X(_1233_));
 sky130_fd_sc_hd__nor2_1 _4164_ (.A(_1233_),
    .B(_0371_),
    .Y(_1234_));
 sky130_fd_sc_hd__a21oi_1 _4165_ (.A1(_0387_),
    .A2(_1234_),
    .B1(_0824_),
    .Y(_1235_));
 sky130_fd_sc_hd__a31o_1 _4166_ (.A1(_1175_),
    .A2(_1200_),
    .A3(_1232_),
    .B1(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__or4_1 _4167_ (.A(_0617_),
    .B(_1050_),
    .C(_1073_),
    .D(_1089_),
    .X(_1237_));
 sky130_fd_sc_hd__nor3_1 _4168_ (.A(_1144_),
    .B(_1160_),
    .C(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__mux2_1 _4169_ (.A0(_0829_),
    .A1(_0838_),
    .S(_1060_),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(_0850_),
    .A1(_0861_),
    .S(_1060_),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(_1239_),
    .A1(_1240_),
    .S(_0600_),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _4172_ (.A0(_0871_),
    .A1(_0902_),
    .S(_1060_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _4173_ (.A0(_0747_),
    .A1(_0892_),
    .S(_0447_),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _4174_ (.A0(_1242_),
    .A1(_1243_),
    .S(_0600_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(_1241_),
    .A1(_1244_),
    .S(_0588_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(_0566_),
    .A1(_0632_),
    .S(_1060_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(_0663_),
    .A1(_0681_),
    .S(_1060_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _4178_ (.A0(_1246_),
    .A1(_1247_),
    .S(_0600_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _4179_ (.A0(_0574_),
    .A1(_0545_),
    .S(_0447_),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(_0694_),
    .A1(_1040_),
    .S(_1060_),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(_1249_),
    .A1(_1250_),
    .S(_0599_),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(_1248_),
    .A1(_1251_),
    .S(_0588_),
    .X(_1252_));
 sky130_fd_sc_hd__nor2_1 _4183_ (.A(_0701_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__a21o_1 _4184_ (.A1(_0701_),
    .A2(_1245_),
    .B1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__and3_1 _4185_ (.A(_0387_),
    .B(_1234_),
    .C(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__a31o_2 _4186_ (.A1(_1127_),
    .A2(_1236_),
    .A3(_1238_),
    .B1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__o21a_1 _4187_ (.A1(_1234_),
    .A2(_1182_),
    .B1(_1023_),
    .X(_1257_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(\cu.alu_f[6] ),
    .A1(_1256_),
    .S(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(_1194_),
    .A1(_1258_),
    .S(_1027_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _4190_ (.A(_1259_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_4 _4191_ (.A(_1110_),
    .X(_1260_));
 sky130_fd_sc_hd__buf_4 _4192_ (.A(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__inv_2 _4193_ (.A(_1184_),
    .Y(_1262_));
 sky130_fd_sc_hd__nor2_4 _4194_ (.A(_0516_),
    .B(_1175_),
    .Y(_1263_));
 sky130_fd_sc_hd__a22o_1 _4195_ (.A1(_0516_),
    .A2(_1260_),
    .B1(_1263_),
    .B2(_1027_),
    .X(_1264_));
 sky130_fd_sc_hd__and3_1 _4196_ (.A(\cu.alu_f[7] ),
    .B(_1027_),
    .C(_1184_),
    .X(_1265_));
 sky130_fd_sc_hd__a221o_1 _4197_ (.A1(_0370_),
    .A2(_1261_),
    .B1(_1262_),
    .B2(_1264_),
    .C1(_1265_),
    .X(_0014_));
 sky130_fd_sc_hd__and3_1 _4198_ (.A(_2877_),
    .B(_0436_),
    .C(_0469_),
    .X(_1266_));
 sky130_fd_sc_hd__o211a_1 _4199_ (.A1(_0323_),
    .A2(_1266_),
    .B1(_2912_),
    .C1(_2937_),
    .X(_1267_));
 sky130_fd_sc_hd__buf_2 _4200_ (.A(\cu.id.state[2] ),
    .X(_1268_));
 sky130_fd_sc_hd__and3b_2 _4201_ (.A_N(\cu.id.state[1] ),
    .B(\cu.id.state[0] ),
    .C(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__or3b_2 _4202_ (.A(_0294_),
    .B(_1267_),
    .C_N(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__buf_2 _4203_ (.A(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__inv_2 _4204_ (.A(_0469_),
    .Y(_1272_));
 sky130_fd_sc_hd__or2_1 _4205_ (.A(_0359_),
    .B(_2937_),
    .X(_1273_));
 sky130_fd_sc_hd__a21o_1 _4206_ (.A1(_0336_),
    .A2(_1266_),
    .B1(_0293_),
    .X(_1274_));
 sky130_fd_sc_hd__a31o_1 _4207_ (.A1(_2912_),
    .A2(_0583_),
    .A3(_1273_),
    .B1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__a31o_2 _4208_ (.A1(_2912_),
    .A2(_2937_),
    .A3(_0583_),
    .B1(_1274_),
    .X(_1276_));
 sky130_fd_sc_hd__or2_1 _4209_ (.A(_2883_),
    .B(_2937_),
    .X(_1277_));
 sky130_fd_sc_hd__a31o_1 _4210_ (.A1(_2877_),
    .A2(_0336_),
    .A3(_0436_),
    .B1(_0293_),
    .X(_1278_));
 sky130_fd_sc_hd__a31o_2 _4211_ (.A1(_2912_),
    .A2(_0583_),
    .A3(_1277_),
    .B1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__nor4b_1 _4212_ (.A(_1272_),
    .B(_1275_),
    .C(_1276_),
    .D_N(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__buf_2 _4213_ (.A(net238),
    .X(_1281_));
 sky130_fd_sc_hd__nor2b_4 _4214_ (.A(_1279_),
    .B_N(_1275_),
    .Y(_1282_));
 sky130_fd_sc_hd__buf_2 _4215_ (.A(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__nor2_4 _4216_ (.A(_1279_),
    .B(_1275_),
    .Y(_1284_));
 sky130_fd_sc_hd__buf_2 _4217_ (.A(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__nor2_4 _4218_ (.A(_0295_),
    .B(_0469_),
    .Y(_1286_));
 sky130_fd_sc_hd__buf_2 _4219_ (.A(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__a22o_1 _4220_ (.A1(\cu.reg_file.reg_a[0] ),
    .A2(_1276_),
    .B1(_1287_),
    .B2(\cu.reg_file.reg_sp[0] ),
    .X(_1288_));
 sky130_fd_sc_hd__a221o_1 _4221_ (.A1(\cu.reg_file.reg_e[0] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[0] ),
    .C1(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__a21oi_1 _4222_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_1281_),
    .B1(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__nor2_1 _4223_ (.A(_1271_),
    .B(_1290_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2_1 _4224_ (.A(_2904_),
    .B(_2924_),
    .Y(_1292_));
 sky130_fd_sc_hd__and3_2 _4225_ (.A(_2950_),
    .B(_1292_),
    .C(_1269_),
    .X(_1293_));
 sky130_fd_sc_hd__buf_2 _4226_ (.A(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__buf_2 _4227_ (.A(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__inv_2 _4228_ (.A(_1271_),
    .Y(_1296_));
 sky130_fd_sc_hd__nor2_2 _4229_ (.A(_1296_),
    .B(_1294_),
    .Y(_1297_));
 sky130_fd_sc_hd__buf_2 _4230_ (.A(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_4 _4231_ (.A(\cu.pc.pc_o[0] ),
    .X(_1299_));
 sky130_fd_sc_hd__buf_2 _4232_ (.A(\cu.id.state[0] ),
    .X(_1300_));
 sky130_fd_sc_hd__buf_2 _4233_ (.A(\cu.id.state[1] ),
    .X(_1301_));
 sky130_fd_sc_hd__and2b_1 _4234_ (.A_N(_1300_),
    .B(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__inv_2 _4235_ (.A(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__nor2_2 _4236_ (.A(_2946_),
    .B(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__clkbuf_8 _4237_ (.A(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_4 _4238_ (.A(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__a221o_1 _4239_ (.A1(_0343_),
    .A2(_1295_),
    .B1(_1298_),
    .B2(_1299_),
    .C1(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__a211oi_1 _4240_ (.A1(_0359_),
    .A2(_0320_),
    .B1(_0336_),
    .C1(_2914_),
    .Y(_1308_));
 sky130_fd_sc_hd__a211o_2 _4241_ (.A1(_0336_),
    .A2(_0436_),
    .B1(_1308_),
    .C1(_0295_),
    .X(_1309_));
 sky130_fd_sc_hd__o31a_1 _4242_ (.A1(_2908_),
    .A2(_0361_),
    .A3(_0968_),
    .B1(_0336_),
    .X(_1310_));
 sky130_fd_sc_hd__a2111o_2 _4243_ (.A1(_2883_),
    .A2(_0320_),
    .B1(_1310_),
    .C1(_0295_),
    .D1(_2914_),
    .X(_1311_));
 sky130_fd_sc_hd__and3b_2 _4244_ (.A_N(_0992_),
    .B(_1309_),
    .C(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_4 _4245_ (.A(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__nor2_2 _4246_ (.A(_1309_),
    .B(_1311_),
    .Y(_1314_));
 sky130_fd_sc_hd__buf_2 _4247_ (.A(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__nor2b_2 _4248_ (.A(_1309_),
    .B_N(_1311_),
    .Y(_1316_));
 sky130_fd_sc_hd__buf_2 _4249_ (.A(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__or4b_4 _4250_ (.A(_2893_),
    .B(_2901_),
    .C(_2923_),
    .D_N(_2936_),
    .X(_1318_));
 sky130_fd_sc_hd__inv_2 _4251_ (.A(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__or4_1 _4252_ (.A(_0295_),
    .B(_2914_),
    .C(_0320_),
    .D(_1310_),
    .X(_1320_));
 sky130_fd_sc_hd__nor2_2 _4253_ (.A(_1319_),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__buf_2 _4254_ (.A(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__nand2_2 _4255_ (.A(_1268_),
    .B(_1302_),
    .Y(_1323_));
 sky130_fd_sc_hd__clkbuf_4 _4256_ (.A(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__a31o_1 _4257_ (.A1(_0343_),
    .A2(_2950_),
    .A3(_1319_),
    .B1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__a221o_1 _4258_ (.A1(\cu.reg_file.reg_sp[0] ),
    .A2(_0993_),
    .B1(_1322_),
    .B2(_1299_),
    .C1(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__a221o_1 _4259_ (.A1(\cu.reg_file.reg_e[0] ),
    .A2(_1315_),
    .B1(_1317_),
    .B2(\cu.reg_file.reg_l[0] ),
    .C1(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__a21oi_1 _4260_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_1313_),
    .B1(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__o21bai_4 _4261_ (.A1(_1291_),
    .A2(_1307_),
    .B1_N(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__buf_4 _4262_ (.A(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__and2_1 _4263_ (.A(\mc.rw.state[2] ),
    .B(_2699_),
    .X(_1331_));
 sky130_fd_sc_hd__clkbuf_4 _4264_ (.A(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_4 _4265_ (.A(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__nor2_1 _4266_ (.A(_2697_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__inv_2 _4267_ (.A(_1329_),
    .Y(_1335_));
 sky130_fd_sc_hd__o211a_1 _4268_ (.A1(\mc.rw.state[2] ),
    .A2(_2705_),
    .B1(_2707_),
    .C1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__a21oi_2 _4269_ (.A1(_1330_),
    .A2(_1334_),
    .B1(_1336_),
    .Y(net35));
 sky130_fd_sc_hd__a22o_1 _4270_ (.A1(\cu.reg_file.reg_a[1] ),
    .A2(_1276_),
    .B1(_1287_),
    .B2(\cu.reg_file.reg_sp[1] ),
    .X(_1337_));
 sky130_fd_sc_hd__a221o_1 _4271_ (.A1(\cu.reg_file.reg_e[1] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[1] ),
    .C1(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__a21oi_1 _4272_ (.A1(\cu.reg_file.reg_c[1] ),
    .A2(_1281_),
    .B1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__nor2_1 _4273_ (.A(_1271_),
    .B(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__a221o_1 _4274_ (.A1(_0340_),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[1] ),
    .C1(_1305_),
    .X(_1341_));
 sky130_fd_sc_hd__and2_1 _4275_ (.A(\cu.reg_file.reg_l[1] ),
    .B(_1317_),
    .X(_1342_));
 sky130_fd_sc_hd__nor2_2 _4276_ (.A(_0295_),
    .B(_1318_),
    .Y(_1343_));
 sky130_fd_sc_hd__buf_2 _4277_ (.A(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__a221o_1 _4278_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(_0340_),
    .C1(_1324_),
    .X(_1345_));
 sky130_fd_sc_hd__a221o_1 _4279_ (.A1(\cu.pc.pc_o[1] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_e[1] ),
    .C1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a211o_1 _4280_ (.A1(\cu.reg_file.reg_c[1] ),
    .A2(_1313_),
    .B1(_1342_),
    .C1(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__o21a_4 _4281_ (.A1(_1340_),
    .A2(_1341_),
    .B1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__xnor2_1 _4282_ (.A(_1332_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_1 _4283_ (.A(_1335_),
    .B(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__or2_2 _4284_ (.A(_2696_),
    .B(_1333_),
    .X(_1351_));
 sky130_fd_sc_hd__o21a_1 _4285_ (.A1(_1335_),
    .A2(_1349_),
    .B1(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__o21a_2 _4286_ (.A1(\mc.rw.state[1] ),
    .A2(\mc.rw.state[0] ),
    .B1(_2698_),
    .X(_1353_));
 sky130_fd_sc_hd__buf_4 _4287_ (.A(_1348_),
    .X(_1354_));
 sky130_fd_sc_hd__or3_1 _4288_ (.A(_2698_),
    .B(\mc.rw.state[1] ),
    .C(\mc.rw.state[0] ),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_4 _4289_ (.A(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__nor2_1 _4290_ (.A(_1356_),
    .B(_1354_),
    .Y(_1357_));
 sky130_fd_sc_hd__a221o_4 _4291_ (.A1(_1350_),
    .A2(_1352_),
    .B1(_1353_),
    .B2(_1354_),
    .C1(_1357_),
    .X(net42));
 sky130_fd_sc_hd__a22o_1 _4292_ (.A1(\cu.reg_file.reg_a[2] ),
    .A2(_1276_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[2] ),
    .X(_1358_));
 sky130_fd_sc_hd__a221o_1 _4293_ (.A1(\cu.reg_file.reg_e[2] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[2] ),
    .C1(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__a21oi_1 _4294_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_1281_),
    .B1(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__nor2_1 _4295_ (.A(_1271_),
    .B(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__a221o_1 _4296_ (.A1(_0341_),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[2] ),
    .C1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__and2_1 _4297_ (.A(\cu.reg_file.reg_e[2] ),
    .B(_1315_),
    .X(_1363_));
 sky130_fd_sc_hd__buf_4 _4298_ (.A(_1324_),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_1 _4299_ (.A1(\cu.reg_file.reg_sp[2] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(_0341_),
    .C1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__a221o_1 _4300_ (.A1(\cu.pc.pc_o[2] ),
    .A2(_1322_),
    .B1(_1317_),
    .B2(\cu.reg_file.reg_l[2] ),
    .C1(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__a211o_1 _4301_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_1313_),
    .B1(_1363_),
    .C1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__o21ai_2 _4302_ (.A1(_1306_),
    .A2(_1362_),
    .B1(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__clkbuf_4 _4303_ (.A(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__a211o_1 _4304_ (.A1(_2701_),
    .A2(_1354_),
    .B1(_1353_),
    .C1(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_4 _4305_ (.A(_2701_),
    .X(_1371_));
 sky130_fd_sc_hd__inv_2 _4306_ (.A(_1348_),
    .Y(_1372_));
 sky130_fd_sc_hd__o21a_2 _4307_ (.A1(_1306_),
    .A2(_1362_),
    .B1(_1367_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_4 _4308_ (.A(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__a21o_1 _4309_ (.A1(_1371_),
    .A2(_1372_),
    .B1(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(\mc.rw.state[2] ),
    .B(_2699_),
    .Y(_1376_));
 sky130_fd_sc_hd__a22o_1 _4311_ (.A1(_1376_),
    .A2(_1348_),
    .B1(_1349_),
    .B2(_1335_),
    .X(_1377_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_1376_),
    .B(_1374_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _4313_ (.A(_1332_),
    .B(_1368_),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_1378_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__xnor2_1 _4315_ (.A(_1377_),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__clkbuf_4 _4316_ (.A(_1351_),
    .X(_1382_));
 sky130_fd_sc_hd__a22o_1 _4317_ (.A1(_1370_),
    .A2(_1375_),
    .B1(_1381_),
    .B2(_1382_),
    .X(net43));
 sky130_fd_sc_hd__a21bo_1 _4318_ (.A1(_1377_),
    .A2(_1379_),
    .B1_N(_1378_),
    .X(_1383_));
 sky130_fd_sc_hd__a22o_1 _4319_ (.A1(\cu.reg_file.reg_a[3] ),
    .A2(_1276_),
    .B1(_1287_),
    .B2(\cu.reg_file.reg_sp[3] ),
    .X(_1384_));
 sky130_fd_sc_hd__a221o_1 _4320_ (.A1(\cu.reg_file.reg_e[3] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[3] ),
    .C1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__a21oi_1 _4321_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_1281_),
    .B1(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__nor2_1 _4322_ (.A(_1271_),
    .B(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__a221o_1 _4323_ (.A1(\cu.id.cb_opcode_y[0] ),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[3] ),
    .C1(_1305_),
    .X(_1388_));
 sky130_fd_sc_hd__and2_1 _4324_ (.A(\cu.reg_file.reg_l[3] ),
    .B(_1317_),
    .X(_1389_));
 sky130_fd_sc_hd__a221o_1 _4325_ (.A1(\cu.reg_file.reg_sp[3] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(\cu.id.cb_opcode_y[0] ),
    .C1(_1324_),
    .X(_1390_));
 sky130_fd_sc_hd__a221o_1 _4326_ (.A1(\cu.pc.pc_o[3] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_e[3] ),
    .C1(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__a211o_1 _4327_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_1313_),
    .B1(_1389_),
    .C1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__o21a_2 _4328_ (.A1(_1387_),
    .A2(_1388_),
    .B1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__or2_1 _4329_ (.A(_1376_),
    .B(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__nand2_1 _4330_ (.A(_1383_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__clkbuf_4 _4331_ (.A(_1376_),
    .X(_1396_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_1396_),
    .B(_1393_),
    .Y(_1397_));
 sky130_fd_sc_hd__or2b_1 _4333_ (.A(_1395_),
    .B_N(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__a21o_1 _4334_ (.A1(_1397_),
    .A2(_1394_),
    .B1(_1383_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_4 _4335_ (.A(_1393_),
    .X(_1400_));
 sky130_fd_sc_hd__nor2_8 _4336_ (.A(_1348_),
    .B(_1373_),
    .Y(_1401_));
 sky130_fd_sc_hd__o21ai_4 _4337_ (.A1(\mc.rw.state[1] ),
    .A2(\mc.rw.state[0] ),
    .B1(_2698_),
    .Y(_1402_));
 sky130_fd_sc_hd__o21ai_1 _4338_ (.A1(_1356_),
    .A2(_1401_),
    .B1(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__and2b_1 _4339_ (.A_N(_1393_),
    .B(_1401_),
    .X(_1404_));
 sky130_fd_sc_hd__a22o_1 _4340_ (.A1(_1400_),
    .A2(_1403_),
    .B1(_1404_),
    .B2(_1371_),
    .X(_1405_));
 sky130_fd_sc_hd__a31o_2 _4341_ (.A1(_1382_),
    .A2(_1398_),
    .A3(_1399_),
    .B1(_1405_),
    .X(net44));
 sky130_fd_sc_hd__a22o_1 _4342_ (.A1(\cu.reg_file.reg_a[4] ),
    .A2(_1276_),
    .B1(_1287_),
    .B2(\cu.reg_file.reg_sp[4] ),
    .X(_1406_));
 sky130_fd_sc_hd__a221o_1 _4343_ (.A1(\cu.reg_file.reg_e[4] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[4] ),
    .C1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__a21oi_1 _4344_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_1281_),
    .B1(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__nor2_1 _4345_ (.A(_1271_),
    .B(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__a221o_2 _4346_ (.A1(_0374_),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[4] ),
    .C1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__and2_1 _4347_ (.A(\cu.reg_file.reg_l[4] ),
    .B(_1317_),
    .X(_1411_));
 sky130_fd_sc_hd__a221o_1 _4348_ (.A1(\cu.reg_file.reg_sp[4] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(_0374_),
    .C1(_1364_),
    .X(_1412_));
 sky130_fd_sc_hd__a221o_1 _4349_ (.A1(\cu.pc.pc_o[4] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_e[4] ),
    .C1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__a211o_2 _4350_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_1313_),
    .B1(_1411_),
    .C1(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__o21a_4 _4351_ (.A1(_1306_),
    .A2(_1410_),
    .B1(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__o21ai_1 _4352_ (.A1(_1356_),
    .A2(_1404_),
    .B1(_1402_),
    .Y(_1416_));
 sky130_fd_sc_hd__o21ai_4 _4353_ (.A1(_1306_),
    .A2(_1410_),
    .B1(_1414_),
    .Y(_1417_));
 sky130_fd_sc_hd__and3_1 _4354_ (.A(_2701_),
    .B(_1404_),
    .C(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__nand2_2 _4355_ (.A(_1396_),
    .B(_1415_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_1332_),
    .B(_1417_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _4357_ (.A(_1419_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__nand3_1 _4358_ (.A(_1397_),
    .B(_1395_),
    .C(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__a21o_1 _4359_ (.A1(_1397_),
    .A2(_1395_),
    .B1(_1421_),
    .X(_1423_));
 sky130_fd_sc_hd__and3_1 _4360_ (.A(_1351_),
    .B(_1422_),
    .C(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__a211o_1 _4361_ (.A1(_1415_),
    .A2(_1416_),
    .B1(_1418_),
    .C1(_1424_),
    .X(net45));
 sky130_fd_sc_hd__a22o_1 _4362_ (.A1(\cu.reg_file.reg_a[5] ),
    .A2(_1276_),
    .B1(_1287_),
    .B2(\cu.reg_file.reg_sp[5] ),
    .X(_1425_));
 sky130_fd_sc_hd__a221o_1 _4363_ (.A1(\cu.reg_file.reg_e[5] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[5] ),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__a21oi_1 _4364_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_1281_),
    .B1(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__nor2_1 _4365_ (.A(_1271_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__a221o_1 _4366_ (.A1(_0373_),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[5] ),
    .C1(_1306_),
    .X(_1429_));
 sky130_fd_sc_hd__and2_1 _4367_ (.A(\cu.reg_file.reg_l[5] ),
    .B(_1317_),
    .X(_1430_));
 sky130_fd_sc_hd__a221o_1 _4368_ (.A1(\cu.reg_file.reg_sp[5] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(_0373_),
    .C1(_1364_),
    .X(_1431_));
 sky130_fd_sc_hd__a221o_1 _4369_ (.A1(\cu.pc.pc_o[5] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_e[5] ),
    .C1(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a211o_1 _4370_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_1313_),
    .B1(_1430_),
    .C1(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__o21a_2 _4371_ (.A1(_1428_),
    .A2(_1429_),
    .B1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__or2_1 _4372_ (.A(_1396_),
    .B(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__nand2_1 _4373_ (.A(_1396_),
    .B(_1434_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _4374_ (.A(_1435_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__a21o_1 _4375_ (.A1(_1419_),
    .A2(_1423_),
    .B1(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__nand3_1 _4376_ (.A(_1419_),
    .B(_1423_),
    .C(_1437_),
    .Y(_1439_));
 sky130_fd_sc_hd__nor2_1 _4377_ (.A(_1415_),
    .B(_1434_),
    .Y(_1440_));
 sky130_fd_sc_hd__nand2_1 _4378_ (.A(_1404_),
    .B(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__a21bo_1 _4379_ (.A1(_1404_),
    .A2(_1417_),
    .B1_N(_1434_),
    .X(_1442_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(_1441_),
    .B(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__a22o_1 _4381_ (.A1(_1353_),
    .A2(_1434_),
    .B1(_1443_),
    .B2(_1371_),
    .X(_1444_));
 sky130_fd_sc_hd__a31o_2 _4382_ (.A1(_1382_),
    .A2(_1438_),
    .A3(_1439_),
    .B1(_1444_),
    .X(net46));
 sky130_fd_sc_hd__or2_1 _4383_ (.A(_1423_),
    .B(_1437_),
    .X(_1445_));
 sky130_fd_sc_hd__a22o_1 _4384_ (.A1(\cu.reg_file.reg_a[6] ),
    .A2(_1276_),
    .B1(_1287_),
    .B2(\cu.reg_file.reg_sp[6] ),
    .X(_1446_));
 sky130_fd_sc_hd__a221o_1 _4385_ (.A1(\cu.reg_file.reg_e[6] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[6] ),
    .C1(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__a21oi_1 _4386_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_1281_),
    .B1(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__nor2_1 _4387_ (.A(_1271_),
    .B(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__a221o_1 _4388_ (.A1(_0387_),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[6] ),
    .C1(_1306_),
    .X(_1450_));
 sky130_fd_sc_hd__and2_1 _4389_ (.A(\cu.reg_file.reg_l[6] ),
    .B(_1317_),
    .X(_1451_));
 sky130_fd_sc_hd__a221o_1 _4390_ (.A1(\cu.reg_file.reg_sp[6] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(_0387_),
    .C1(_1324_),
    .X(_1452_));
 sky130_fd_sc_hd__a221o_1 _4391_ (.A1(\cu.pc.pc_o[6] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_e[6] ),
    .C1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__a211o_1 _4392_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_1313_),
    .B1(_1451_),
    .C1(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__o21a_2 _4393_ (.A1(_1449_),
    .A2(_1450_),
    .B1(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__xnor2_1 _4394_ (.A(_1396_),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__a31o_1 _4395_ (.A1(_1419_),
    .A2(_1436_),
    .A3(_1445_),
    .B1(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__nand4_1 _4396_ (.A(_1419_),
    .B(_1436_),
    .C(_1456_),
    .D(_1445_),
    .Y(_1458_));
 sky130_fd_sc_hd__a21o_1 _4397_ (.A1(_2701_),
    .A2(_1441_),
    .B1(_1353_),
    .X(_1459_));
 sky130_fd_sc_hd__nor2_1 _4398_ (.A(_1441_),
    .B(_1455_),
    .Y(_1460_));
 sky130_fd_sc_hd__a22o_1 _4399_ (.A1(_1455_),
    .A2(_1459_),
    .B1(_1460_),
    .B2(_1371_),
    .X(_1461_));
 sky130_fd_sc_hd__a31o_2 _4400_ (.A1(_1382_),
    .A2(_1457_),
    .A3(_1458_),
    .B1(_1461_),
    .X(net47));
 sky130_fd_sc_hd__inv_2 _4401_ (.A(_1455_),
    .Y(_1462_));
 sky130_fd_sc_hd__o21a_1 _4402_ (.A1(_1333_),
    .A2(_1462_),
    .B1(_1457_),
    .X(_1463_));
 sky130_fd_sc_hd__a22o_1 _4403_ (.A1(\cu.reg_file.reg_a[7] ),
    .A2(_1276_),
    .B1(_1287_),
    .B2(\cu.reg_file.reg_sp[7] ),
    .X(_1464_));
 sky130_fd_sc_hd__a221o_1 _4404_ (.A1(\cu.reg_file.reg_e[7] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_l[7] ),
    .C1(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__a21oi_1 _4405_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_1281_),
    .B1(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__nor2_1 _4406_ (.A(_1271_),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__a221o_1 _4407_ (.A1(\cu.id.cb_opcode_x[1] ),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[7] ),
    .C1(_1306_),
    .X(_1468_));
 sky130_fd_sc_hd__and2_1 _4408_ (.A(\cu.reg_file.reg_l[7] ),
    .B(_1317_),
    .X(_1469_));
 sky130_fd_sc_hd__a221o_1 _4409_ (.A1(\cu.reg_file.reg_sp[7] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(\cu.id.cb_opcode_x[1] ),
    .C1(_1324_),
    .X(_1470_));
 sky130_fd_sc_hd__a221o_1 _4410_ (.A1(\cu.pc.pc_o[7] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_e[7] ),
    .C1(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__a211o_1 _4411_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_1313_),
    .B1(_1469_),
    .C1(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__o21ai_4 _4412_ (.A1(_1467_),
    .A2(_1468_),
    .B1(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__xnor2_1 _4413_ (.A(_1332_),
    .B(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__or2_1 _4414_ (.A(_1463_),
    .B(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__nand2_1 _4415_ (.A(_1463_),
    .B(_1474_),
    .Y(_1476_));
 sky130_fd_sc_hd__o21a_1 _4416_ (.A1(_1356_),
    .A2(_1460_),
    .B1(_1402_),
    .X(_1477_));
 sky130_fd_sc_hd__nand2_1 _4417_ (.A(_1460_),
    .B(_1473_),
    .Y(_1478_));
 sky130_fd_sc_hd__o22ai_1 _4418_ (.A1(_1473_),
    .A2(_1477_),
    .B1(_1478_),
    .B2(_1356_),
    .Y(_1479_));
 sky130_fd_sc_hd__a31o_1 _4419_ (.A1(_1382_),
    .A2(_1475_),
    .A3(_1476_),
    .B1(_1479_),
    .X(net48));
 sky130_fd_sc_hd__a31o_1 _4420_ (.A1(_1440_),
    .A2(_1462_),
    .A3(_1473_),
    .B1(_1332_),
    .X(_1480_));
 sky130_fd_sc_hd__or4_1 _4421_ (.A(_1423_),
    .B(_1437_),
    .C(_1456_),
    .D(_1474_),
    .X(_1481_));
 sky130_fd_sc_hd__or2_1 _4422_ (.A(_1301_),
    .B(_1300_),
    .X(_1482_));
 sky130_fd_sc_hd__or2_2 _4423_ (.A(_1268_),
    .B(_2947_),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_2 _4424_ (.A(_1482_),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__or2_4 _4425_ (.A(_1269_),
    .B(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__a22o_1 _4426_ (.A1(\cu.reg_file.reg_d[0] ),
    .A2(_1282_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[8] ),
    .X(_1486_));
 sky130_fd_sc_hd__a221o_1 _4427_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(net144),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[0] ),
    .C1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__nor2_1 _4428_ (.A(_1269_),
    .B(_1484_),
    .Y(_1488_));
 sky130_fd_sc_hd__buf_4 _4429_ (.A(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__a221o_1 _4430_ (.A1(\cu.id.imm_i[8] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[8] ),
    .C1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__a21o_1 _4431_ (.A1(_1296_),
    .A2(_1487_),
    .B1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__o21a_1 _4432_ (.A1(\cu.pc.pc_o[8] ),
    .A2(_1485_),
    .B1(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__a221o_1 _4433_ (.A1(\cu.reg_file.reg_sp[8] ),
    .A2(_0992_),
    .B1(_1343_),
    .B2(\cu.id.imm_i[8] ),
    .C1(_1323_),
    .X(_1493_));
 sky130_fd_sc_hd__a221o_1 _4434_ (.A1(\cu.pc.pc_o[8] ),
    .A2(_1321_),
    .B1(_1314_),
    .B2(\cu.reg_file.reg_d[0] ),
    .C1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__a221o_1 _4435_ (.A1(\cu.reg_file.reg_h[0] ),
    .A2(_1316_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_b[0] ),
    .C1(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__o21a_2 _4436_ (.A1(_1305_),
    .A2(_1492_),
    .B1(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__xnor2_1 _4437_ (.A(_1396_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__a21o_1 _4438_ (.A1(_1480_),
    .A2(_1481_),
    .B1(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__nand3_1 _4439_ (.A(_1497_),
    .B(_1480_),
    .C(_1481_),
    .Y(_1499_));
 sky130_fd_sc_hd__a21o_1 _4440_ (.A1(_2701_),
    .A2(_1478_),
    .B1(_1353_),
    .X(_1500_));
 sky130_fd_sc_hd__nor2_1 _4441_ (.A(_1478_),
    .B(_1496_),
    .Y(_1501_));
 sky130_fd_sc_hd__a22o_1 _4442_ (.A1(_1496_),
    .A2(_1500_),
    .B1(_1501_),
    .B2(_1371_),
    .X(_1502_));
 sky130_fd_sc_hd__a31o_2 _4443_ (.A1(_1382_),
    .A2(_1498_),
    .A3(_1499_),
    .B1(_1502_),
    .X(net49));
 sky130_fd_sc_hd__a22o_1 _4444_ (.A1(\cu.reg_file.reg_sp[9] ),
    .A2(_1287_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_h[1] ),
    .X(_1503_));
 sky130_fd_sc_hd__a22o_1 _4445_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_1281_),
    .B1(_1283_),
    .B2(\cu.reg_file.reg_d[1] ),
    .X(_1504_));
 sky130_fd_sc_hd__o21a_1 _4446_ (.A1(_1503_),
    .A2(_1504_),
    .B1(_1296_),
    .X(_1505_));
 sky130_fd_sc_hd__a221o_1 _4447_ (.A1(\cu.id.imm_i[9] ),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[9] ),
    .C1(_1305_),
    .X(_1506_));
 sky130_fd_sc_hd__and2_1 _4448_ (.A(\cu.reg_file.reg_h[1] ),
    .B(_1316_),
    .X(_1507_));
 sky130_fd_sc_hd__a221o_1 _4449_ (.A1(\cu.reg_file.reg_sp[9] ),
    .A2(_0993_),
    .B1(_1344_),
    .B2(\cu.id.imm_i[9] ),
    .C1(_1324_),
    .X(_1508_));
 sky130_fd_sc_hd__a221o_1 _4450_ (.A1(\cu.pc.pc_o[9] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_d[1] ),
    .C1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__a211o_1 _4451_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_1313_),
    .B1(_1507_),
    .C1(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__o21ai_4 _4452_ (.A1(_1505_),
    .A2(_1506_),
    .B1(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__or2_1 _4453_ (.A(_1332_),
    .B(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__nand2_1 _4454_ (.A(_1332_),
    .B(_1511_),
    .Y(_1513_));
 sky130_fd_sc_hd__a21bo_1 _4455_ (.A1(_1396_),
    .A2(_1496_),
    .B1_N(_1498_),
    .X(_1514_));
 sky130_fd_sc_hd__a21oi_1 _4456_ (.A1(_1512_),
    .A2(_1513_),
    .B1(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__a31o_1 _4457_ (.A1(_1512_),
    .A2(_1513_),
    .A3(_1514_),
    .B1(_1334_),
    .X(_1516_));
 sky130_fd_sc_hd__and2_1 _4458_ (.A(_1501_),
    .B(_1511_),
    .X(_1517_));
 sky130_fd_sc_hd__o21a_1 _4459_ (.A1(_1356_),
    .A2(_1501_),
    .B1(_1402_),
    .X(_1518_));
 sky130_fd_sc_hd__o2bb2a_1 _4460_ (.A1_N(_1371_),
    .A2_N(_1517_),
    .B1(_1518_),
    .B2(_1511_),
    .X(_1519_));
 sky130_fd_sc_hd__o21ai_4 _4461_ (.A1(_1515_),
    .A2(_1516_),
    .B1(_1519_),
    .Y(net50));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(_1513_),
    .B(_1514_),
    .Y(_1520_));
 sky130_fd_sc_hd__clkbuf_4 _4463_ (.A(\cu.pc.pc_o[10] ),
    .X(_1521_));
 sky130_fd_sc_hd__a22o_1 _4464_ (.A1(\cu.reg_file.reg_d[2] ),
    .A2(_1282_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[10] ),
    .X(_1522_));
 sky130_fd_sc_hd__a221o_1 _4465_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(net238),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[2] ),
    .C1(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__a221o_1 _4466_ (.A1(\cu.id.imm_i[10] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(_1521_),
    .C1(_1489_),
    .X(_1524_));
 sky130_fd_sc_hd__a21o_1 _4467_ (.A1(_1296_),
    .A2(_1523_),
    .B1(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__o21a_1 _4468_ (.A1(_1521_),
    .A2(_1485_),
    .B1(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__a221o_1 _4469_ (.A1(\cu.reg_file.reg_sp[10] ),
    .A2(_0992_),
    .B1(_1344_),
    .B2(\cu.id.imm_i[10] ),
    .C1(_1324_),
    .X(_1527_));
 sky130_fd_sc_hd__a221o_1 _4470_ (.A1(_1521_),
    .A2(_1321_),
    .B1(_1314_),
    .B2(\cu.reg_file.reg_d[2] ),
    .C1(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__a221o_1 _4471_ (.A1(\cu.reg_file.reg_h[2] ),
    .A2(_1317_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_b[2] ),
    .C1(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__o21ai_4 _4472_ (.A1(_1305_),
    .A2(_1526_),
    .B1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__xnor2_1 _4473_ (.A(_1332_),
    .B(_1530_),
    .Y(_1531_));
 sky130_fd_sc_hd__a21o_1 _4474_ (.A1(_1512_),
    .A2(_1520_),
    .B1(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__nand3_1 _4475_ (.A(_1512_),
    .B(_1531_),
    .C(_1520_),
    .Y(_1533_));
 sky130_fd_sc_hd__o21a_1 _4476_ (.A1(_1356_),
    .A2(_1517_),
    .B1(_1402_),
    .X(_1534_));
 sky130_fd_sc_hd__nand2_1 _4477_ (.A(_1517_),
    .B(_1530_),
    .Y(_1535_));
 sky130_fd_sc_hd__o22ai_1 _4478_ (.A1(_1530_),
    .A2(_1534_),
    .B1(_1535_),
    .B2(_1356_),
    .Y(_1536_));
 sky130_fd_sc_hd__a31o_1 _4479_ (.A1(_1382_),
    .A2(_1532_),
    .A3(_1533_),
    .B1(_1536_),
    .X(net36));
 sky130_fd_sc_hd__a22o_1 _4480_ (.A1(\cu.reg_file.reg_d[3] ),
    .A2(_1282_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[11] ),
    .X(_1537_));
 sky130_fd_sc_hd__a221o_1 _4481_ (.A1(\cu.reg_file.reg_b[3] ),
    .A2(net144),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[3] ),
    .C1(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__a221o_1 _4482_ (.A1(\cu.id.imm_i[11] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[11] ),
    .C1(_1489_),
    .X(_1539_));
 sky130_fd_sc_hd__a21o_1 _4483_ (.A1(_1296_),
    .A2(_1538_),
    .B1(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__o21a_1 _4484_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_1485_),
    .B1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__a221o_1 _4485_ (.A1(\cu.reg_file.reg_sp[11] ),
    .A2(_0992_),
    .B1(_1343_),
    .B2(\cu.id.imm_i[11] ),
    .C1(_1324_),
    .X(_1542_));
 sky130_fd_sc_hd__a221o_1 _4486_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_1321_),
    .B1(_1314_),
    .B2(\cu.reg_file.reg_d[3] ),
    .C1(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__a221o_1 _4487_ (.A1(\cu.reg_file.reg_h[3] ),
    .A2(_1316_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_b[3] ),
    .C1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__o21ai_4 _4488_ (.A1(_1305_),
    .A2(_1541_),
    .B1(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__or2_1 _4489_ (.A(_1333_),
    .B(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__nand2_1 _4490_ (.A(_1333_),
    .B(_1545_),
    .Y(_1547_));
 sky130_fd_sc_hd__and2_1 _4491_ (.A(_1546_),
    .B(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__o21a_1 _4492_ (.A1(_1332_),
    .A2(_1530_),
    .B1(_1532_),
    .X(_1549_));
 sky130_fd_sc_hd__xnor2_1 _4493_ (.A(_1548_),
    .B(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__xor2_1 _4494_ (.A(_1535_),
    .B(_1545_),
    .X(_1551_));
 sky130_fd_sc_hd__nor2_1 _4495_ (.A(_1402_),
    .B(_1545_),
    .Y(_1552_));
 sky130_fd_sc_hd__a221o_1 _4496_ (.A1(_1351_),
    .A2(_1550_),
    .B1(_1551_),
    .B2(_1371_),
    .C1(_1552_),
    .X(net37));
 sky130_fd_sc_hd__a22o_1 _4497_ (.A1(\cu.reg_file.reg_d[4] ),
    .A2(_1282_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[12] ),
    .X(_1553_));
 sky130_fd_sc_hd__a221o_1 _4498_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(net144),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[4] ),
    .C1(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__a221o_1 _4499_ (.A1(\cu.id.imm_i[12] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[12] ),
    .C1(_1488_),
    .X(_1555_));
 sky130_fd_sc_hd__a21o_1 _4500_ (.A1(_1296_),
    .A2(_1554_),
    .B1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__o21a_1 _4501_ (.A1(\cu.pc.pc_o[12] ),
    .A2(_1485_),
    .B1(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__a221o_1 _4502_ (.A1(\cu.reg_file.reg_sp[12] ),
    .A2(_0992_),
    .B1(_1343_),
    .B2(\cu.id.imm_i[12] ),
    .C1(_1323_),
    .X(_1558_));
 sky130_fd_sc_hd__a221o_1 _4503_ (.A1(\cu.pc.pc_o[12] ),
    .A2(_1321_),
    .B1(_1314_),
    .B2(\cu.reg_file.reg_d[4] ),
    .C1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__a221o_1 _4504_ (.A1(\cu.reg_file.reg_h[4] ),
    .A2(_1316_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_b[4] ),
    .C1(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__o21ai_4 _4505_ (.A1(_1305_),
    .A2(_1557_),
    .B1(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__xnor2_1 _4506_ (.A(_1333_),
    .B(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__a21o_1 _4507_ (.A1(_1333_),
    .A2(_1545_),
    .B1(_1549_),
    .X(_1563_));
 sky130_fd_sc_hd__nand3_1 _4508_ (.A(_1546_),
    .B(_1562_),
    .C(_1563_),
    .Y(_1564_));
 sky130_fd_sc_hd__a21o_1 _4509_ (.A1(_1546_),
    .A2(_1563_),
    .B1(_1562_),
    .X(_1565_));
 sky130_fd_sc_hd__and3_1 _4510_ (.A(_1517_),
    .B(_1530_),
    .C(_1545_),
    .X(_1566_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_1566_),
    .B(_1561_),
    .Y(_1567_));
 sky130_fd_sc_hd__or2_1 _4512_ (.A(_1566_),
    .B(_1561_),
    .X(_1568_));
 sky130_fd_sc_hd__nand2_1 _4513_ (.A(_1567_),
    .B(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__a2bb2o_1 _4514_ (.A1_N(_1402_),
    .A2_N(_1561_),
    .B1(_1569_),
    .B2(_1371_),
    .X(_1570_));
 sky130_fd_sc_hd__a31o_1 _4515_ (.A1(_1382_),
    .A2(_1564_),
    .A3(_1565_),
    .B1(_1570_),
    .X(net38));
 sky130_fd_sc_hd__a22o_1 _4516_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_1282_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[13] ),
    .X(_1571_));
 sky130_fd_sc_hd__a221o_1 _4517_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(net144),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[5] ),
    .C1(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__a221o_1 _4518_ (.A1(\cu.id.imm_i[13] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[13] ),
    .C1(_1488_),
    .X(_1573_));
 sky130_fd_sc_hd__a21o_1 _4519_ (.A1(_1296_),
    .A2(_1572_),
    .B1(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__o21a_1 _4520_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_1485_),
    .B1(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__a221o_1 _4521_ (.A1(\cu.reg_file.reg_sp[13] ),
    .A2(_0992_),
    .B1(_1343_),
    .B2(\cu.id.imm_i[13] ),
    .C1(_1323_),
    .X(_1576_));
 sky130_fd_sc_hd__a221o_1 _4522_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_1321_),
    .B1(_1314_),
    .B2(\cu.reg_file.reg_d[5] ),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__a221o_1 _4523_ (.A1(\cu.reg_file.reg_h[5] ),
    .A2(_1316_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_b[5] ),
    .C1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__o21a_2 _4524_ (.A1(_1304_),
    .A2(_1575_),
    .B1(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__or2_1 _4525_ (.A(_1396_),
    .B(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(_1396_),
    .B(_1579_),
    .Y(_1581_));
 sky130_fd_sc_hd__o21ai_1 _4527_ (.A1(_1333_),
    .A2(_1561_),
    .B1(_1565_),
    .Y(_1582_));
 sky130_fd_sc_hd__a21o_1 _4528_ (.A1(_1580_),
    .A2(_1581_),
    .B1(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__a31oi_1 _4529_ (.A1(_1580_),
    .A2(_1581_),
    .A3(_1582_),
    .B1(_1334_),
    .Y(_1584_));
 sky130_fd_sc_hd__or2_1 _4530_ (.A(_1567_),
    .B(_1579_),
    .X(_1585_));
 sky130_fd_sc_hd__nand2_1 _4531_ (.A(_1567_),
    .B(_1579_),
    .Y(_1586_));
 sky130_fd_sc_hd__a21oi_1 _4532_ (.A1(_1585_),
    .A2(_1586_),
    .B1(_1356_),
    .Y(_1587_));
 sky130_fd_sc_hd__a221o_1 _4533_ (.A1(_1353_),
    .A2(_1579_),
    .B1(_1583_),
    .B2(_1584_),
    .C1(_1587_),
    .X(net39));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_1580_),
    .B(_1582_),
    .Y(_1588_));
 sky130_fd_sc_hd__nand2_1 _4535_ (.A(\cu.reg_file.reg_sp[14] ),
    .B(_1286_),
    .Y(_1589_));
 sky130_fd_sc_hd__a21bo_1 _4536_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_1283_),
    .B1_N(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__a221o_1 _4537_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(_1281_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_h[6] ),
    .C1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__a221o_1 _4538_ (.A1(\cu.id.imm_i[14] ),
    .A2(_1295_),
    .B1(_1298_),
    .B2(\cu.pc.pc_o[14] ),
    .C1(_1489_),
    .X(_1592_));
 sky130_fd_sc_hd__a21o_1 _4539_ (.A1(_1296_),
    .A2(_1591_),
    .B1(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__o21a_1 _4540_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_1485_),
    .B1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__a221o_1 _4541_ (.A1(\cu.reg_file.reg_sp[14] ),
    .A2(_0992_),
    .B1(_1344_),
    .B2(\cu.id.imm_i[14] ),
    .C1(_1324_),
    .X(_1595_));
 sky130_fd_sc_hd__a221o_1 _4542_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_1322_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_d[6] ),
    .C1(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__a221o_1 _4543_ (.A1(\cu.reg_file.reg_h[6] ),
    .A2(_1317_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_b[6] ),
    .C1(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__o21ai_4 _4544_ (.A1(_1305_),
    .A2(_1594_),
    .B1(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__or2_1 _4545_ (.A(_1333_),
    .B(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(_1333_),
    .B(_1598_),
    .Y(_1600_));
 sky130_fd_sc_hd__nand2_1 _4547_ (.A(_1599_),
    .B(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__a21o_1 _4548_ (.A1(_1581_),
    .A2(_1588_),
    .B1(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__nand3_1 _4549_ (.A(_1581_),
    .B(_1601_),
    .C(_1588_),
    .Y(_1603_));
 sky130_fd_sc_hd__xor2_1 _4550_ (.A(_1585_),
    .B(_1598_),
    .X(_1604_));
 sky130_fd_sc_hd__a2bb2o_1 _4551_ (.A1_N(_1402_),
    .A2_N(_1598_),
    .B1(_1604_),
    .B2(_1371_),
    .X(_1605_));
 sky130_fd_sc_hd__a31o_2 _4552_ (.A1(_1382_),
    .A2(_1602_),
    .A3(_1603_),
    .B1(_1605_),
    .X(net40));
 sky130_fd_sc_hd__a22o_1 _4553_ (.A1(\cu.reg_file.reg_d[7] ),
    .A2(_1282_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[15] ),
    .X(_1606_));
 sky130_fd_sc_hd__a221o_1 _4554_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(net144),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[7] ),
    .C1(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__a221o_1 _4555_ (.A1(\cu.id.imm_i[15] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[15] ),
    .C1(_1489_),
    .X(_1608_));
 sky130_fd_sc_hd__a21o_1 _4556_ (.A1(_1296_),
    .A2(_1607_),
    .B1(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__o21a_1 _4557_ (.A1(\cu.pc.pc_o[15] ),
    .A2(_1485_),
    .B1(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__a221o_1 _4558_ (.A1(\cu.reg_file.reg_sp[15] ),
    .A2(_0992_),
    .B1(_1343_),
    .B2(\cu.id.imm_i[15] ),
    .C1(_1323_),
    .X(_1611_));
 sky130_fd_sc_hd__a221o_1 _4559_ (.A1(\cu.pc.pc_o[15] ),
    .A2(_1321_),
    .B1(_1314_),
    .B2(\cu.reg_file.reg_d[7] ),
    .C1(_1611_),
    .X(_1612_));
 sky130_fd_sc_hd__a221o_1 _4560_ (.A1(\cu.reg_file.reg_h[7] ),
    .A2(_1316_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_b[7] ),
    .C1(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__o21a_1 _4561_ (.A1(_1305_),
    .A2(_1610_),
    .B1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__xnor2_1 _4562_ (.A(_1396_),
    .B(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__a21o_1 _4563_ (.A1(_1599_),
    .A2(_1602_),
    .B1(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__nand3_1 _4564_ (.A(_1599_),
    .B(_1602_),
    .C(_1615_),
    .Y(_1617_));
 sky130_fd_sc_hd__or3b_1 _4565_ (.A(_1567_),
    .B(_1579_),
    .C_N(_1598_),
    .X(_1618_));
 sky130_fd_sc_hd__or2_1 _4566_ (.A(_1356_),
    .B(_1614_),
    .X(_1619_));
 sky130_fd_sc_hd__a21o_1 _4567_ (.A1(_2701_),
    .A2(_1618_),
    .B1(_1353_),
    .X(_1620_));
 sky130_fd_sc_hd__a2bb2o_1 _4568_ (.A1_N(_1618_),
    .A2_N(_1619_),
    .B1(_1620_),
    .B2(_1614_),
    .X(_1621_));
 sky130_fd_sc_hd__a31o_1 _4569_ (.A1(_1382_),
    .A2(_1616_),
    .A3(_1617_),
    .B1(_1621_),
    .X(net41));
 sky130_fd_sc_hd__and2_4 _4570_ (.A(_0824_),
    .B(_0819_),
    .X(_1622_));
 sky130_fd_sc_hd__a22o_1 _4571_ (.A1(_2702_),
    .A2(_0619_),
    .B1(_1622_),
    .B2(_2697_),
    .X(net51));
 sky130_fd_sc_hd__nor2_8 _4572_ (.A(_0516_),
    .B(_1230_),
    .Y(_1623_));
 sky130_fd_sc_hd__a22o_1 _4573_ (.A1(_2702_),
    .A2(_1052_),
    .B1(_1623_),
    .B2(_2697_),
    .X(net52));
 sky130_fd_sc_hd__a22o_1 _4574_ (.A1(_2702_),
    .A2(_1075_),
    .B1(_1226_),
    .B2(_2697_),
    .X(net53));
 sky130_fd_sc_hd__a22o_1 _4575_ (.A1(_2702_),
    .A2(_1188_),
    .B1(_1222_),
    .B2(_2697_),
    .X(net54));
 sky130_fd_sc_hd__a22o_1 _4576_ (.A1(_2702_),
    .A2(_1190_),
    .B1(_1213_),
    .B2(_2697_),
    .X(net55));
 sky130_fd_sc_hd__a22o_1 _4577_ (.A1(_2702_),
    .A2(_1192_),
    .B1(_1209_),
    .B2(_2697_),
    .X(net56));
 sky130_fd_sc_hd__nor2_4 _4578_ (.A(_0516_),
    .B(_1200_),
    .Y(_1624_));
 sky130_fd_sc_hd__a22o_1 _4579_ (.A1(_2702_),
    .A2(_1194_),
    .B1(_1624_),
    .B2(_2697_),
    .X(net57));
 sky130_fd_sc_hd__a22o_1 _4580_ (.A1(_2702_),
    .A2(_1261_),
    .B1(_1263_),
    .B2(_2697_),
    .X(net58));
 sky130_fd_sc_hd__nand2_2 _4581_ (.A(_1329_),
    .B(_1372_),
    .Y(_1625_));
 sky130_fd_sc_hd__inv_2 _4582_ (.A(_1579_),
    .Y(_1626_));
 sky130_fd_sc_hd__or4b_1 _4583_ (.A(_1561_),
    .B(_1626_),
    .C(_1598_),
    .D_N(_1614_),
    .X(_1627_));
 sky130_fd_sc_hd__or4b_1 _4584_ (.A(_1511_),
    .B(_1530_),
    .C(_1545_),
    .D_N(_1496_),
    .X(_1628_));
 sky130_fd_sc_hd__or3_4 _4585_ (.A(_1393_),
    .B(_1627_),
    .C(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__or4_2 _4586_ (.A(_1434_),
    .B(_1462_),
    .C(_1473_),
    .D(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__a211o_1 _4587_ (.A1(_1374_),
    .A2(_1625_),
    .B1(_1630_),
    .C1(_1417_),
    .X(_1631_));
 sky130_fd_sc_hd__or2b_2 _4588_ (.A(\mc.cl.cmp_o ),
    .B_N(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__nand2_4 _4589_ (.A(_1329_),
    .B(_1401_),
    .Y(_1633_));
 sky130_fd_sc_hd__or3_2 _4590_ (.A(_1415_),
    .B(_1630_),
    .C(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__nor2_1 _4591_ (.A(_1455_),
    .B(_1473_),
    .Y(_1635_));
 sky130_fd_sc_hd__or3b_2 _4592_ (.A(_1434_),
    .B(_1629_),
    .C_N(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_1434_),
    .B(_1635_),
    .Y(_1637_));
 sky130_fd_sc_hd__nor2_1 _4594_ (.A(_1329_),
    .B(_1372_),
    .Y(_1638_));
 sky130_fd_sc_hd__or4_1 _4595_ (.A(_1373_),
    .B(_1417_),
    .C(_1637_),
    .D(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__nor2_1 _4596_ (.A(_1629_),
    .B(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__clkinv_4 _4597_ (.A(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__or3_2 _4598_ (.A(_1415_),
    .B(_1629_),
    .C(_1637_),
    .X(_1642_));
 sky130_fd_sc_hd__nand4_4 _4599_ (.A(_1634_),
    .B(_1636_),
    .C(_1641_),
    .D(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__nor2_4 _4600_ (.A(_1632_),
    .B(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__a21o_1 _4601_ (.A1(_1364_),
    .A2(_1489_),
    .B1(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__buf_4 _4602_ (.A(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__buf_2 _4603_ (.A(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_4 _4604_ (.A(_1485_),
    .X(_1648_));
 sky130_fd_sc_hd__buf_2 _4605_ (.A(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_4 _4606_ (.A(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__nor3_1 _4607_ (.A(\mc.rw.state[2] ),
    .B(\mc.rw.state[1] ),
    .C(\mc.rw.state[0] ),
    .Y(_1651_));
 sky130_fd_sc_hd__or3_1 _4608_ (.A(\mc.cc.count[2] ),
    .B(\mc.cc.count[1] ),
    .C(\mc.cc.count[0] ),
    .X(_1652_));
 sky130_fd_sc_hd__or3b_2 _4609_ (.A(_1652_),
    .B(\mc.cc.count[3] ),
    .C_N(\mc.cc.enable_edge_detector.prev_data ),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_1 _4610_ (.A0(_2701_),
    .A1(_2706_),
    .S(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__a31o_1 _4611_ (.A1(_1650_),
    .A2(_1644_),
    .A3(_1651_),
    .B1(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__a21o_1 _4612_ (.A1(_2704_),
    .A2(_1647_),
    .B1(_1655_),
    .X(\mc.rw.next_state[0] ));
 sky130_fd_sc_hd__or3b_1 _4613_ (.A(\mc.cl.cmp_o ),
    .B(_1364_),
    .C_N(_1613_),
    .X(_1656_));
 sky130_fd_sc_hd__inv_2 _4614_ (.A(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__or3_2 _4615_ (.A(_0350_),
    .B(_2940_),
    .C(_0379_),
    .X(_1658_));
 sky130_fd_sc_hd__or2_1 _4616_ (.A(_2923_),
    .B(_2903_),
    .X(_1659_));
 sky130_fd_sc_hd__nor3b_4 _4617_ (.A(_0315_),
    .B(_1658_),
    .C_N(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__clkbuf_4 _4618_ (.A(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__mux2_1 _4619_ (.A0(_1650_),
    .A1(_1657_),
    .S(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__a21o_1 _4620_ (.A1(_1651_),
    .A2(_1662_),
    .B1(_2699_),
    .X(_1663_));
 sky130_fd_sc_hd__a21o_1 _4621_ (.A1(_1647_),
    .A2(_1663_),
    .B1(_2706_),
    .X(\mc.rw.next_state[1] ));
 sky130_fd_sc_hd__inv_2 _4622_ (.A(_1653_),
    .Y(_1664_));
 sky130_fd_sc_hd__or3b_4 _4623_ (.A(_0315_),
    .B(_1658_),
    .C_N(_1659_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_4 _4624_ (.A(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_8 _4625_ (.A(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__a31o_1 _4626_ (.A1(_1651_),
    .A2(_1667_),
    .A3(_1657_),
    .B1(_1351_),
    .X(_1668_));
 sky130_fd_sc_hd__a221o_1 _4627_ (.A1(_2706_),
    .A2(_1664_),
    .B1(_1668_),
    .B2(_1647_),
    .C1(_1371_),
    .X(\mc.rw.next_state[2] ));
 sky130_fd_sc_hd__and2_1 _4628_ (.A(\ih.t.enable ),
    .B(_2869_),
    .X(_1669_));
 sky130_fd_sc_hd__clkbuf_4 _4629_ (.A(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__and2b_1 _4630_ (.A_N(\ih.t.count[0] ),
    .B(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__clkbuf_1 _4631_ (.A(_1671_),
    .X(\ih.t.next_count[0] ));
 sky130_fd_sc_hd__clkbuf_4 _4632_ (.A(_1669_),
    .X(_1672_));
 sky130_fd_sc_hd__nand2_1 _4633_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .Y(_1673_));
 sky130_fd_sc_hd__or2_1 _4634_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .X(_1674_));
 sky130_fd_sc_hd__and3_1 _4635_ (.A(_1672_),
    .B(_1673_),
    .C(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _4636_ (.A(_1675_),
    .X(\ih.t.next_count[1] ));
 sky130_fd_sc_hd__a21o_1 _4637_ (.A1(\ih.t.count[0] ),
    .A2(\ih.t.count[1] ),
    .B1(\ih.t.count[2] ),
    .X(_1676_));
 sky130_fd_sc_hd__nand3_1 _4638_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .C(\ih.t.count[2] ),
    .Y(_1677_));
 sky130_fd_sc_hd__and3_1 _4639_ (.A(_1672_),
    .B(_1676_),
    .C(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__clkbuf_1 _4640_ (.A(_1678_),
    .X(\ih.t.next_count[2] ));
 sky130_fd_sc_hd__and4_1 _4641_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .C(\ih.t.count[2] ),
    .D(\ih.t.count[3] ),
    .X(_1679_));
 sky130_fd_sc_hd__a31o_1 _4642_ (.A1(\ih.t.count[0] ),
    .A2(\ih.t.count[1] ),
    .A3(\ih.t.count[2] ),
    .B1(\ih.t.count[3] ),
    .X(_1680_));
 sky130_fd_sc_hd__and3b_1 _4643_ (.A_N(_1679_),
    .B(_1680_),
    .C(_1672_),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_1 _4644_ (.A(_1681_),
    .X(\ih.t.next_count[3] ));
 sky130_fd_sc_hd__o21ai_1 _4645_ (.A1(\ih.t.count[4] ),
    .A2(_1679_),
    .B1(_1670_),
    .Y(_1682_));
 sky130_fd_sc_hd__a21oi_1 _4646_ (.A1(net220),
    .A2(_1679_),
    .B1(_1682_),
    .Y(\ih.t.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _4647_ (.A(\ih.t.count[4] ),
    .B(\ih.t.count[5] ),
    .C(_1679_),
    .X(_1683_));
 sky130_fd_sc_hd__a21o_1 _4648_ (.A1(\ih.t.count[4] ),
    .A2(_1679_),
    .B1(\ih.t.count[5] ),
    .X(_1684_));
 sky130_fd_sc_hd__and3b_1 _4649_ (.A_N(_1683_),
    .B(_1684_),
    .C(_1672_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _4650_ (.A(_1685_),
    .X(\ih.t.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _4651_ (.A(\ih.t.count[6] ),
    .B(_1683_),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_4 _4652_ (.A(_1669_),
    .X(_1687_));
 sky130_fd_sc_hd__o21ai_1 _4653_ (.A1(net229),
    .A2(_1683_),
    .B1(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__nor2_1 _4654_ (.A(_1686_),
    .B(_1688_),
    .Y(\ih.t.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _4655_ (.A(\ih.t.count[6] ),
    .B(\ih.t.count[7] ),
    .C(_1683_),
    .X(_1689_));
 sky130_fd_sc_hd__o21ai_1 _4656_ (.A1(net227),
    .A2(_1686_),
    .B1(_1687_),
    .Y(_1690_));
 sky130_fd_sc_hd__nor2_1 _4657_ (.A(_1689_),
    .B(_1690_),
    .Y(\ih.t.next_count[7] ));
 sky130_fd_sc_hd__and2_1 _4658_ (.A(\ih.t.count[8] ),
    .B(_1689_),
    .X(_1691_));
 sky130_fd_sc_hd__o21ai_1 _4659_ (.A1(\ih.t.count[8] ),
    .A2(_1689_),
    .B1(_1687_),
    .Y(_1692_));
 sky130_fd_sc_hd__nor2_1 _4660_ (.A(_1691_),
    .B(_1692_),
    .Y(\ih.t.next_count[8] ));
 sky130_fd_sc_hd__and3_1 _4661_ (.A(\ih.t.count[8] ),
    .B(\ih.t.count[9] ),
    .C(_1689_),
    .X(_1693_));
 sky130_fd_sc_hd__o21ai_1 _4662_ (.A1(net226),
    .A2(_1691_),
    .B1(_1687_),
    .Y(_1694_));
 sky130_fd_sc_hd__nor2_1 _4663_ (.A(_1693_),
    .B(_1694_),
    .Y(\ih.t.next_count[9] ));
 sky130_fd_sc_hd__o21ai_1 _4664_ (.A1(\ih.t.count[10] ),
    .A2(_1693_),
    .B1(_1670_),
    .Y(_1695_));
 sky130_fd_sc_hd__a21oi_1 _4665_ (.A1(net215),
    .A2(_1693_),
    .B1(_1695_),
    .Y(\ih.t.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _4666_ (.A(\ih.t.count[10] ),
    .B(\ih.t.count[11] ),
    .C(_1693_),
    .X(_1696_));
 sky130_fd_sc_hd__a21o_1 _4667_ (.A1(\ih.t.count[10] ),
    .A2(_1693_),
    .B1(\ih.t.count[11] ),
    .X(_1697_));
 sky130_fd_sc_hd__and3b_1 _4668_ (.A_N(_1696_),
    .B(_1697_),
    .C(_1672_),
    .X(_1698_));
 sky130_fd_sc_hd__clkbuf_1 _4669_ (.A(_1698_),
    .X(\ih.t.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _4670_ (.A(\ih.t.count[12] ),
    .B(_1696_),
    .X(_1699_));
 sky130_fd_sc_hd__o21ai_1 _4671_ (.A1(\ih.t.count[12] ),
    .A2(_1696_),
    .B1(_1687_),
    .Y(_1700_));
 sky130_fd_sc_hd__nor2_1 _4672_ (.A(_1699_),
    .B(_1700_),
    .Y(\ih.t.next_count[12] ));
 sky130_fd_sc_hd__o21ai_1 _4673_ (.A1(\ih.t.count[13] ),
    .A2(_1699_),
    .B1(_1670_),
    .Y(_1701_));
 sky130_fd_sc_hd__a21oi_1 _4674_ (.A1(net218),
    .A2(_1699_),
    .B1(_1701_),
    .Y(\ih.t.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _4675_ (.A(\ih.t.count[13] ),
    .B(\ih.t.count[14] ),
    .C(_1699_),
    .X(_1702_));
 sky130_fd_sc_hd__a31o_1 _4676_ (.A1(\ih.t.count[12] ),
    .A2(\ih.t.count[13] ),
    .A3(_1696_),
    .B1(\ih.t.count[14] ),
    .X(_1703_));
 sky130_fd_sc_hd__and3b_1 _4677_ (.A_N(_1702_),
    .B(_1703_),
    .C(_1672_),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _4678_ (.A(_1704_),
    .X(\ih.t.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _4679_ (.A(\ih.t.count[15] ),
    .B(_1702_),
    .X(_1705_));
 sky130_fd_sc_hd__o21ai_1 _4680_ (.A1(net235),
    .A2(_1702_),
    .B1(_1687_),
    .Y(_1706_));
 sky130_fd_sc_hd__nor2_1 _4681_ (.A(_1705_),
    .B(_1706_),
    .Y(\ih.t.next_count[15] ));
 sky130_fd_sc_hd__o21ai_1 _4682_ (.A1(\ih.t.count[16] ),
    .A2(_1705_),
    .B1(_1670_),
    .Y(_1707_));
 sky130_fd_sc_hd__a21oi_1 _4683_ (.A1(net217),
    .A2(_1705_),
    .B1(_1707_),
    .Y(\ih.t.next_count[16] ));
 sky130_fd_sc_hd__and3_1 _4684_ (.A(\ih.t.count[16] ),
    .B(\ih.t.count[17] ),
    .C(_1705_),
    .X(_1708_));
 sky130_fd_sc_hd__a31o_1 _4685_ (.A1(\ih.t.count[15] ),
    .A2(\ih.t.count[16] ),
    .A3(_1702_),
    .B1(\ih.t.count[17] ),
    .X(_1709_));
 sky130_fd_sc_hd__and3b_1 _4686_ (.A_N(_1708_),
    .B(_1709_),
    .C(_1672_),
    .X(_1710_));
 sky130_fd_sc_hd__clkbuf_1 _4687_ (.A(_1710_),
    .X(\ih.t.next_count[17] ));
 sky130_fd_sc_hd__and2_1 _4688_ (.A(\ih.t.count[18] ),
    .B(_1708_),
    .X(_1711_));
 sky130_fd_sc_hd__o21ai_1 _4689_ (.A1(\ih.t.count[18] ),
    .A2(_1708_),
    .B1(_1687_),
    .Y(_1712_));
 sky130_fd_sc_hd__nor2_1 _4690_ (.A(_1711_),
    .B(_1712_),
    .Y(\ih.t.next_count[18] ));
 sky130_fd_sc_hd__o21ai_1 _4691_ (.A1(\ih.t.count[19] ),
    .A2(_1711_),
    .B1(_1670_),
    .Y(_1713_));
 sky130_fd_sc_hd__a21oi_1 _4692_ (.A1(net213),
    .A2(_1711_),
    .B1(_1713_),
    .Y(\ih.t.next_count[19] ));
 sky130_fd_sc_hd__and3_1 _4693_ (.A(\ih.t.count[19] ),
    .B(\ih.t.count[20] ),
    .C(_1711_),
    .X(_1714_));
 sky130_fd_sc_hd__a31o_1 _4694_ (.A1(\ih.t.count[18] ),
    .A2(\ih.t.count[19] ),
    .A3(_1708_),
    .B1(\ih.t.count[20] ),
    .X(_1715_));
 sky130_fd_sc_hd__and3b_1 _4695_ (.A_N(_1714_),
    .B(_1715_),
    .C(_1672_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _4696_ (.A(_1716_),
    .X(\ih.t.next_count[20] ));
 sky130_fd_sc_hd__and2_1 _4697_ (.A(\ih.t.count[21] ),
    .B(_1714_),
    .X(_1717_));
 sky130_fd_sc_hd__o21ai_1 _4698_ (.A1(net230),
    .A2(_1714_),
    .B1(_1687_),
    .Y(_1718_));
 sky130_fd_sc_hd__nor2_1 _4699_ (.A(_1717_),
    .B(_1718_),
    .Y(\ih.t.next_count[21] ));
 sky130_fd_sc_hd__o21ai_1 _4700_ (.A1(\ih.t.count[22] ),
    .A2(_1717_),
    .B1(_1670_),
    .Y(_1719_));
 sky130_fd_sc_hd__a21oi_1 _4701_ (.A1(net219),
    .A2(_1717_),
    .B1(_1719_),
    .Y(\ih.t.next_count[22] ));
 sky130_fd_sc_hd__and3_1 _4702_ (.A(\ih.t.count[22] ),
    .B(\ih.t.count[23] ),
    .C(_1717_),
    .X(_1720_));
 sky130_fd_sc_hd__a31o_1 _4703_ (.A1(\ih.t.count[21] ),
    .A2(\ih.t.count[22] ),
    .A3(_1714_),
    .B1(\ih.t.count[23] ),
    .X(_1721_));
 sky130_fd_sc_hd__and3b_1 _4704_ (.A_N(_1720_),
    .B(_1721_),
    .C(_1672_),
    .X(_1722_));
 sky130_fd_sc_hd__clkbuf_1 _4705_ (.A(_1722_),
    .X(\ih.t.next_count[23] ));
 sky130_fd_sc_hd__and2_1 _4706_ (.A(\ih.t.count[24] ),
    .B(_1720_),
    .X(_1723_));
 sky130_fd_sc_hd__o21ai_1 _4707_ (.A1(net232),
    .A2(_1720_),
    .B1(_1687_),
    .Y(_1724_));
 sky130_fd_sc_hd__nor2_1 _4708_ (.A(_1723_),
    .B(_1724_),
    .Y(\ih.t.next_count[24] ));
 sky130_fd_sc_hd__o21ai_1 _4709_ (.A1(\ih.t.count[25] ),
    .A2(_1723_),
    .B1(_1670_),
    .Y(_1725_));
 sky130_fd_sc_hd__a21oi_1 _4710_ (.A1(net222),
    .A2(_1723_),
    .B1(_1725_),
    .Y(\ih.t.next_count[25] ));
 sky130_fd_sc_hd__and3_1 _4711_ (.A(\ih.t.count[25] ),
    .B(\ih.t.count[26] ),
    .C(_1723_),
    .X(_1726_));
 sky130_fd_sc_hd__a31o_1 _4712_ (.A1(\ih.t.count[24] ),
    .A2(\ih.t.count[25] ),
    .A3(_1720_),
    .B1(\ih.t.count[26] ),
    .X(_1727_));
 sky130_fd_sc_hd__and3b_1 _4713_ (.A_N(_1726_),
    .B(_1727_),
    .C(_1669_),
    .X(_1728_));
 sky130_fd_sc_hd__clkbuf_1 _4714_ (.A(_1728_),
    .X(\ih.t.next_count[26] ));
 sky130_fd_sc_hd__and2_1 _4715_ (.A(\ih.t.count[27] ),
    .B(_1726_),
    .X(_1729_));
 sky130_fd_sc_hd__o21ai_1 _4716_ (.A1(net231),
    .A2(_1726_),
    .B1(_1687_),
    .Y(_1730_));
 sky130_fd_sc_hd__nor2_1 _4717_ (.A(_1729_),
    .B(_1730_),
    .Y(\ih.t.next_count[27] ));
 sky130_fd_sc_hd__o21ai_1 _4718_ (.A1(\ih.t.count[28] ),
    .A2(_1729_),
    .B1(_1670_),
    .Y(_1731_));
 sky130_fd_sc_hd__a21oi_1 _4719_ (.A1(net221),
    .A2(_1729_),
    .B1(_1731_),
    .Y(\ih.t.next_count[28] ));
 sky130_fd_sc_hd__and3_1 _4720_ (.A(\ih.t.count[28] ),
    .B(\ih.t.count[29] ),
    .C(_1729_),
    .X(_1732_));
 sky130_fd_sc_hd__a31o_1 _4721_ (.A1(\ih.t.count[27] ),
    .A2(\ih.t.count[28] ),
    .A3(_1726_),
    .B1(\ih.t.count[29] ),
    .X(_1733_));
 sky130_fd_sc_hd__and3b_1 _4722_ (.A_N(_1732_),
    .B(_1733_),
    .C(_1669_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _4723_ (.A(_1734_),
    .X(\ih.t.next_count[29] ));
 sky130_fd_sc_hd__o21ai_1 _4724_ (.A1(net207),
    .A2(_1732_),
    .B1(_1670_),
    .Y(_1735_));
 sky130_fd_sc_hd__a21oi_1 _4725_ (.A1(net207),
    .A2(_1732_),
    .B1(_1735_),
    .Y(\ih.t.next_count[30] ));
 sky130_fd_sc_hd__a21o_1 _4726_ (.A1(\ih.t.count[30] ),
    .A2(_1732_),
    .B1(\ih.t.count[31] ),
    .X(_1736_));
 sky130_fd_sc_hd__nand3_1 _4727_ (.A(\ih.t.count[30] ),
    .B(\ih.t.count[31] ),
    .C(_1732_),
    .Y(_1737_));
 sky130_fd_sc_hd__and3_1 _4728_ (.A(_1672_),
    .B(_1736_),
    .C(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__clkbuf_1 _4729_ (.A(_1738_),
    .X(\ih.t.next_count[31] ));
 sky130_fd_sc_hd__a21oi_4 _4730_ (.A1(_1364_),
    .A2(_1489_),
    .B1(_1644_),
    .Y(_1739_));
 sky130_fd_sc_hd__a21oi_1 _4731_ (.A1(_2946_),
    .A2(_1301_),
    .B1(_1300_),
    .Y(_1740_));
 sky130_fd_sc_hd__mux2_1 _4732_ (.A0(\cu.alu_f[6] ),
    .A1(\alu.Cin ),
    .S(_0359_),
    .X(_1741_));
 sky130_fd_sc_hd__xnor2_1 _4733_ (.A(_2893_),
    .B(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__o21ai_1 _4734_ (.A1(_2939_),
    .A2(_2916_),
    .B1(_2878_),
    .Y(_1743_));
 sky130_fd_sc_hd__or3_1 _4735_ (.A(_0303_),
    .B(_0449_),
    .C(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__a31o_1 _4736_ (.A1(_2897_),
    .A2(_2941_),
    .A3(_1742_),
    .B1(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__nor3b_1 _4737_ (.A(_0302_),
    .B(_1266_),
    .C_N(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__o21ai_2 _4738_ (.A1(_0456_),
    .A2(_1746_),
    .B1(_2950_),
    .Y(_1747_));
 sky130_fd_sc_hd__or2_1 _4739_ (.A(_1012_),
    .B(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__o32a_1 _4740_ (.A1(_2908_),
    .A2(_0361_),
    .A3(_0968_),
    .B1(_0313_),
    .B2(_0326_),
    .X(_1749_));
 sky130_fd_sc_hd__and2b_1 _4741_ (.A_N(_2922_),
    .B(_0303_),
    .X(_1750_));
 sky130_fd_sc_hd__nor2_1 _4742_ (.A(_0314_),
    .B(_1741_),
    .Y(_1751_));
 sky130_fd_sc_hd__or4_1 _4743_ (.A(_2907_),
    .B(_0311_),
    .C(_0379_),
    .D(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__o22a_1 _4744_ (.A1(_0338_),
    .A2(_1749_),
    .B1(_1750_),
    .B2(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__or4_1 _4745_ (.A(_0296_),
    .B(_0320_),
    .C(_1319_),
    .D(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__o21ai_1 _4746_ (.A1(_1483_),
    .A2(_1748_),
    .B1(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_1754_),
    .B(_1747_),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _4748_ (.A(_0371_),
    .B(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__a21oi_1 _4749_ (.A1(_1739_),
    .A2(_1757_),
    .B1(_1483_),
    .Y(_1758_));
 sky130_fd_sc_hd__o22a_1 _4750_ (.A1(_1645_),
    .A2(_1755_),
    .B1(_1758_),
    .B2(_1269_),
    .X(_1759_));
 sky130_fd_sc_hd__o22a_1 _4751_ (.A1(_1300_),
    .A2(_1739_),
    .B1(_1740_),
    .B2(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__a41o_1 _4752_ (.A1(_2880_),
    .A2(_2913_),
    .A3(_2935_),
    .A4(_0977_),
    .B1(_0350_),
    .X(_1761_));
 sky130_fd_sc_hd__and3b_1 _4753_ (.A_N(net150),
    .B(_2952_),
    .C(_0307_),
    .X(_1762_));
 sky130_fd_sc_hd__a41o_1 _4754_ (.A1(_2904_),
    .A2(_2924_),
    .A3(_1318_),
    .A4(_1762_),
    .B1(_0350_),
    .X(_1763_));
 sky130_fd_sc_hd__nand2_1 _4755_ (.A(_1756_),
    .B(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__or3b_1 _4756_ (.A(_1268_),
    .B(_1301_),
    .C_N(_1300_),
    .X(_1765_));
 sky130_fd_sc_hd__a21oi_1 _4757_ (.A1(_1761_),
    .A2(_1764_),
    .B1(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__and4bb_1 _4758_ (.A_N(_1268_),
    .B_N(_1300_),
    .C(_1756_),
    .D(_1301_),
    .X(_1767_));
 sky130_fd_sc_hd__or3_1 _4759_ (.A(_1760_),
    .B(_1766_),
    .C(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__or2_1 _4760_ (.A(net236),
    .B(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__clkbuf_1 _4761_ (.A(_1769_),
    .X(_0004_));
 sky130_fd_sc_hd__a31o_1 _4762_ (.A1(_1301_),
    .A2(_1300_),
    .A3(_1748_),
    .B1(_1268_),
    .X(_1770_));
 sky130_fd_sc_hd__nand2_1 _4763_ (.A(_1739_),
    .B(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__nor2_1 _4764_ (.A(_1268_),
    .B(_1747_),
    .Y(_1772_));
 sky130_fd_sc_hd__a21boi_1 _4765_ (.A1(_1747_),
    .A2(_1763_),
    .B1_N(_1761_),
    .Y(_1773_));
 sky130_fd_sc_hd__o22a_1 _4766_ (.A1(_1303_),
    .A2(_1772_),
    .B1(_1773_),
    .B2(_1765_),
    .X(_1774_));
 sky130_fd_sc_hd__o311a_1 _4767_ (.A1(_1483_),
    .A2(_1632_),
    .A3(_1643_),
    .B1(_1771_),
    .C1(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__nor2_1 _4768_ (.A(net206),
    .B(_1775_),
    .Y(_0005_));
 sky130_fd_sc_hd__o21a_1 _4769_ (.A1(_1300_),
    .A2(_1644_),
    .B1(_1268_),
    .X(_1776_));
 sky130_fd_sc_hd__a21oi_1 _4770_ (.A1(_1300_),
    .A2(_1761_),
    .B1(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__or4b_1 _4771_ (.A(_1268_),
    .B(_1012_),
    .C(_1646_),
    .D_N(_1301_),
    .X(_1778_));
 sky130_fd_sc_hd__o211a_1 _4772_ (.A1(_1301_),
    .A2(_1777_),
    .B1(_1778_),
    .C1(_1303_),
    .X(_1779_));
 sky130_fd_sc_hd__nor2_1 _4773_ (.A(net206),
    .B(_1779_),
    .Y(_0006_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_2948_),
    .B(_0986_),
    .Y(_1780_));
 sky130_fd_sc_hd__or4b_1 _4775_ (.A(_0976_),
    .B(_0989_),
    .C(_1780_),
    .D_N(_0994_),
    .X(_1781_));
 sky130_fd_sc_hd__or2_1 _4776_ (.A(_0980_),
    .B(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__nand2_1 _4777_ (.A(net200),
    .B(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__a21boi_1 _4778_ (.A1(net140),
    .A2(_1783_),
    .B1_N(net203),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(_1775_),
    .B(_1779_),
    .Y(_1784_));
 sky130_fd_sc_hd__o21a_1 _4780_ (.A1(_1768_),
    .A2(_1784_),
    .B1(_0350_),
    .X(_1785_));
 sky130_fd_sc_hd__o21ba_1 _4781_ (.A1(net200),
    .A2(_1785_),
    .B1_N(net204),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _4782_ (.A1(_0350_),
    .A2(_2948_),
    .B1(_1782_),
    .B2(net204),
    .X(_0002_));
 sky130_fd_sc_hd__and3_1 _4783_ (.A(_0986_),
    .B(_0989_),
    .C(_0994_),
    .X(_1786_));
 sky130_fd_sc_hd__a21oi_1 _4784_ (.A1(_1000_),
    .A2(_1786_),
    .B1(\cu.id.is_halted ),
    .Y(_1787_));
 sky130_fd_sc_hd__nor2_1 _4785_ (.A(net200),
    .B(_1787_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _4786_ (.A(_1299_),
    .Y(_1788_));
 sky130_fd_sc_hd__xor2_1 _4787_ (.A(_0343_),
    .B(_1299_),
    .X(_1789_));
 sky130_fd_sc_hd__nor2_2 _4788_ (.A(_2953_),
    .B(_0339_),
    .Y(_1790_));
 sky130_fd_sc_hd__nor2_1 _4789_ (.A(_0350_),
    .B(_0358_),
    .Y(_1791_));
 sky130_fd_sc_hd__or2_2 _4790_ (.A(_1791_),
    .B(_0366_),
    .X(_1792_));
 sky130_fd_sc_hd__or4_2 _4791_ (.A(_1186_),
    .B(_1790_),
    .C(_0352_),
    .D(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__buf_2 _4792_ (.A(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__buf_4 _4793_ (.A(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__mux2_1 _4794_ (.A0(_0617_),
    .A1(_1788_),
    .S(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__a2bb2o_2 _4795_ (.A1_N(_0986_),
    .A2_N(_1005_),
    .B1(_1786_),
    .B2(_0983_),
    .X(_1797_));
 sky130_fd_sc_hd__nand2_8 _4796_ (.A(_2948_),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__clkbuf_4 _4797_ (.A(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__mux2_1 _4798_ (.A0(_1789_),
    .A1(_1796_),
    .S(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__nor2_1 _4799_ (.A(_0310_),
    .B(_0311_),
    .Y(_1801_));
 sky130_fd_sc_hd__or2_1 _4800_ (.A(_2932_),
    .B(_0330_),
    .X(_1802_));
 sky130_fd_sc_hd__o311a_1 _4801_ (.A1(_2923_),
    .A2(_2899_),
    .A3(_2879_),
    .B1(_0314_),
    .C1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__or2b_1 _4802_ (.A(_1803_),
    .B_N(_1742_),
    .X(_1804_));
 sky130_fd_sc_hd__o22a_1 _4803_ (.A1(_2939_),
    .A2(_2916_),
    .B1(_2932_),
    .B2(_0331_),
    .X(_1805_));
 sky130_fd_sc_hd__o211a_1 _4804_ (.A1(_0306_),
    .A2(_0305_),
    .B1(_1805_),
    .C1(_2950_),
    .X(_1806_));
 sky130_fd_sc_hd__o2111a_2 _4805_ (.A1(_0359_),
    .A2(_0304_),
    .B1(_1801_),
    .C1(_1804_),
    .D1(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__o21ai_4 _4806_ (.A1(_2935_),
    .A2(_1256_),
    .B1(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__buf_4 _4807_ (.A(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__mux2_1 _4808_ (.A0(_1788_),
    .A1(_1800_),
    .S(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__o22ai_1 _4809_ (.A1(_1301_),
    .A2(_1775_),
    .B1(_1779_),
    .B2(_1268_),
    .Y(_1811_));
 sky130_fd_sc_hd__xor2_1 _4810_ (.A(_1300_),
    .B(_1768_),
    .X(_1812_));
 sky130_fd_sc_hd__a211o_1 _4811_ (.A1(_1301_),
    .A2(_1775_),
    .B1(_1811_),
    .C1(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__a22o_4 _4812_ (.A1(_2948_),
    .A2(_1808_),
    .B1(_1813_),
    .B2(_1484_),
    .X(_1814_));
 sky130_fd_sc_hd__buf_4 _4813_ (.A(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__mux2_1 _4814_ (.A0(_1299_),
    .A1(_1810_),
    .S(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_1 _4815_ (.A(_1816_),
    .X(_0016_));
 sky130_fd_sc_hd__xor2_1 _4816_ (.A(_1299_),
    .B(\cu.pc.pc_o[1] ),
    .X(_1817_));
 sky130_fd_sc_hd__xor2_1 _4817_ (.A(_0340_),
    .B(\cu.pc.pc_o[1] ),
    .X(_1818_));
 sky130_fd_sc_hd__and3_1 _4818_ (.A(_0343_),
    .B(_1299_),
    .C(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__a21oi_1 _4819_ (.A1(_0343_),
    .A2(_1299_),
    .B1(_1818_),
    .Y(_1820_));
 sky130_fd_sc_hd__nor2_1 _4820_ (.A(_1819_),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__mux2_1 _4821_ (.A0(_1050_),
    .A1(_1817_),
    .S(_1795_),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_1821_),
    .A1(_1822_),
    .S(_1799_),
    .X(_1823_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(_1817_),
    .A1(_1823_),
    .S(_1809_),
    .X(_1824_));
 sky130_fd_sc_hd__mux2_1 _4824_ (.A0(\cu.pc.pc_o[1] ),
    .A1(_1824_),
    .S(_1815_),
    .X(_1825_));
 sky130_fd_sc_hd__clkbuf_1 _4825_ (.A(_1825_),
    .X(_0017_));
 sky130_fd_sc_hd__and3_1 _4826_ (.A(_1299_),
    .B(\cu.pc.pc_o[1] ),
    .C(\cu.pc.pc_o[2] ),
    .X(_1826_));
 sky130_fd_sc_hd__a21oi_1 _4827_ (.A1(_1299_),
    .A2(\cu.pc.pc_o[1] ),
    .B1(\cu.pc.pc_o[2] ),
    .Y(_1827_));
 sky130_fd_sc_hd__nor2_1 _4828_ (.A(_1826_),
    .B(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nor2_1 _4829_ (.A(_0341_),
    .B(\cu.pc.pc_o[2] ),
    .Y(_1829_));
 sky130_fd_sc_hd__nand2_1 _4830_ (.A(_0341_),
    .B(\cu.pc.pc_o[2] ),
    .Y(_1830_));
 sky130_fd_sc_hd__and2b_1 _4831_ (.A_N(_1829_),
    .B(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__a21oi_1 _4832_ (.A1(_0340_),
    .A2(\cu.pc.pc_o[1] ),
    .B1(_1819_),
    .Y(_1832_));
 sky130_fd_sc_hd__xnor2_1 _4833_ (.A(_1831_),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(_1073_),
    .A1(_1828_),
    .S(_1795_),
    .X(_1834_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(_1833_),
    .A1(_1834_),
    .S(_1799_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _4836_ (.A0(_1828_),
    .A1(_1835_),
    .S(_1809_),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _4837_ (.A0(\cu.pc.pc_o[2] ),
    .A1(_1836_),
    .S(_1815_),
    .X(_1837_));
 sky130_fd_sc_hd__clkbuf_1 _4838_ (.A(_1837_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _4839_ (.A(\cu.pc.pc_o[3] ),
    .B(_1826_),
    .X(_1838_));
 sky130_fd_sc_hd__nor2_1 _4840_ (.A(\cu.pc.pc_o[3] ),
    .B(_1826_),
    .Y(_1839_));
 sky130_fd_sc_hd__nor2_1 _4841_ (.A(_1838_),
    .B(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__nor2_1 _4842_ (.A(\cu.id.cb_opcode_y[0] ),
    .B(\cu.pc.pc_o[3] ),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _4843_ (.A(\cu.id.cb_opcode_y[0] ),
    .B(\cu.pc.pc_o[3] ),
    .Y(_1842_));
 sky130_fd_sc_hd__and2b_1 _4844_ (.A_N(_1841_),
    .B(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__o21a_1 _4845_ (.A1(_1829_),
    .A2(_1832_),
    .B1(_1830_),
    .X(_1844_));
 sky130_fd_sc_hd__xnor2_1 _4846_ (.A(_1843_),
    .B(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__mux2_1 _4847_ (.A0(_1089_),
    .A1(_1840_),
    .S(_1795_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(_1845_),
    .A1(_1846_),
    .S(_1799_),
    .X(_1847_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(_1840_),
    .A1(_1847_),
    .S(_1809_),
    .X(_1848_));
 sky130_fd_sc_hd__mux2_1 _4850_ (.A0(\cu.pc.pc_o[3] ),
    .A1(_1848_),
    .S(_1815_),
    .X(_1849_));
 sky130_fd_sc_hd__clkbuf_1 _4851_ (.A(_1849_),
    .X(_0019_));
 sky130_fd_sc_hd__xor2_1 _4852_ (.A(\cu.pc.pc_o[4] ),
    .B(_1838_),
    .X(_1850_));
 sky130_fd_sc_hd__nor2_1 _4853_ (.A(_0374_),
    .B(\cu.pc.pc_o[4] ),
    .Y(_1851_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_0374_),
    .B(\cu.pc.pc_o[4] ),
    .Y(_1852_));
 sky130_fd_sc_hd__and2b_1 _4855_ (.A_N(_1851_),
    .B(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__o21a_1 _4856_ (.A1(_1841_),
    .A2(_1844_),
    .B1(_1842_),
    .X(_1854_));
 sky130_fd_sc_hd__xnor2_1 _4857_ (.A(_1853_),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__mux2_1 _4858_ (.A0(_1160_),
    .A1(_1850_),
    .S(_1795_),
    .X(_1856_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(_1855_),
    .A1(_1856_),
    .S(_1799_),
    .X(_1857_));
 sky130_fd_sc_hd__mux2_1 _4860_ (.A0(_1850_),
    .A1(_1857_),
    .S(_1809_),
    .X(_1858_));
 sky130_fd_sc_hd__mux2_1 _4861_ (.A0(\cu.pc.pc_o[4] ),
    .A1(_1858_),
    .S(_1815_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _4862_ (.A(_1859_),
    .X(_0020_));
 sky130_fd_sc_hd__and3_1 _4863_ (.A(\cu.pc.pc_o[5] ),
    .B(\cu.pc.pc_o[4] ),
    .C(_1838_),
    .X(_1860_));
 sky130_fd_sc_hd__a21oi_1 _4864_ (.A1(\cu.pc.pc_o[4] ),
    .A2(_1838_),
    .B1(\cu.pc.pc_o[5] ),
    .Y(_1861_));
 sky130_fd_sc_hd__nor2_1 _4865_ (.A(_1860_),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__nor2_1 _4866_ (.A(_0373_),
    .B(\cu.pc.pc_o[5] ),
    .Y(_1863_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(_0373_),
    .B(\cu.pc.pc_o[5] ),
    .Y(_1864_));
 sky130_fd_sc_hd__and2b_1 _4868_ (.A_N(_1863_),
    .B(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__o21a_1 _4869_ (.A1(_1851_),
    .A2(_1854_),
    .B1(_1852_),
    .X(_1866_));
 sky130_fd_sc_hd__xnor2_1 _4870_ (.A(_1865_),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__mux2_1 _4871_ (.A0(_1144_),
    .A1(_1862_),
    .S(_1795_),
    .X(_1868_));
 sky130_fd_sc_hd__mux2_1 _4872_ (.A0(_1867_),
    .A1(_1868_),
    .S(_1799_),
    .X(_1869_));
 sky130_fd_sc_hd__mux2_1 _4873_ (.A0(_1862_),
    .A1(_1869_),
    .S(_1809_),
    .X(_1870_));
 sky130_fd_sc_hd__mux2_1 _4874_ (.A0(\cu.pc.pc_o[5] ),
    .A1(_1870_),
    .S(_1815_),
    .X(_1871_));
 sky130_fd_sc_hd__clkbuf_1 _4875_ (.A(_1871_),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _4876_ (.A(\cu.pc.pc_o[6] ),
    .B(_1860_),
    .X(_1872_));
 sky130_fd_sc_hd__nor2_1 _4877_ (.A(\cu.pc.pc_o[6] ),
    .B(_1860_),
    .Y(_1873_));
 sky130_fd_sc_hd__nor2_1 _4878_ (.A(_1872_),
    .B(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__nor2_1 _4879_ (.A(_0387_),
    .B(\cu.pc.pc_o[6] ),
    .Y(_1875_));
 sky130_fd_sc_hd__nand2_1 _4880_ (.A(_0387_),
    .B(\cu.pc.pc_o[6] ),
    .Y(_1876_));
 sky130_fd_sc_hd__or2b_1 _4881_ (.A(_1875_),
    .B_N(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__o21a_1 _4882_ (.A1(_1863_),
    .A2(_1866_),
    .B1(_1864_),
    .X(_1878_));
 sky130_fd_sc_hd__xor2_1 _4883_ (.A(_1877_),
    .B(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__mux2_1 _4884_ (.A0(_1126_),
    .A1(_1874_),
    .S(_1795_),
    .X(_1880_));
 sky130_fd_sc_hd__mux2_1 _4885_ (.A0(_1879_),
    .A1(_1880_),
    .S(_1799_),
    .X(_1881_));
 sky130_fd_sc_hd__mux2_1 _4886_ (.A0(_1874_),
    .A1(_1881_),
    .S(_1809_),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(\cu.pc.pc_o[6] ),
    .A1(_1882_),
    .S(_1815_),
    .X(_1883_));
 sky130_fd_sc_hd__clkbuf_1 _4888_ (.A(_1883_),
    .X(_0022_));
 sky130_fd_sc_hd__xor2_1 _4889_ (.A(\cu.pc.pc_o[7] ),
    .B(_1872_),
    .X(_1884_));
 sky130_fd_sc_hd__nor2_1 _4890_ (.A(_2920_),
    .B(\cu.pc.pc_o[7] ),
    .Y(_1885_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_2920_),
    .B(\cu.pc.pc_o[7] ),
    .Y(_1886_));
 sky130_fd_sc_hd__and2b_1 _4892_ (.A_N(_1885_),
    .B(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__o21a_1 _4893_ (.A1(_1875_),
    .A2(_1878_),
    .B1(_1876_),
    .X(_1888_));
 sky130_fd_sc_hd__xnor2_1 _4894_ (.A(_1887_),
    .B(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__mux2_1 _4895_ (.A0(_1110_),
    .A1(_1884_),
    .S(_1794_),
    .X(_1890_));
 sky130_fd_sc_hd__mux2_1 _4896_ (.A0(_1889_),
    .A1(_1890_),
    .S(_1798_),
    .X(_1891_));
 sky130_fd_sc_hd__mux2_1 _4897_ (.A0(_1884_),
    .A1(_1891_),
    .S(_1809_),
    .X(_1892_));
 sky130_fd_sc_hd__mux2_1 _4898_ (.A0(\cu.pc.pc_o[7] ),
    .A1(_1892_),
    .S(_1815_),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _4899_ (.A(_1893_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _4900_ (.A(\cu.pc.pc_o[7] ),
    .B(\cu.pc.pc_o[8] ),
    .C(_1872_),
    .X(_1894_));
 sky130_fd_sc_hd__a21oi_1 _4901_ (.A1(\cu.pc.pc_o[7] ),
    .A2(_1872_),
    .B1(\cu.pc.pc_o[8] ),
    .Y(_1895_));
 sky130_fd_sc_hd__nor2_1 _4902_ (.A(_1894_),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__mux2_1 _4903_ (.A0(_1622_),
    .A1(_1896_),
    .S(_1795_),
    .X(_1897_));
 sky130_fd_sc_hd__nor2_1 _4904_ (.A(_2920_),
    .B(\cu.pc.pc_o[8] ),
    .Y(_1898_));
 sky130_fd_sc_hd__and2_1 _4905_ (.A(\cu.id.cb_opcode_x[1] ),
    .B(\cu.pc.pc_o[8] ),
    .X(_1899_));
 sky130_fd_sc_hd__or2_1 _4906_ (.A(_1898_),
    .B(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__o21a_1 _4907_ (.A1(_1885_),
    .A2(_1888_),
    .B1(_1886_),
    .X(_1901_));
 sky130_fd_sc_hd__or2_1 _4908_ (.A(_1900_),
    .B(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__a21oi_1 _4909_ (.A1(_1900_),
    .A2(_1901_),
    .B1(_1798_),
    .Y(_1903_));
 sky130_fd_sc_hd__a22o_1 _4910_ (.A1(_1799_),
    .A2(_1897_),
    .B1(_1902_),
    .B2(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _4911_ (.A0(_1896_),
    .A1(_1904_),
    .S(_1809_),
    .X(_1905_));
 sky130_fd_sc_hd__mux2_1 _4912_ (.A0(\cu.pc.pc_o[8] ),
    .A1(_1905_),
    .S(_1815_),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_1 _4913_ (.A(_1906_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _4914_ (.A(\cu.pc.pc_o[9] ),
    .B(_1894_),
    .X(_1907_));
 sky130_fd_sc_hd__nor2_1 _4915_ (.A(\cu.pc.pc_o[9] ),
    .B(_1894_),
    .Y(_1908_));
 sky130_fd_sc_hd__nor2_1 _4916_ (.A(_1907_),
    .B(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__xor2_1 _4917_ (.A(_2920_),
    .B(\cu.pc.pc_o[9] ),
    .X(_1910_));
 sky130_fd_sc_hd__or2b_1 _4918_ (.A(_1899_),
    .B_N(_1902_),
    .X(_1911_));
 sky130_fd_sc_hd__xor2_1 _4919_ (.A(_1910_),
    .B(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_1 _4920_ (.A0(_1623_),
    .A1(_1909_),
    .S(_1794_),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _4921_ (.A0(_1912_),
    .A1(_1913_),
    .S(_1798_),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _4922_ (.A0(_1909_),
    .A1(_1914_),
    .S(_1809_),
    .X(_1915_));
 sky130_fd_sc_hd__mux2_1 _4923_ (.A0(\cu.pc.pc_o[9] ),
    .A1(_1915_),
    .S(_1815_),
    .X(_1916_));
 sky130_fd_sc_hd__clkbuf_1 _4924_ (.A(_1916_),
    .X(_0025_));
 sky130_fd_sc_hd__xor2_1 _4925_ (.A(_1521_),
    .B(_1907_),
    .X(_1917_));
 sky130_fd_sc_hd__or2_1 _4926_ (.A(_2920_),
    .B(_1521_),
    .X(_1918_));
 sky130_fd_sc_hd__nand2_1 _4927_ (.A(_2920_),
    .B(_1521_),
    .Y(_1919_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_1918_),
    .B(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__o21ai_1 _4929_ (.A1(\cu.pc.pc_o[9] ),
    .A2(\cu.pc.pc_o[8] ),
    .B1(_1233_),
    .Y(_1921_));
 sky130_fd_sc_hd__or2b_1 _4930_ (.A(_1902_),
    .B_N(_1910_),
    .X(_1922_));
 sky130_fd_sc_hd__nand2_1 _4931_ (.A(_1921_),
    .B(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__xnor2_1 _4932_ (.A(_1920_),
    .B(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__mux2_1 _4933_ (.A0(_1226_),
    .A1(_1917_),
    .S(_1794_),
    .X(_1925_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(_1924_),
    .A1(_1925_),
    .S(_1798_),
    .X(_1926_));
 sky130_fd_sc_hd__mux2_1 _4935_ (.A0(_1917_),
    .A1(_1926_),
    .S(_1808_),
    .X(_1927_));
 sky130_fd_sc_hd__mux2_1 _4936_ (.A0(_1521_),
    .A1(_1927_),
    .S(_1814_),
    .X(_1928_));
 sky130_fd_sc_hd__clkbuf_1 _4937_ (.A(_1928_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _4938_ (.A(\cu.pc.pc_o[11] ),
    .B(_1521_),
    .C(_1907_),
    .X(_1929_));
 sky130_fd_sc_hd__a21oi_1 _4939_ (.A1(_1521_),
    .A2(_1907_),
    .B1(\cu.pc.pc_o[11] ),
    .Y(_1930_));
 sky130_fd_sc_hd__nor2_1 _4940_ (.A(_1929_),
    .B(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__xnor2_1 _4941_ (.A(_2920_),
    .B(\cu.pc.pc_o[11] ),
    .Y(_1932_));
 sky130_fd_sc_hd__a21bo_1 _4942_ (.A1(_1918_),
    .A2(_1923_),
    .B1_N(_1919_),
    .X(_1933_));
 sky130_fd_sc_hd__xnor2_1 _4943_ (.A(_1932_),
    .B(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__mux2_1 _4944_ (.A0(_1222_),
    .A1(_1931_),
    .S(_1794_),
    .X(_1935_));
 sky130_fd_sc_hd__mux2_1 _4945_ (.A0(_1934_),
    .A1(_1935_),
    .S(_1798_),
    .X(_1936_));
 sky130_fd_sc_hd__mux2_1 _4946_ (.A0(_1931_),
    .A1(_1936_),
    .S(_1808_),
    .X(_1937_));
 sky130_fd_sc_hd__mux2_1 _4947_ (.A0(\cu.pc.pc_o[11] ),
    .A1(_1937_),
    .S(_1814_),
    .X(_1938_));
 sky130_fd_sc_hd__clkbuf_1 _4948_ (.A(_1938_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _4949_ (.A(\cu.pc.pc_o[12] ),
    .B(_1929_),
    .X(_1939_));
 sky130_fd_sc_hd__nor2_1 _4950_ (.A(\cu.pc.pc_o[12] ),
    .B(_1929_),
    .Y(_1940_));
 sky130_fd_sc_hd__nor2_1 _4951_ (.A(_1939_),
    .B(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__mux2_1 _4952_ (.A0(_1213_),
    .A1(_1941_),
    .S(_1795_),
    .X(_1942_));
 sky130_fd_sc_hd__and2_1 _4953_ (.A(_2920_),
    .B(\cu.pc.pc_o[12] ),
    .X(_1943_));
 sky130_fd_sc_hd__nor2_1 _4954_ (.A(_1233_),
    .B(\cu.pc.pc_o[12] ),
    .Y(_1944_));
 sky130_fd_sc_hd__or2_1 _4955_ (.A(_1943_),
    .B(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__o21ai_1 _4956_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_1521_),
    .B1(_1233_),
    .Y(_1946_));
 sky130_fd_sc_hd__o311a_1 _4957_ (.A1(_1920_),
    .A2(_1922_),
    .A3(_1932_),
    .B1(_1946_),
    .C1(_1921_),
    .X(_1947_));
 sky130_fd_sc_hd__or2_1 _4958_ (.A(_1945_),
    .B(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__a21oi_1 _4959_ (.A1(_1945_),
    .A2(_1947_),
    .B1(_1798_),
    .Y(_1949_));
 sky130_fd_sc_hd__a22o_1 _4960_ (.A1(_1799_),
    .A2(_1942_),
    .B1(_1948_),
    .B2(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__mux2_1 _4961_ (.A0(_1941_),
    .A1(_1950_),
    .S(_1808_),
    .X(_1951_));
 sky130_fd_sc_hd__mux2_1 _4962_ (.A0(\cu.pc.pc_o[12] ),
    .A1(_1951_),
    .S(_1814_),
    .X(_1952_));
 sky130_fd_sc_hd__clkbuf_1 _4963_ (.A(_1952_),
    .X(_0028_));
 sky130_fd_sc_hd__xor2_1 _4964_ (.A(\cu.pc.pc_o[13] ),
    .B(_1939_),
    .X(_1953_));
 sky130_fd_sc_hd__nor2_1 _4965_ (.A(_1233_),
    .B(\cu.pc.pc_o[13] ),
    .Y(_1954_));
 sky130_fd_sc_hd__and2_1 _4966_ (.A(_1233_),
    .B(\cu.pc.pc_o[13] ),
    .X(_1955_));
 sky130_fd_sc_hd__nor2_1 _4967_ (.A(_1954_),
    .B(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__and2b_1 _4968_ (.A_N(_1943_),
    .B(_1948_),
    .X(_1957_));
 sky130_fd_sc_hd__xnor2_1 _4969_ (.A(_1956_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__mux2_1 _4970_ (.A0(_1209_),
    .A1(_1953_),
    .S(_1794_),
    .X(_1959_));
 sky130_fd_sc_hd__mux2_1 _4971_ (.A0(_1958_),
    .A1(_1959_),
    .S(_1798_),
    .X(_1960_));
 sky130_fd_sc_hd__mux2_1 _4972_ (.A0(_1953_),
    .A1(_1960_),
    .S(_1808_),
    .X(_1961_));
 sky130_fd_sc_hd__mux2_1 _4973_ (.A0(\cu.pc.pc_o[13] ),
    .A1(_1961_),
    .S(_1814_),
    .X(_1962_));
 sky130_fd_sc_hd__clkbuf_1 _4974_ (.A(_1962_),
    .X(_0029_));
 sky130_fd_sc_hd__and3_1 _4975_ (.A(\cu.pc.pc_o[14] ),
    .B(\cu.pc.pc_o[13] ),
    .C(_1939_),
    .X(_1963_));
 sky130_fd_sc_hd__a21oi_1 _4976_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_1939_),
    .B1(\cu.pc.pc_o[14] ),
    .Y(_1964_));
 sky130_fd_sc_hd__nor2_1 _4977_ (.A(_1963_),
    .B(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hd__xor2_1 _4978_ (.A(_1233_),
    .B(\cu.pc.pc_o[14] ),
    .X(_1966_));
 sky130_fd_sc_hd__and2b_1 _4979_ (.A_N(_1948_),
    .B(_1956_),
    .X(_1967_));
 sky130_fd_sc_hd__or3_1 _4980_ (.A(_1943_),
    .B(_1955_),
    .C(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__and2_1 _4981_ (.A(_1966_),
    .B(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__o21bai_1 _4982_ (.A1(_1966_),
    .A2(_1968_),
    .B1_N(_1798_),
    .Y(_1970_));
 sky130_fd_sc_hd__mux2_1 _4983_ (.A0(_1624_),
    .A1(_1965_),
    .S(_1795_),
    .X(_1971_));
 sky130_fd_sc_hd__a2bb2o_1 _4984_ (.A1_N(_1969_),
    .A2_N(_1970_),
    .B1(_1971_),
    .B2(_1799_),
    .X(_1972_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(_1965_),
    .A1(_1972_),
    .S(_1808_),
    .X(_1973_));
 sky130_fd_sc_hd__mux2_1 _4986_ (.A0(\cu.pc.pc_o[14] ),
    .A1(_1973_),
    .S(_1814_),
    .X(_1974_));
 sky130_fd_sc_hd__clkbuf_1 _4987_ (.A(_1974_),
    .X(_0030_));
 sky130_fd_sc_hd__xor2_1 _4988_ (.A(\cu.pc.pc_o[15] ),
    .B(_1963_),
    .X(_1975_));
 sky130_fd_sc_hd__o21a_1 _4989_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_1968_),
    .B1(_1233_),
    .X(_1976_));
 sky130_fd_sc_hd__o21ba_1 _4990_ (.A1(_1233_),
    .A2(_1969_),
    .B1_N(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__xor2_1 _4991_ (.A(\cu.pc.pc_o[15] ),
    .B(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _4992_ (.A0(_1263_),
    .A1(_1975_),
    .S(_1794_),
    .X(_1979_));
 sky130_fd_sc_hd__mux2_1 _4993_ (.A0(_1978_),
    .A1(_1979_),
    .S(_1798_),
    .X(_1980_));
 sky130_fd_sc_hd__mux2_1 _4994_ (.A0(_1975_),
    .A1(_1980_),
    .S(_1808_),
    .X(_1981_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(\cu.pc.pc_o[15] ),
    .A1(_1981_),
    .S(_1814_),
    .X(_1982_));
 sky130_fd_sc_hd__clkbuf_1 _4996_ (.A(_1982_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _4997_ (.A0(_0618_),
    .A1(_1622_),
    .S(_0368_),
    .X(_1983_));
 sky130_fd_sc_hd__and3_1 _4998_ (.A(_2951_),
    .B(_0367_),
    .C(_0352_),
    .X(_1984_));
 sky130_fd_sc_hd__clkbuf_4 _4999_ (.A(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__mux2_1 _5000_ (.A0(\cu.reg_file.reg_a[0] ),
    .A1(_1983_),
    .S(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__clkbuf_1 _5001_ (.A(_1986_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _5002_ (.A0(_1051_),
    .A1(_1623_),
    .S(_0368_),
    .X(_1987_));
 sky130_fd_sc_hd__mux2_1 _5003_ (.A0(\cu.reg_file.reg_a[1] ),
    .A1(_1987_),
    .S(_1985_),
    .X(_1988_));
 sky130_fd_sc_hd__clkbuf_1 _5004_ (.A(_1988_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _5005_ (.A0(_1074_),
    .A1(_1226_),
    .S(_0368_),
    .X(_1989_));
 sky130_fd_sc_hd__mux2_1 _5006_ (.A0(\cu.reg_file.reg_a[2] ),
    .A1(_1989_),
    .S(_1985_),
    .X(_1990_));
 sky130_fd_sc_hd__clkbuf_1 _5007_ (.A(_1990_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _5008_ (.A0(_1187_),
    .A1(_1222_),
    .S(_0368_),
    .X(_1991_));
 sky130_fd_sc_hd__mux2_1 _5009_ (.A0(\cu.reg_file.reg_a[3] ),
    .A1(_1991_),
    .S(_1985_),
    .X(_1992_));
 sky130_fd_sc_hd__clkbuf_1 _5010_ (.A(_1992_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(_1189_),
    .A1(_1213_),
    .S(_0368_),
    .X(_1993_));
 sky130_fd_sc_hd__mux2_1 _5012_ (.A0(\cu.reg_file.reg_a[4] ),
    .A1(_1993_),
    .S(_1985_),
    .X(_1994_));
 sky130_fd_sc_hd__clkbuf_1 _5013_ (.A(_1994_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _5014_ (.A0(_1191_),
    .A1(_1209_),
    .S(_0368_),
    .X(_1995_));
 sky130_fd_sc_hd__mux2_1 _5015_ (.A0(\cu.reg_file.reg_a[5] ),
    .A1(_1995_),
    .S(_1985_),
    .X(_1996_));
 sky130_fd_sc_hd__clkbuf_1 _5016_ (.A(_1996_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _5017_ (.A0(_1193_),
    .A1(_1624_),
    .S(_0368_),
    .X(_1997_));
 sky130_fd_sc_hd__mux2_1 _5018_ (.A0(\cu.reg_file.reg_a[6] ),
    .A1(_1997_),
    .S(_1985_),
    .X(_1998_));
 sky130_fd_sc_hd__clkbuf_1 _5019_ (.A(_1998_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _5020_ (.A0(_1260_),
    .A1(_1263_),
    .S(_0368_),
    .X(_1999_));
 sky130_fd_sc_hd__mux2_1 _5021_ (.A0(\cu.reg_file.reg_a[7] ),
    .A1(_1999_),
    .S(_1985_),
    .X(_2000_));
 sky130_fd_sc_hd__clkbuf_1 _5022_ (.A(_2000_),
    .X(_0039_));
 sky130_fd_sc_hd__and4b_1 _5023_ (.A_N(_1790_),
    .B(_0352_),
    .C(_1791_),
    .D(_0366_),
    .X(_2001_));
 sky130_fd_sc_hd__buf_4 _5024_ (.A(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _5025_ (.A0(_0618_),
    .A1(_1622_),
    .S(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_1790_),
    .B(_0352_),
    .Y(_2004_));
 sky130_fd_sc_hd__nor2_1 _5027_ (.A(_1792_),
    .B(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__o21a_4 _5028_ (.A1(_2002_),
    .A2(_2005_),
    .B1(_2951_),
    .X(_2006_));
 sky130_fd_sc_hd__mux2_1 _5029_ (.A0(\cu.reg_file.reg_b[0] ),
    .A1(_2003_),
    .S(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__clkbuf_1 _5030_ (.A(_2007_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _5031_ (.A0(_1051_),
    .A1(_1623_),
    .S(_2002_),
    .X(_2008_));
 sky130_fd_sc_hd__mux2_1 _5032_ (.A0(\cu.reg_file.reg_b[1] ),
    .A1(_2008_),
    .S(_2006_),
    .X(_2009_));
 sky130_fd_sc_hd__clkbuf_1 _5033_ (.A(_2009_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _5034_ (.A0(_1074_),
    .A1(_1226_),
    .S(_2002_),
    .X(_2010_));
 sky130_fd_sc_hd__mux2_1 _5035_ (.A0(\cu.reg_file.reg_b[2] ),
    .A1(_2010_),
    .S(_2006_),
    .X(_2011_));
 sky130_fd_sc_hd__clkbuf_1 _5036_ (.A(_2011_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _5037_ (.A0(_1187_),
    .A1(_1222_),
    .S(_2002_),
    .X(_2012_));
 sky130_fd_sc_hd__mux2_1 _5038_ (.A0(\cu.reg_file.reg_b[3] ),
    .A1(_2012_),
    .S(_2006_),
    .X(_2013_));
 sky130_fd_sc_hd__clkbuf_1 _5039_ (.A(_2013_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _5040_ (.A0(_1189_),
    .A1(_1213_),
    .S(_2002_),
    .X(_2014_));
 sky130_fd_sc_hd__mux2_1 _5041_ (.A0(\cu.reg_file.reg_b[4] ),
    .A1(_2014_),
    .S(_2006_),
    .X(_2015_));
 sky130_fd_sc_hd__clkbuf_1 _5042_ (.A(_2015_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _5043_ (.A0(_1191_),
    .A1(_1209_),
    .S(_2002_),
    .X(_2016_));
 sky130_fd_sc_hd__mux2_1 _5044_ (.A0(\cu.reg_file.reg_b[5] ),
    .A1(_2016_),
    .S(_2006_),
    .X(_2017_));
 sky130_fd_sc_hd__clkbuf_1 _5045_ (.A(_2017_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _5046_ (.A0(_1193_),
    .A1(_1624_),
    .S(_2002_),
    .X(_2018_));
 sky130_fd_sc_hd__mux2_1 _5047_ (.A0(\cu.reg_file.reg_b[6] ),
    .A1(_2018_),
    .S(_2006_),
    .X(_2019_));
 sky130_fd_sc_hd__clkbuf_1 _5048_ (.A(_2019_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(_1260_),
    .A1(_1263_),
    .S(_2002_),
    .X(_2020_));
 sky130_fd_sc_hd__mux2_1 _5050_ (.A0(\cu.reg_file.reg_b[7] ),
    .A1(_2020_),
    .S(_2006_),
    .X(_2021_));
 sky130_fd_sc_hd__clkbuf_1 _5051_ (.A(_2021_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_4 _5052_ (.A(_0618_),
    .X(_2022_));
 sky130_fd_sc_hd__or3_1 _5053_ (.A(_0350_),
    .B(_0358_),
    .C(_0366_),
    .X(_2023_));
 sky130_fd_sc_hd__nor2_1 _5054_ (.A(_2004_),
    .B(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__o21a_4 _5055_ (.A1(_2002_),
    .A2(_2024_),
    .B1(_2951_),
    .X(_2025_));
 sky130_fd_sc_hd__mux2_1 _5056_ (.A0(\cu.reg_file.reg_c[0] ),
    .A1(_2022_),
    .S(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__clkbuf_1 _5057_ (.A(_2026_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _5058_ (.A0(\cu.reg_file.reg_c[1] ),
    .A1(_1051_),
    .S(_2025_),
    .X(_2027_));
 sky130_fd_sc_hd__clkbuf_1 _5059_ (.A(_2027_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _5060_ (.A0(\cu.reg_file.reg_c[2] ),
    .A1(_1074_),
    .S(_2025_),
    .X(_2028_));
 sky130_fd_sc_hd__clkbuf_1 _5061_ (.A(_2028_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _5062_ (.A0(\cu.reg_file.reg_c[3] ),
    .A1(_1187_),
    .S(_2025_),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _5063_ (.A(_2029_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _5064_ (.A0(\cu.reg_file.reg_c[4] ),
    .A1(_1189_),
    .S(_2025_),
    .X(_2030_));
 sky130_fd_sc_hd__clkbuf_1 _5065_ (.A(_2030_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _5066_ (.A0(\cu.reg_file.reg_c[5] ),
    .A1(_1191_),
    .S(_2025_),
    .X(_2031_));
 sky130_fd_sc_hd__clkbuf_1 _5067_ (.A(_2031_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _5068_ (.A0(\cu.reg_file.reg_c[6] ),
    .A1(_1193_),
    .S(_2025_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _5069_ (.A(_2032_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(\cu.reg_file.reg_c[7] ),
    .A1(_1260_),
    .S(_2025_),
    .X(_2033_));
 sky130_fd_sc_hd__clkbuf_1 _5071_ (.A(_2033_),
    .X(_0055_));
 sky130_fd_sc_hd__or3_2 _5072_ (.A(_1790_),
    .B(_0348_),
    .C(_0351_),
    .X(_2034_));
 sky130_fd_sc_hd__nor2_8 _5073_ (.A(_2034_),
    .B(_1792_),
    .Y(_2035_));
 sky130_fd_sc_hd__mux2_1 _5074_ (.A0(_0617_),
    .A1(_1622_),
    .S(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__and2b_1 _5075_ (.A_N(_0352_),
    .B(_1790_),
    .X(_2037_));
 sky130_fd_sc_hd__and2_1 _5076_ (.A(_0367_),
    .B(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__o21a_4 _5077_ (.A1(_2035_),
    .A2(_2038_),
    .B1(_2951_),
    .X(_2039_));
 sky130_fd_sc_hd__mux2_1 _5078_ (.A0(\cu.reg_file.reg_d[0] ),
    .A1(_2036_),
    .S(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__clkbuf_1 _5079_ (.A(_2040_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _5080_ (.A0(_1051_),
    .A1(_1623_),
    .S(_2035_),
    .X(_2041_));
 sky130_fd_sc_hd__mux2_1 _5081_ (.A0(\cu.reg_file.reg_d[1] ),
    .A1(_2041_),
    .S(_2039_),
    .X(_2042_));
 sky130_fd_sc_hd__clkbuf_1 _5082_ (.A(_2042_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _5083_ (.A0(_1074_),
    .A1(_1226_),
    .S(_2035_),
    .X(_2043_));
 sky130_fd_sc_hd__mux2_1 _5084_ (.A0(\cu.reg_file.reg_d[2] ),
    .A1(_2043_),
    .S(_2039_),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _5085_ (.A(_2044_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _5086_ (.A0(_1187_),
    .A1(_1222_),
    .S(_2035_),
    .X(_2045_));
 sky130_fd_sc_hd__mux2_1 _5087_ (.A0(\cu.reg_file.reg_d[3] ),
    .A1(_2045_),
    .S(_2039_),
    .X(_2046_));
 sky130_fd_sc_hd__clkbuf_1 _5088_ (.A(_2046_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _5089_ (.A0(_1189_),
    .A1(_1213_),
    .S(_2035_),
    .X(_2047_));
 sky130_fd_sc_hd__mux2_1 _5090_ (.A0(\cu.reg_file.reg_d[4] ),
    .A1(_2047_),
    .S(_2039_),
    .X(_2048_));
 sky130_fd_sc_hd__clkbuf_1 _5091_ (.A(_2048_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _5092_ (.A0(_1191_),
    .A1(_1209_),
    .S(_2035_),
    .X(_2049_));
 sky130_fd_sc_hd__mux2_1 _5093_ (.A0(\cu.reg_file.reg_d[5] ),
    .A1(_2049_),
    .S(_2039_),
    .X(_2050_));
 sky130_fd_sc_hd__clkbuf_1 _5094_ (.A(_2050_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _5095_ (.A0(_1193_),
    .A1(_1624_),
    .S(_2035_),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_1 _5096_ (.A0(\cu.reg_file.reg_d[6] ),
    .A1(_2051_),
    .S(_2039_),
    .X(_2052_));
 sky130_fd_sc_hd__clkbuf_1 _5097_ (.A(_2052_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _5098_ (.A0(_1110_),
    .A1(_1263_),
    .S(_2035_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2_1 _5099_ (.A0(\cu.reg_file.reg_d[7] ),
    .A1(_2053_),
    .S(_2039_),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _5100_ (.A(_2054_),
    .X(_0063_));
 sky130_fd_sc_hd__and3_1 _5101_ (.A(_1791_),
    .B(_0366_),
    .C(_2037_),
    .X(_2055_));
 sky130_fd_sc_hd__o21a_4 _5102_ (.A1(_2035_),
    .A2(_2055_),
    .B1(_2951_),
    .X(_2056_));
 sky130_fd_sc_hd__mux2_1 _5103_ (.A0(\cu.reg_file.reg_e[0] ),
    .A1(_2022_),
    .S(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__clkbuf_1 _5104_ (.A(_2057_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(\cu.reg_file.reg_e[1] ),
    .A1(_1051_),
    .S(_2056_),
    .X(_2058_));
 sky130_fd_sc_hd__clkbuf_1 _5106_ (.A(_2058_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(\cu.reg_file.reg_e[2] ),
    .A1(_1074_),
    .S(_2056_),
    .X(_2059_));
 sky130_fd_sc_hd__clkbuf_1 _5108_ (.A(_2059_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _5109_ (.A0(\cu.reg_file.reg_e[3] ),
    .A1(_1187_),
    .S(_2056_),
    .X(_2060_));
 sky130_fd_sc_hd__clkbuf_1 _5110_ (.A(_2060_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(\cu.reg_file.reg_e[4] ),
    .A1(_1189_),
    .S(_2056_),
    .X(_2061_));
 sky130_fd_sc_hd__clkbuf_1 _5112_ (.A(_2061_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(\cu.reg_file.reg_e[5] ),
    .A1(_1191_),
    .S(_2056_),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _5114_ (.A(_2062_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(\cu.reg_file.reg_e[6] ),
    .A1(_1193_),
    .S(_2056_),
    .X(_2063_));
 sky130_fd_sc_hd__clkbuf_1 _5116_ (.A(_2063_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(\cu.reg_file.reg_e[7] ),
    .A1(_1260_),
    .S(_2056_),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _5118_ (.A(_2064_),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _5119_ (.A(_2034_),
    .B(_2023_),
    .X(_2065_));
 sky130_fd_sc_hd__buf_4 _5120_ (.A(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__mux2_1 _5121_ (.A0(_1622_),
    .A1(_0617_),
    .S(_2066_),
    .X(_2067_));
 sky130_fd_sc_hd__or3b_1 _5122_ (.A(_0352_),
    .B(_1792_),
    .C_N(_1790_),
    .X(_2068_));
 sky130_fd_sc_hd__a21bo_4 _5123_ (.A1(_2066_),
    .A2(_2068_),
    .B1_N(_2951_),
    .X(_2069_));
 sky130_fd_sc_hd__mux2_1 _5124_ (.A0(_2067_),
    .A1(\cu.reg_file.reg_h[0] ),
    .S(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__clkbuf_1 _5125_ (.A(_2070_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _5126_ (.A0(_1623_),
    .A1(_1050_),
    .S(_2066_),
    .X(_2071_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(_2071_),
    .A1(\cu.reg_file.reg_h[1] ),
    .S(_2069_),
    .X(_2072_));
 sky130_fd_sc_hd__clkbuf_1 _5128_ (.A(_2072_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(_1226_),
    .A1(_1073_),
    .S(_2066_),
    .X(_2073_));
 sky130_fd_sc_hd__mux2_1 _5130_ (.A0(_2073_),
    .A1(\cu.reg_file.reg_h[2] ),
    .S(_2069_),
    .X(_2074_));
 sky130_fd_sc_hd__clkbuf_1 _5131_ (.A(_2074_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _5132_ (.A0(_1222_),
    .A1(_1089_),
    .S(_2066_),
    .X(_2075_));
 sky130_fd_sc_hd__mux2_1 _5133_ (.A0(_2075_),
    .A1(\cu.reg_file.reg_h[3] ),
    .S(_2069_),
    .X(_2076_));
 sky130_fd_sc_hd__clkbuf_1 _5134_ (.A(_2076_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _5135_ (.A0(_1213_),
    .A1(_1160_),
    .S(_2066_),
    .X(_2077_));
 sky130_fd_sc_hd__mux2_1 _5136_ (.A0(_2077_),
    .A1(\cu.reg_file.reg_h[4] ),
    .S(_2069_),
    .X(_2078_));
 sky130_fd_sc_hd__clkbuf_1 _5137_ (.A(_2078_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _5138_ (.A0(_1209_),
    .A1(_1144_),
    .S(_2066_),
    .X(_2079_));
 sky130_fd_sc_hd__mux2_1 _5139_ (.A0(_2079_),
    .A1(\cu.reg_file.reg_h[5] ),
    .S(_2069_),
    .X(_2080_));
 sky130_fd_sc_hd__clkbuf_1 _5140_ (.A(_2080_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _5141_ (.A0(_1624_),
    .A1(_1126_),
    .S(_2066_),
    .X(_2081_));
 sky130_fd_sc_hd__mux2_1 _5142_ (.A0(_2081_),
    .A1(\cu.reg_file.reg_h[6] ),
    .S(_2069_),
    .X(_2082_));
 sky130_fd_sc_hd__clkbuf_1 _5143_ (.A(_2082_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _5144_ (.A0(_1263_),
    .A1(_1110_),
    .S(_2066_),
    .X(_2083_));
 sky130_fd_sc_hd__mux2_1 _5145_ (.A0(_2083_),
    .A1(\cu.reg_file.reg_h[7] ),
    .S(_2069_),
    .X(_2084_));
 sky130_fd_sc_hd__clkbuf_1 _5146_ (.A(_2084_),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_4 _5147_ (.A(_0618_),
    .X(_2085_));
 sky130_fd_sc_hd__inv_2 _5148_ (.A(_2023_),
    .Y(_2086_));
 sky130_fd_sc_hd__and3_1 _5149_ (.A(_2951_),
    .B(_2004_),
    .C(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__clkbuf_4 _5150_ (.A(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(\cu.reg_file.reg_l[0] ),
    .A1(_2085_),
    .S(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__clkbuf_1 _5152_ (.A(_2089_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(\cu.reg_file.reg_l[1] ),
    .A1(_1051_),
    .S(_2088_),
    .X(_2090_));
 sky130_fd_sc_hd__clkbuf_1 _5154_ (.A(_2090_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(\cu.reg_file.reg_l[2] ),
    .A1(_1074_),
    .S(_2088_),
    .X(_2091_));
 sky130_fd_sc_hd__clkbuf_1 _5156_ (.A(_2091_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _5157_ (.A0(\cu.reg_file.reg_l[3] ),
    .A1(_1187_),
    .S(_2088_),
    .X(_2092_));
 sky130_fd_sc_hd__clkbuf_1 _5158_ (.A(_2092_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _5159_ (.A0(\cu.reg_file.reg_l[4] ),
    .A1(_1189_),
    .S(_2088_),
    .X(_2093_));
 sky130_fd_sc_hd__clkbuf_1 _5160_ (.A(_2093_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _5161_ (.A0(\cu.reg_file.reg_l[5] ),
    .A1(_1191_),
    .S(_2088_),
    .X(_2094_));
 sky130_fd_sc_hd__clkbuf_1 _5162_ (.A(_2094_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _5163_ (.A0(\cu.reg_file.reg_l[6] ),
    .A1(_1193_),
    .S(_2088_),
    .X(_2095_));
 sky130_fd_sc_hd__clkbuf_1 _5164_ (.A(_2095_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(\cu.reg_file.reg_l[7] ),
    .A1(_1260_),
    .S(_2088_),
    .X(_2096_));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(_2096_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _5167_ (.A0(\mc.cl.next_data[8] ),
    .A1(net18),
    .S(\mc.count ),
    .X(_2097_));
 sky130_fd_sc_hd__and2_1 _5168_ (.A(_1647_),
    .B(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__clkbuf_1 _5169_ (.A(_2098_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _5170_ (.A0(\mc.cl.next_data[9] ),
    .A1(net19),
    .S(\mc.count ),
    .X(_2099_));
 sky130_fd_sc_hd__and2_1 _5171_ (.A(_1647_),
    .B(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__clkbuf_1 _5172_ (.A(_2100_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _5173_ (.A0(\mc.cl.next_data[10] ),
    .A1(net20),
    .S(\mc.count ),
    .X(_2101_));
 sky130_fd_sc_hd__and2_1 _5174_ (.A(_1647_),
    .B(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__clkbuf_1 _5175_ (.A(_2102_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _5176_ (.A0(\mc.cl.next_data[11] ),
    .A1(net21),
    .S(\mc.count ),
    .X(_2103_));
 sky130_fd_sc_hd__and2_1 _5177_ (.A(_1647_),
    .B(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__clkbuf_1 _5178_ (.A(_2104_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _5179_ (.A0(\mc.cl.next_data[12] ),
    .A1(net22),
    .S(\mc.count ),
    .X(_2105_));
 sky130_fd_sc_hd__and2_1 _5180_ (.A(_1647_),
    .B(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__clkbuf_1 _5181_ (.A(_2106_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _5182_ (.A0(\mc.cl.next_data[13] ),
    .A1(net23),
    .S(\mc.count ),
    .X(_2107_));
 sky130_fd_sc_hd__and2_1 _5183_ (.A(_1647_),
    .B(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__clkbuf_1 _5184_ (.A(_2108_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _5185_ (.A0(\mc.cl.next_data[14] ),
    .A1(net24),
    .S(\mc.count ),
    .X(_2109_));
 sky130_fd_sc_hd__and2_1 _5186_ (.A(_1647_),
    .B(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__clkbuf_1 _5187_ (.A(_2110_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_2 _5188_ (.A(_1646_),
    .X(_2111_));
 sky130_fd_sc_hd__mux2_1 _5189_ (.A0(\mc.cl.next_data[15] ),
    .A1(net25),
    .S(\mc.count ),
    .X(_2112_));
 sky130_fd_sc_hd__and2_1 _5190_ (.A(_2111_),
    .B(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__clkbuf_1 _5191_ (.A(_2113_),
    .X(_0095_));
 sky130_fd_sc_hd__or3b_1 _5192_ (.A(_1790_),
    .B(_0352_),
    .C_N(_2951_),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_2 _5193_ (.A(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__inv_2 _5194_ (.A(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__mux2_1 _5195_ (.A0(\cu.reg_file.reg_sp[0] ),
    .A1(_2085_),
    .S(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_1 _5196_ (.A(_2117_),
    .X(_0096_));
 sky130_fd_sc_hd__or2_2 _5197_ (.A(\mc.cc.count[0] ),
    .B(_2708_),
    .X(_2118_));
 sky130_fd_sc_hd__o21ba_1 _5198_ (.A1(\mc.cc.count[3] ),
    .A2(_1652_),
    .B1_N(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__a22o_1 _5199_ (.A1(net210),
    .A2(_2708_),
    .B1(_2119_),
    .B2(\mc.cc.enable_edge_detector.prev_data ),
    .X(_0097_));
 sky130_fd_sc_hd__or2_1 _5200_ (.A(\mc.cc.enable_edge_detector.prev_data ),
    .B(_2708_),
    .X(_2120_));
 sky130_fd_sc_hd__o21ai_1 _5201_ (.A1(\mc.cc.count[1] ),
    .A2(_2118_),
    .B1(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__a21o_1 _5202_ (.A1(net228),
    .A2(_2118_),
    .B1(_2121_),
    .X(_0098_));
 sky130_fd_sc_hd__nor3_1 _5203_ (.A(\mc.cc.count[2] ),
    .B(\mc.cc.count[1] ),
    .C(_2118_),
    .Y(_2122_));
 sky130_fd_sc_hd__o211a_1 _5204_ (.A1(\mc.cc.count[1] ),
    .A2(_2118_),
    .B1(_2120_),
    .C1(\mc.cc.count[2] ),
    .X(_2123_));
 sky130_fd_sc_hd__a31o_1 _5205_ (.A1(net223),
    .A2(\mc.cc.enable_edge_detector.prev_data ),
    .A3(_2122_),
    .B1(_2123_),
    .X(_0099_));
 sky130_fd_sc_hd__and3b_1 _5206_ (.A_N(_2122_),
    .B(\mc.cc.count[3] ),
    .C(_2120_),
    .X(_2124_));
 sky130_fd_sc_hd__clkbuf_1 _5207_ (.A(_2124_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_4 _5208_ (.A(_1634_),
    .X(_2125_));
 sky130_fd_sc_hd__or2_1 _5209_ (.A(_1364_),
    .B(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__clkbuf_4 _5210_ (.A(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(_0619_),
    .A1(\ih.gpio_interrupt_mask[0] ),
    .S(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _5212_ (.A(_2128_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _5213_ (.A0(_1052_),
    .A1(\ih.gpio_interrupt_mask[1] ),
    .S(_2127_),
    .X(_2129_));
 sky130_fd_sc_hd__clkbuf_1 _5214_ (.A(_2129_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _5215_ (.A0(_1075_),
    .A1(\ih.gpio_interrupt_mask[2] ),
    .S(_2127_),
    .X(_2130_));
 sky130_fd_sc_hd__clkbuf_1 _5216_ (.A(_2130_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _5217_ (.A0(_1188_),
    .A1(\ih.gpio_interrupt_mask[3] ),
    .S(_2127_),
    .X(_2131_));
 sky130_fd_sc_hd__clkbuf_1 _5218_ (.A(_2131_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(_1190_),
    .A1(\ih.gpio_interrupt_mask[4] ),
    .S(_2127_),
    .X(_2132_));
 sky130_fd_sc_hd__clkbuf_1 _5220_ (.A(_2132_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _5221_ (.A0(_1192_),
    .A1(\ih.gpio_interrupt_mask[5] ),
    .S(_2127_),
    .X(_2133_));
 sky130_fd_sc_hd__clkbuf_1 _5222_ (.A(_2133_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _5223_ (.A0(_1194_),
    .A1(\ih.gpio_interrupt_mask[6] ),
    .S(_2127_),
    .X(_2134_));
 sky130_fd_sc_hd__clkbuf_1 _5224_ (.A(_2134_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _5225_ (.A0(_1261_),
    .A1(\ih.gpio_interrupt_mask[7] ),
    .S(_2127_),
    .X(_2135_));
 sky130_fd_sc_hd__clkbuf_1 _5226_ (.A(_2135_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_4 _5227_ (.A(_1636_),
    .X(_2136_));
 sky130_fd_sc_hd__nor2_4 _5228_ (.A(_1415_),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__and2_1 _5229_ (.A(_1306_),
    .B(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__buf_2 _5230_ (.A(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__or3_2 _5231_ (.A(_1367_),
    .B(_1625_),
    .C(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__or2_1 _5232_ (.A(_1364_),
    .B(_1631_),
    .X(_2141_));
 sky130_fd_sc_hd__nor2_1 _5233_ (.A(_2140_),
    .B(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__mux2_1 _5234_ (.A0(\ih.t.enable ),
    .A1(_2085_),
    .S(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__clkbuf_1 _5235_ (.A(_2143_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _5236_ (.A0(_0617_),
    .A1(_1622_),
    .S(_1667_),
    .X(_2144_));
 sky130_fd_sc_hd__nor2_1 _5237_ (.A(_1369_),
    .B(_1625_),
    .Y(_2145_));
 sky130_fd_sc_hd__clkbuf_4 _5238_ (.A(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_8 _5239_ (.A(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__or2_2 _5240_ (.A(_1329_),
    .B(_1372_),
    .X(_2148_));
 sky130_fd_sc_hd__nor2_1 _5241_ (.A(_1374_),
    .B(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__or2_2 _5242_ (.A(_2145_),
    .B(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__buf_2 _5243_ (.A(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__o21ba_1 _5244_ (.A1(_1661_),
    .A2(_2151_),
    .B1_N(_2141_),
    .X(_2152_));
 sky130_fd_sc_hd__o21a_4 _5245_ (.A1(_1667_),
    .A2(_2147_),
    .B1(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__mux2_1 _5246_ (.A0(\ih.t.timer_max[24] ),
    .A1(_2144_),
    .S(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__clkbuf_1 _5247_ (.A(_2154_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(_1050_),
    .A1(_1623_),
    .S(_1667_),
    .X(_2155_));
 sky130_fd_sc_hd__mux2_1 _5249_ (.A0(\ih.t.timer_max[25] ),
    .A1(_2155_),
    .S(_2153_),
    .X(_2156_));
 sky130_fd_sc_hd__clkbuf_1 _5250_ (.A(_2156_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _5251_ (.A0(_1073_),
    .A1(_1226_),
    .S(_1667_),
    .X(_2157_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(\ih.t.timer_max[26] ),
    .A1(_2157_),
    .S(_2153_),
    .X(_2158_));
 sky130_fd_sc_hd__clkbuf_1 _5253_ (.A(_2158_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(_1089_),
    .A1(_1222_),
    .S(_1667_),
    .X(_2159_));
 sky130_fd_sc_hd__mux2_1 _5255_ (.A0(\ih.t.timer_max[27] ),
    .A1(_2159_),
    .S(_2153_),
    .X(_2160_));
 sky130_fd_sc_hd__clkbuf_1 _5256_ (.A(_2160_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(_1160_),
    .A1(_1213_),
    .S(_1667_),
    .X(_2161_));
 sky130_fd_sc_hd__mux2_1 _5258_ (.A0(\ih.t.timer_max[28] ),
    .A1(_2161_),
    .S(_2153_),
    .X(_2162_));
 sky130_fd_sc_hd__clkbuf_1 _5259_ (.A(_2162_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(_1144_),
    .A1(_1209_),
    .S(_1666_),
    .X(_2163_));
 sky130_fd_sc_hd__mux2_1 _5261_ (.A0(\ih.t.timer_max[29] ),
    .A1(_2163_),
    .S(_2153_),
    .X(_2164_));
 sky130_fd_sc_hd__clkbuf_1 _5262_ (.A(_2164_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(_1126_),
    .A1(_1624_),
    .S(_1666_),
    .X(_2165_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(\ih.t.timer_max[30] ),
    .A1(_2165_),
    .S(_2153_),
    .X(_2166_));
 sky130_fd_sc_hd__clkbuf_1 _5265_ (.A(_2166_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(_1110_),
    .A1(_1263_),
    .S(_1666_),
    .X(_2167_));
 sky130_fd_sc_hd__mux2_1 _5267_ (.A0(\ih.t.timer_max[31] ),
    .A1(_2167_),
    .S(_2153_),
    .X(_2168_));
 sky130_fd_sc_hd__clkbuf_1 _5268_ (.A(_2168_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_4 _5269_ (.A(_1642_),
    .X(_2169_));
 sky130_fd_sc_hd__nor2_4 _5270_ (.A(_2169_),
    .B(_2140_),
    .Y(_2170_));
 sky130_fd_sc_hd__mux2_1 _5271_ (.A0(net76),
    .A1(_2085_),
    .S(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__clkbuf_1 _5272_ (.A(_2171_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _5273_ (.A0(net77),
    .A1(_1051_),
    .S(_2170_),
    .X(_2172_));
 sky130_fd_sc_hd__clkbuf_1 _5274_ (.A(_2172_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _5275_ (.A0(net78),
    .A1(_1074_),
    .S(_2170_),
    .X(_2173_));
 sky130_fd_sc_hd__clkbuf_1 _5276_ (.A(_2173_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(net79),
    .A1(_1187_),
    .S(_2170_),
    .X(_2174_));
 sky130_fd_sc_hd__clkbuf_1 _5278_ (.A(_2174_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _5279_ (.A0(net80),
    .A1(_1189_),
    .S(_2170_),
    .X(_2175_));
 sky130_fd_sc_hd__clkbuf_1 _5280_ (.A(_2175_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(net81),
    .A1(_1191_),
    .S(_2170_),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_1 _5282_ (.A(_2176_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(net82),
    .A1(_1193_),
    .S(_2170_),
    .X(_2177_));
 sky130_fd_sc_hd__clkbuf_1 _5284_ (.A(_2177_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _5285_ (.A0(net83),
    .A1(_1260_),
    .S(_2170_),
    .X(_2178_));
 sky130_fd_sc_hd__clkbuf_1 _5286_ (.A(_2178_),
    .X(_0125_));
 sky130_fd_sc_hd__nor2_2 _5287_ (.A(_1329_),
    .B(_1354_),
    .Y(_2179_));
 sky130_fd_sc_hd__and2_4 _5288_ (.A(_1369_),
    .B(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__nor2_2 _5289_ (.A(_1364_),
    .B(_2169_),
    .Y(_2181_));
 sky130_fd_sc_hd__nand2_8 _5290_ (.A(_2180_),
    .B(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(_0619_),
    .A1(net84),
    .S(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__clkbuf_1 _5292_ (.A(_2183_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(_1052_),
    .A1(net85),
    .S(_2182_),
    .X(_2184_));
 sky130_fd_sc_hd__clkbuf_1 _5294_ (.A(_2184_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(_1075_),
    .A1(net86),
    .S(_2182_),
    .X(_2185_));
 sky130_fd_sc_hd__clkbuf_1 _5296_ (.A(_2185_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(_1188_),
    .A1(net87),
    .S(_2182_),
    .X(_2186_));
 sky130_fd_sc_hd__clkbuf_1 _5298_ (.A(_2186_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(_1190_),
    .A1(net88),
    .S(_2182_),
    .X(_2187_));
 sky130_fd_sc_hd__clkbuf_1 _5300_ (.A(_2187_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _5301_ (.A0(_1192_),
    .A1(net89),
    .S(_2182_),
    .X(_2188_));
 sky130_fd_sc_hd__clkbuf_1 _5302_ (.A(_2188_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(_1194_),
    .A1(net90),
    .S(_2182_),
    .X(_2189_));
 sky130_fd_sc_hd__clkbuf_1 _5304_ (.A(_2189_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(_1261_),
    .A1(net91),
    .S(_2182_),
    .X(_2190_));
 sky130_fd_sc_hd__clkbuf_1 _5306_ (.A(_2190_),
    .X(_0133_));
 sky130_fd_sc_hd__nand2_1 _5307_ (.A(_1329_),
    .B(_1354_),
    .Y(_2191_));
 sky130_fd_sc_hd__nor2_1 _5308_ (.A(_1374_),
    .B(_2191_),
    .Y(_2192_));
 sky130_fd_sc_hd__clkbuf_4 _5309_ (.A(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_8 _5310_ (.A(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__nand2_8 _5311_ (.A(net141),
    .B(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(_0619_),
    .A1(net92),
    .S(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__clkbuf_1 _5313_ (.A(_2196_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(_1052_),
    .A1(net93),
    .S(_2195_),
    .X(_2197_));
 sky130_fd_sc_hd__clkbuf_1 _5315_ (.A(_2197_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(_1075_),
    .A1(net94),
    .S(_2195_),
    .X(_2198_));
 sky130_fd_sc_hd__clkbuf_1 _5317_ (.A(_2198_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _5318_ (.A0(_1188_),
    .A1(net95),
    .S(_2195_),
    .X(_2199_));
 sky130_fd_sc_hd__clkbuf_1 _5319_ (.A(_2199_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _5320_ (.A0(_1190_),
    .A1(net96),
    .S(_2195_),
    .X(_2200_));
 sky130_fd_sc_hd__clkbuf_1 _5321_ (.A(_2200_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _5322_ (.A0(_1192_),
    .A1(net97),
    .S(_2195_),
    .X(_2201_));
 sky130_fd_sc_hd__clkbuf_1 _5323_ (.A(_2201_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(_1194_),
    .A1(net98),
    .S(_2195_),
    .X(_2202_));
 sky130_fd_sc_hd__clkbuf_1 _5325_ (.A(_2202_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _5326_ (.A0(_1261_),
    .A1(net99),
    .S(_2195_),
    .X(_2203_));
 sky130_fd_sc_hd__clkbuf_1 _5327_ (.A(_2203_),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_4 _5328_ (.A(_2149_),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_8 _5329_ (.A(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__nand2_8 _5330_ (.A(_2205_),
    .B(net141),
    .Y(_2206_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(_0619_),
    .A1(net100),
    .S(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_1 _5332_ (.A(_2207_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _5333_ (.A0(_1052_),
    .A1(net101),
    .S(_2206_),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_1 _5334_ (.A(_2208_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _5335_ (.A0(_1075_),
    .A1(net102),
    .S(_2206_),
    .X(_2209_));
 sky130_fd_sc_hd__clkbuf_1 _5336_ (.A(_2209_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(_1188_),
    .A1(net103),
    .S(_2206_),
    .X(_2210_));
 sky130_fd_sc_hd__clkbuf_1 _5338_ (.A(_2210_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _5339_ (.A0(_1190_),
    .A1(net104),
    .S(_2206_),
    .X(_2211_));
 sky130_fd_sc_hd__clkbuf_1 _5340_ (.A(_2211_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _5341_ (.A0(_1192_),
    .A1(net105),
    .S(_2206_),
    .X(_2212_));
 sky130_fd_sc_hd__clkbuf_1 _5342_ (.A(_2212_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(_1194_),
    .A1(net106),
    .S(_2206_),
    .X(_2213_));
 sky130_fd_sc_hd__clkbuf_1 _5344_ (.A(_2213_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(_1261_),
    .A1(net107),
    .S(_2206_),
    .X(_2214_));
 sky130_fd_sc_hd__clkbuf_1 _5346_ (.A(_2214_),
    .X(_0149_));
 sky130_fd_sc_hd__nand2_8 _5347_ (.A(_2147_),
    .B(net141),
    .Y(_2215_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(_0619_),
    .A1(net108),
    .S(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__clkbuf_1 _5349_ (.A(_2216_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(_1052_),
    .A1(net109),
    .S(_2215_),
    .X(_2217_));
 sky130_fd_sc_hd__clkbuf_1 _5351_ (.A(_2217_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _5352_ (.A0(_1075_),
    .A1(net110),
    .S(_2215_),
    .X(_2218_));
 sky130_fd_sc_hd__clkbuf_1 _5353_ (.A(_2218_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _5354_ (.A0(_1188_),
    .A1(net111),
    .S(_2215_),
    .X(_2219_));
 sky130_fd_sc_hd__clkbuf_1 _5355_ (.A(_2219_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(_1190_),
    .A1(net112),
    .S(_2215_),
    .X(_2220_));
 sky130_fd_sc_hd__clkbuf_1 _5357_ (.A(_2220_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _5358_ (.A0(_1192_),
    .A1(net113),
    .S(_2215_),
    .X(_2221_));
 sky130_fd_sc_hd__clkbuf_1 _5359_ (.A(_2221_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _5360_ (.A0(_1194_),
    .A1(net114),
    .S(_2215_),
    .X(_2222_));
 sky130_fd_sc_hd__clkbuf_1 _5361_ (.A(_2222_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(_1261_),
    .A1(net115),
    .S(_2215_),
    .X(_2223_));
 sky130_fd_sc_hd__clkbuf_1 _5363_ (.A(_2223_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _5364_ (.A(_1374_),
    .B(_2179_),
    .X(_2224_));
 sky130_fd_sc_hd__buf_4 _5365_ (.A(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__nand2_8 _5366_ (.A(net141),
    .B(_2225_),
    .Y(_2226_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(_0619_),
    .A1(net116),
    .S(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__clkbuf_1 _5368_ (.A(_2227_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(_1052_),
    .A1(net117),
    .S(_2226_),
    .X(_2228_));
 sky130_fd_sc_hd__clkbuf_1 _5370_ (.A(_2228_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(_1075_),
    .A1(net118),
    .S(_2226_),
    .X(_2229_));
 sky130_fd_sc_hd__clkbuf_1 _5372_ (.A(_2229_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(_1188_),
    .A1(net119),
    .S(_2226_),
    .X(_2230_));
 sky130_fd_sc_hd__clkbuf_1 _5374_ (.A(_2230_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(_1190_),
    .A1(net120),
    .S(_2226_),
    .X(_2231_));
 sky130_fd_sc_hd__clkbuf_1 _5376_ (.A(_2231_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(_1192_),
    .A1(net121),
    .S(_2226_),
    .X(_2232_));
 sky130_fd_sc_hd__clkbuf_1 _5378_ (.A(_2232_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5379_ (.A0(_1194_),
    .A1(net122),
    .S(_2226_),
    .X(_2233_));
 sky130_fd_sc_hd__clkbuf_1 _5380_ (.A(_2233_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(_1261_),
    .A1(net123),
    .S(_2226_),
    .X(_2234_));
 sky130_fd_sc_hd__clkbuf_1 _5382_ (.A(_2234_),
    .X(_0165_));
 sky130_fd_sc_hd__nor2_1 _5383_ (.A(_1369_),
    .B(_2191_),
    .Y(_2235_));
 sky130_fd_sc_hd__clkbuf_8 _5384_ (.A(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__nand2_8 _5385_ (.A(net141),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__mux2_1 _5386_ (.A0(_0619_),
    .A1(net124),
    .S(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__clkbuf_1 _5387_ (.A(_2238_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5388_ (.A0(_1052_),
    .A1(net125),
    .S(_2237_),
    .X(_2239_));
 sky130_fd_sc_hd__clkbuf_1 _5389_ (.A(_2239_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5390_ (.A0(_1075_),
    .A1(net126),
    .S(_2237_),
    .X(_2240_));
 sky130_fd_sc_hd__clkbuf_1 _5391_ (.A(_2240_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5392_ (.A0(_1188_),
    .A1(net127),
    .S(_2237_),
    .X(_2241_));
 sky130_fd_sc_hd__clkbuf_1 _5393_ (.A(_2241_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5394_ (.A0(_1190_),
    .A1(net128),
    .S(_2237_),
    .X(_2242_));
 sky130_fd_sc_hd__clkbuf_1 _5395_ (.A(_2242_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(_1192_),
    .A1(net129),
    .S(_2237_),
    .X(_2243_));
 sky130_fd_sc_hd__clkbuf_1 _5397_ (.A(_2243_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5398_ (.A0(_1194_),
    .A1(net130),
    .S(_2237_),
    .X(_2244_));
 sky130_fd_sc_hd__clkbuf_1 _5399_ (.A(_2244_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5400_ (.A0(_1261_),
    .A1(net131),
    .S(_2237_),
    .X(_2245_));
 sky130_fd_sc_hd__clkbuf_1 _5401_ (.A(_2245_),
    .X(_0173_));
 sky130_fd_sc_hd__nor2_1 _5402_ (.A(_1369_),
    .B(_2148_),
    .Y(_2246_));
 sky130_fd_sc_hd__clkbuf_8 _5403_ (.A(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__nand2_8 _5404_ (.A(net141),
    .B(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(_0619_),
    .A1(net132),
    .S(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__clkbuf_1 _5406_ (.A(_2249_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(_1052_),
    .A1(net133),
    .S(_2248_),
    .X(_2250_));
 sky130_fd_sc_hd__clkbuf_1 _5408_ (.A(_2250_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _5409_ (.A0(_1075_),
    .A1(net134),
    .S(_2248_),
    .X(_2251_));
 sky130_fd_sc_hd__clkbuf_1 _5410_ (.A(_2251_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(_1188_),
    .A1(net135),
    .S(_2248_),
    .X(_2252_));
 sky130_fd_sc_hd__clkbuf_1 _5412_ (.A(_2252_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _5413_ (.A0(_1190_),
    .A1(net136),
    .S(_2248_),
    .X(_2253_));
 sky130_fd_sc_hd__clkbuf_1 _5414_ (.A(_2253_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _5415_ (.A0(_1192_),
    .A1(net137),
    .S(_2248_),
    .X(_2254_));
 sky130_fd_sc_hd__clkbuf_1 _5416_ (.A(_2254_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _5417_ (.A0(_1194_),
    .A1(net138),
    .S(_2248_),
    .X(_2255_));
 sky130_fd_sc_hd__clkbuf_1 _5418_ (.A(_2255_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(_1261_),
    .A1(net139),
    .S(_2248_),
    .X(_2256_));
 sky130_fd_sc_hd__clkbuf_1 _5420_ (.A(_2256_),
    .X(_0181_));
 sky130_fd_sc_hd__and3_1 _5421_ (.A(_1329_),
    .B(_1372_),
    .C(_1369_),
    .X(_2257_));
 sky130_fd_sc_hd__and3_1 _5422_ (.A(_1306_),
    .B(_2257_),
    .C(_2137_),
    .X(_2258_));
 sky130_fd_sc_hd__mux2_1 _5423_ (.A0(net68),
    .A1(_2085_),
    .S(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__clkbuf_1 _5424_ (.A(_2259_),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _5425_ (.A(_2139_),
    .B(_2180_),
    .Y(_2260_));
 sky130_fd_sc_hd__mux2_1 _5426_ (.A0(_2022_),
    .A1(net69),
    .S(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__clkbuf_1 _5427_ (.A(_2261_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_2139_),
    .B(_2194_),
    .Y(_2262_));
 sky130_fd_sc_hd__mux2_1 _5429_ (.A0(_2022_),
    .A1(net70),
    .S(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__clkbuf_1 _5430_ (.A(_2263_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_2139_),
    .B(_2205_),
    .Y(_2264_));
 sky130_fd_sc_hd__mux2_1 _5432_ (.A0(_2022_),
    .A1(net71),
    .S(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__clkbuf_1 _5433_ (.A(_2265_),
    .X(_0185_));
 sky130_fd_sc_hd__nand2_1 _5434_ (.A(_2139_),
    .B(_2147_),
    .Y(_2266_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(_2022_),
    .A1(net72),
    .S(_2266_),
    .X(_2267_));
 sky130_fd_sc_hd__clkbuf_1 _5436_ (.A(_2267_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_2139_),
    .B(_2225_),
    .Y(_2268_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(_2022_),
    .A1(net73),
    .S(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__clkbuf_1 _5439_ (.A(_2269_),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(_2139_),
    .B(_2236_),
    .Y(_2270_));
 sky130_fd_sc_hd__mux2_1 _5441_ (.A0(_2022_),
    .A1(net74),
    .S(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__clkbuf_1 _5442_ (.A(_2271_),
    .X(_0188_));
 sky130_fd_sc_hd__nand2_1 _5443_ (.A(_2139_),
    .B(_2247_),
    .Y(_2272_));
 sky130_fd_sc_hd__mux2_1 _5444_ (.A0(_2022_),
    .A1(net75),
    .S(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__clkbuf_1 _5445_ (.A(_2273_),
    .X(_0189_));
 sky130_fd_sc_hd__buf_2 _5446_ (.A(_1640_),
    .X(_2274_));
 sky130_fd_sc_hd__or2_1 _5447_ (.A(_1417_),
    .B(_2136_),
    .X(_2275_));
 sky130_fd_sc_hd__mux4_1 _5448_ (.A0(net73),
    .A1(net75),
    .A2(net72),
    .A3(net74),
    .S0(_1354_),
    .S1(_1330_),
    .X(_2276_));
 sky130_fd_sc_hd__nor2_1 _5449_ (.A(_1335_),
    .B(_1354_),
    .Y(_2277_));
 sky130_fd_sc_hd__a22o_1 _5450_ (.A1(net68),
    .A2(_2277_),
    .B1(_2179_),
    .B2(net69),
    .X(_2278_));
 sky130_fd_sc_hd__nor2_1 _5451_ (.A(_1335_),
    .B(_1372_),
    .Y(_2279_));
 sky130_fd_sc_hd__a22o_1 _5452_ (.A1(net71),
    .A2(_1638_),
    .B1(_2279_),
    .B2(net70),
    .X(_2280_));
 sky130_fd_sc_hd__or3_1 _5453_ (.A(_1374_),
    .B(_2278_),
    .C(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__o21ai_1 _5454_ (.A1(_1369_),
    .A2(_2276_),
    .B1(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__or4_1 _5455_ (.A(_1364_),
    .B(_2274_),
    .C(_2275_),
    .D(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__buf_2 _5456_ (.A(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__nor2_1 _5457_ (.A(_1633_),
    .B(_2284_),
    .Y(_2285_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(net60),
    .A1(_2085_),
    .S(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__clkbuf_1 _5459_ (.A(_2286_),
    .X(_0190_));
 sky130_fd_sc_hd__nand2_1 _5460_ (.A(_1369_),
    .B(_2179_),
    .Y(_2287_));
 sky130_fd_sc_hd__nor2_1 _5461_ (.A(_2287_),
    .B(_2284_),
    .Y(_2288_));
 sky130_fd_sc_hd__mux2_1 _5462_ (.A0(net61),
    .A1(_2085_),
    .S(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__clkbuf_1 _5463_ (.A(_2289_),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _5464_ (.A(_2194_),
    .Y(_2290_));
 sky130_fd_sc_hd__nor2_1 _5465_ (.A(_2290_),
    .B(_2284_),
    .Y(_2291_));
 sky130_fd_sc_hd__mux2_1 _5466_ (.A0(net62),
    .A1(_2085_),
    .S(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__clkbuf_1 _5467_ (.A(_2292_),
    .X(_0192_));
 sky130_fd_sc_hd__inv_2 _5468_ (.A(_2205_),
    .Y(_2293_));
 sky130_fd_sc_hd__nor2_1 _5469_ (.A(_2293_),
    .B(_2284_),
    .Y(_2294_));
 sky130_fd_sc_hd__mux2_1 _5470_ (.A0(net63),
    .A1(_2085_),
    .S(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__clkbuf_1 _5471_ (.A(_2295_),
    .X(_0193_));
 sky130_fd_sc_hd__inv_2 _5472_ (.A(_2147_),
    .Y(_2296_));
 sky130_fd_sc_hd__nor2_1 _5473_ (.A(_2296_),
    .B(_2284_),
    .Y(_2297_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(net64),
    .A1(_2085_),
    .S(_2297_),
    .X(_2298_));
 sky130_fd_sc_hd__clkbuf_1 _5475_ (.A(_2298_),
    .X(_0194_));
 sky130_fd_sc_hd__inv_2 _5476_ (.A(_2225_),
    .Y(_2299_));
 sky130_fd_sc_hd__nor2_1 _5477_ (.A(_2299_),
    .B(_2284_),
    .Y(_2300_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(net65),
    .A1(_0618_),
    .S(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _5479_ (.A(_2301_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _5480_ (.A(_2236_),
    .Y(_2302_));
 sky130_fd_sc_hd__nor2_1 _5481_ (.A(_2302_),
    .B(_2284_),
    .Y(_2303_));
 sky130_fd_sc_hd__mux2_1 _5482_ (.A0(net66),
    .A1(_0618_),
    .S(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__clkbuf_1 _5483_ (.A(_2304_),
    .X(_0196_));
 sky130_fd_sc_hd__inv_2 _5484_ (.A(_2247_),
    .Y(_2305_));
 sky130_fd_sc_hd__nor2_1 _5485_ (.A(_2305_),
    .B(_2284_),
    .Y(_2306_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(net67),
    .A1(_0618_),
    .S(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__clkbuf_1 _5487_ (.A(_2307_),
    .X(_0197_));
 sky130_fd_sc_hd__a22o_1 _5488_ (.A1(net84),
    .A2(_2180_),
    .B1(_2224_),
    .B2(net116),
    .X(_2308_));
 sky130_fd_sc_hd__a221o_1 _5489_ (.A1(net124),
    .A2(_2236_),
    .B1(_2247_),
    .B2(net132),
    .C1(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__a22o_1 _5490_ (.A1(net108),
    .A2(_2146_),
    .B1(_2193_),
    .B2(net92),
    .X(_2310_));
 sky130_fd_sc_hd__a211o_1 _5491_ (.A1(net100),
    .A2(_2205_),
    .B1(_2310_),
    .C1(_2257_),
    .X(_2311_));
 sky130_fd_sc_hd__o22a_1 _5492_ (.A1(net76),
    .A2(_1633_),
    .B1(_2309_),
    .B2(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__and3_2 _5493_ (.A(\mc.cl.cmp_o ),
    .B(_1648_),
    .C(_1631_),
    .X(_2313_));
 sky130_fd_sc_hd__nor2_2 _5494_ (.A(_1400_),
    .B(_2287_),
    .Y(_2314_));
 sky130_fd_sc_hd__a22o_1 _5495_ (.A1(\ih.t.enable ),
    .A2(_2257_),
    .B1(_2192_),
    .B2(\ih.t.timer_max[8] ),
    .X(_2315_));
 sky130_fd_sc_hd__a22o_1 _5496_ (.A1(\ih.t.timer_max[24] ),
    .A2(_2146_),
    .B1(_2204_),
    .B2(\ih.t.timer_max[16] ),
    .X(_2316_));
 sky130_fd_sc_hd__nor2_1 _5497_ (.A(_2315_),
    .B(_2316_),
    .Y(_2317_));
 sky130_fd_sc_hd__o2bb2a_1 _5498_ (.A1_N(\ih.t.timer_max[0] ),
    .A2_N(_2314_),
    .B1(_2317_),
    .B2(_1400_),
    .X(_2318_));
 sky130_fd_sc_hd__or2_2 _5499_ (.A(_2180_),
    .B(_2193_),
    .X(_2319_));
 sky130_fd_sc_hd__buf_2 _5500_ (.A(_2319_),
    .X(_2320_));
 sky130_fd_sc_hd__a221o_1 _5501_ (.A1(\ih.t.enable ),
    .A2(_2257_),
    .B1(_2150_),
    .B2(\ih.t.timer_max[16] ),
    .C1(_1660_),
    .X(_2321_));
 sky130_fd_sc_hd__a21oi_1 _5502_ (.A1(\ih.t.timer_max[0] ),
    .A2(_2320_),
    .B1(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__a21oi_1 _5503_ (.A1(_1661_),
    .A2(_2318_),
    .B1(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__a2111oi_1 _5504_ (.A1(_1374_),
    .A2(_1625_),
    .B1(_1630_),
    .C1(_1489_),
    .D1(_1417_),
    .Y(_2324_));
 sky130_fd_sc_hd__a22o_1 _5505_ (.A1(\mc.cl.next_data[0] ),
    .A2(_2313_),
    .B1(_2323_),
    .B2(net237),
    .X(_2325_));
 sky130_fd_sc_hd__nor2_2 _5506_ (.A(_1489_),
    .B(_2125_),
    .Y(_2326_));
 sky130_fd_sc_hd__nor3_4 _5507_ (.A(_1415_),
    .B(_1629_),
    .C(_1637_),
    .Y(_2327_));
 sky130_fd_sc_hd__a221o_1 _5508_ (.A1(_2125_),
    .A2(_2325_),
    .B1(_2326_),
    .B2(\ih.gpio_interrupt_mask[0] ),
    .C1(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__o211a_1 _5509_ (.A1(_2169_),
    .A2(_2312_),
    .B1(_2328_),
    .C1(_2136_),
    .X(_2329_));
 sky130_fd_sc_hd__a31o_1 _5510_ (.A1(net68),
    .A2(_1648_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2330_));
 sky130_fd_sc_hd__a22o_1 _5511_ (.A1(net64),
    .A2(_2277_),
    .B1(_2179_),
    .B2(net65),
    .X(_2331_));
 sky130_fd_sc_hd__a22o_1 _5512_ (.A1(net67),
    .A2(_1638_),
    .B1(_2279_),
    .B2(net66),
    .X(_2332_));
 sky130_fd_sc_hd__a22o_1 _5513_ (.A1(net60),
    .A2(_2277_),
    .B1(_2179_),
    .B2(net61),
    .X(_2333_));
 sky130_fd_sc_hd__a22o_1 _5514_ (.A1(net63),
    .A2(_1638_),
    .B1(_2279_),
    .B2(net62),
    .X(_2334_));
 sky130_fd_sc_hd__or3_1 _5515_ (.A(_1374_),
    .B(_2333_),
    .C(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__o31a_1 _5516_ (.A1(_1369_),
    .A2(_2331_),
    .A3(_2332_),
    .B1(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__or3_1 _5517_ (.A(net32),
    .B(_1330_),
    .C(_1354_),
    .X(_2337_));
 sky130_fd_sc_hd__o21a_1 _5518_ (.A1(net33),
    .A2(_2191_),
    .B1(_1374_),
    .X(_2338_));
 sky130_fd_sc_hd__o22a_1 _5519_ (.A1(net31),
    .A2(_1625_),
    .B1(_2148_),
    .B2(net34),
    .X(_2339_));
 sky130_fd_sc_hd__mux4_1 _5520_ (.A0(net28),
    .A1(net30),
    .A2(net27),
    .A3(net29),
    .S0(_1354_),
    .S1(_1330_),
    .X(_2340_));
 sky130_fd_sc_hd__a32o_1 _5521_ (.A1(_2337_),
    .A2(_2338_),
    .A3(_2339_),
    .B1(_2340_),
    .B2(_1369_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(_2336_),
    .A1(_2341_),
    .S(_2282_),
    .X(_2342_));
 sky130_fd_sc_hd__and3b_1 _5523_ (.A_N(_2275_),
    .B(_2342_),
    .C(_1648_),
    .X(_2343_));
 sky130_fd_sc_hd__nand2_1 _5524_ (.A(_1666_),
    .B(_2191_),
    .Y(_2344_));
 sky130_fd_sc_hd__nand2_2 _5525_ (.A(_1625_),
    .B(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__a22o_1 _5526_ (.A1(net16),
    .A2(_2179_),
    .B1(_2279_),
    .B2(\ih.input_handler_enable ),
    .X(_2346_));
 sky130_fd_sc_hd__a21o_1 _5527_ (.A1(net2),
    .A2(_2345_),
    .B1(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _5528_ (.A0(net2),
    .A1(_2148_),
    .S(_2344_),
    .X(_2348_));
 sky130_fd_sc_hd__a31o_1 _5529_ (.A1(_1649_),
    .A2(_2347_),
    .A3(_2348_),
    .B1(_1641_),
    .X(_2349_));
 sky130_fd_sc_hd__o31a_2 _5530_ (.A1(_2329_),
    .A2(_2330_),
    .A3(_2343_),
    .B1(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__clkbuf_8 _5531_ (.A(_1739_),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(\cu.reg_file.reg_mem[0] ),
    .A1(_2350_),
    .S(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__clkbuf_1 _5533_ (.A(_2352_),
    .X(_0198_));
 sky130_fd_sc_hd__a22o_1 _5534_ (.A1(net125),
    .A2(_2236_),
    .B1(_2247_),
    .B2(net133),
    .X(_2353_));
 sky130_fd_sc_hd__a21o_1 _5535_ (.A1(net93),
    .A2(_2194_),
    .B1(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__or2_1 _5536_ (.A(net85),
    .B(_1330_),
    .X(_2355_));
 sky130_fd_sc_hd__a22o_1 _5537_ (.A1(net101),
    .A2(_2205_),
    .B1(_2355_),
    .B2(_1401_),
    .X(_2356_));
 sky130_fd_sc_hd__a221o_1 _5538_ (.A1(net109),
    .A2(_2147_),
    .B1(_2225_),
    .B2(net117),
    .C1(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__o22a_1 _5539_ (.A1(net77),
    .A2(_1633_),
    .B1(_2354_),
    .B2(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__buf_2 _5540_ (.A(_2313_),
    .X(_2359_));
 sky130_fd_sc_hd__a22o_1 _5541_ (.A1(\ih.t.timer_max[25] ),
    .A2(_2146_),
    .B1(_2204_),
    .B2(\ih.t.timer_max[17] ),
    .X(_2360_));
 sky130_fd_sc_hd__a221o_1 _5542_ (.A1(\ih.t.timer_max[9] ),
    .A2(_2193_),
    .B1(_2314_),
    .B2(\ih.t.timer_max[1] ),
    .C1(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__and2b_1 _5543_ (.A_N(_1400_),
    .B(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__a221o_1 _5544_ (.A1(\ih.t.timer_max[17] ),
    .A2(_2151_),
    .B1(_2319_),
    .B2(\ih.t.timer_max[1] ),
    .C1(_1661_),
    .X(_2363_));
 sky130_fd_sc_hd__o21a_1 _5545_ (.A1(_1666_),
    .A2(_2362_),
    .B1(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__a22o_1 _5546_ (.A1(\mc.cl.next_data[1] ),
    .A2(_2359_),
    .B1(_2324_),
    .B2(_2364_),
    .X(_2365_));
 sky130_fd_sc_hd__a221o_1 _5547_ (.A1(\ih.gpio_interrupt_mask[1] ),
    .A2(_2326_),
    .B1(_2365_),
    .B2(_2125_),
    .C1(_2327_),
    .X(_2366_));
 sky130_fd_sc_hd__o211a_1 _5548_ (.A1(_2169_),
    .A2(_2358_),
    .B1(_2366_),
    .C1(_2136_),
    .X(_2367_));
 sky130_fd_sc_hd__a31o_1 _5549_ (.A1(net69),
    .A2(_1649_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2368_));
 sky130_fd_sc_hd__and3_2 _5550_ (.A(_1335_),
    .B(_1372_),
    .C(_1661_),
    .X(_2369_));
 sky130_fd_sc_hd__a22o_1 _5551_ (.A1(net9),
    .A2(_2345_),
    .B1(_2369_),
    .B2(net17),
    .X(_2370_));
 sky130_fd_sc_hd__and2_1 _5552_ (.A(_1649_),
    .B(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__o22a_2 _5553_ (.A1(_2367_),
    .A2(_2368_),
    .B1(_2371_),
    .B2(_1641_),
    .X(_2372_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(\cu.reg_file.reg_mem[1] ),
    .A1(_2372_),
    .S(_2351_),
    .X(_2373_));
 sky130_fd_sc_hd__clkbuf_1 _5555_ (.A(_2373_),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_1 _5556_ (.A1(net126),
    .A2(_2236_),
    .B1(_2247_),
    .B2(net134),
    .X(_2374_));
 sky130_fd_sc_hd__a21o_1 _5557_ (.A1(net94),
    .A2(_2194_),
    .B1(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__or2_1 _5558_ (.A(net86),
    .B(_1330_),
    .X(_2376_));
 sky130_fd_sc_hd__a22o_1 _5559_ (.A1(net102),
    .A2(_2205_),
    .B1(_2376_),
    .B2(_1401_),
    .X(_2377_));
 sky130_fd_sc_hd__a221o_1 _5560_ (.A1(net110),
    .A2(_2147_),
    .B1(_2225_),
    .B2(net118),
    .C1(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__o22a_1 _5561_ (.A1(net78),
    .A2(_1633_),
    .B1(_2375_),
    .B2(_2378_),
    .X(_2379_));
 sky130_fd_sc_hd__a22o_1 _5562_ (.A1(\ih.t.timer_max[26] ),
    .A2(_2146_),
    .B1(_2204_),
    .B2(\ih.t.timer_max[18] ),
    .X(_2380_));
 sky130_fd_sc_hd__a221o_1 _5563_ (.A1(\ih.t.timer_max[10] ),
    .A2(_2193_),
    .B1(_2314_),
    .B2(\ih.t.timer_max[2] ),
    .C1(_2380_),
    .X(_2381_));
 sky130_fd_sc_hd__and2b_1 _5564_ (.A_N(_1400_),
    .B(_2381_),
    .X(_2382_));
 sky130_fd_sc_hd__a221o_1 _5565_ (.A1(\ih.t.timer_max[18] ),
    .A2(_2150_),
    .B1(_2319_),
    .B2(\ih.t.timer_max[2] ),
    .C1(_1661_),
    .X(_2383_));
 sky130_fd_sc_hd__o21a_1 _5566_ (.A1(_1666_),
    .A2(_2382_),
    .B1(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__a22o_1 _5567_ (.A1(\mc.cl.next_data[2] ),
    .A2(_2359_),
    .B1(net237),
    .B2(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__a221o_1 _5568_ (.A1(\ih.gpio_interrupt_mask[2] ),
    .A2(_2326_),
    .B1(_2385_),
    .B2(_2125_),
    .C1(_2327_),
    .X(_2386_));
 sky130_fd_sc_hd__o211a_1 _5569_ (.A1(_2169_),
    .A2(_2379_),
    .B1(_2386_),
    .C1(_2136_),
    .X(_2387_));
 sky130_fd_sc_hd__a31o_1 _5570_ (.A1(net70),
    .A2(_1648_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2388_));
 sky130_fd_sc_hd__a22o_1 _5571_ (.A1(net10),
    .A2(_2345_),
    .B1(_2369_),
    .B2(net3),
    .X(_2389_));
 sky130_fd_sc_hd__and2_1 _5572_ (.A(_1649_),
    .B(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__o22a_2 _5573_ (.A1(_2387_),
    .A2(_2388_),
    .B1(_2390_),
    .B2(_1641_),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(\cu.reg_file.reg_mem[2] ),
    .A1(_2391_),
    .S(_2351_),
    .X(_2392_));
 sky130_fd_sc_hd__clkbuf_1 _5575_ (.A(_2392_),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _5576_ (.A1(net127),
    .A2(_2236_),
    .B1(_2247_),
    .B2(net135),
    .X(_2393_));
 sky130_fd_sc_hd__a21o_1 _5577_ (.A1(net95),
    .A2(_2194_),
    .B1(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__or2_1 _5578_ (.A(net87),
    .B(_1330_),
    .X(_2395_));
 sky130_fd_sc_hd__a22o_1 _5579_ (.A1(net103),
    .A2(_2205_),
    .B1(_2395_),
    .B2(_1401_),
    .X(_2396_));
 sky130_fd_sc_hd__a221o_1 _5580_ (.A1(net111),
    .A2(_2147_),
    .B1(_2225_),
    .B2(net119),
    .C1(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__o22a_1 _5581_ (.A1(net79),
    .A2(_1633_),
    .B1(_2394_),
    .B2(_2397_),
    .X(_2398_));
 sky130_fd_sc_hd__a22o_1 _5582_ (.A1(\ih.t.timer_max[27] ),
    .A2(_2146_),
    .B1(_2204_),
    .B2(\ih.t.timer_max[19] ),
    .X(_2399_));
 sky130_fd_sc_hd__a221o_1 _5583_ (.A1(\ih.t.timer_max[11] ),
    .A2(_2193_),
    .B1(_2314_),
    .B2(\ih.t.timer_max[3] ),
    .C1(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__and2b_1 _5584_ (.A_N(_1400_),
    .B(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__a221o_1 _5585_ (.A1(\ih.t.timer_max[19] ),
    .A2(_2150_),
    .B1(_2319_),
    .B2(\ih.t.timer_max[3] ),
    .C1(_1661_),
    .X(_2402_));
 sky130_fd_sc_hd__o21a_1 _5586_ (.A1(_1666_),
    .A2(_2401_),
    .B1(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__a22o_1 _5587_ (.A1(\mc.cl.next_data[3] ),
    .A2(_2313_),
    .B1(net142),
    .B2(_2403_),
    .X(_2404_));
 sky130_fd_sc_hd__a221o_1 _5588_ (.A1(\ih.gpio_interrupt_mask[3] ),
    .A2(_2326_),
    .B1(_2404_),
    .B2(_2125_),
    .C1(_2327_),
    .X(_2405_));
 sky130_fd_sc_hd__o211a_1 _5589_ (.A1(_2169_),
    .A2(_2398_),
    .B1(_2405_),
    .C1(_2136_),
    .X(_2406_));
 sky130_fd_sc_hd__a31o_1 _5590_ (.A1(net71),
    .A2(_1648_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2407_));
 sky130_fd_sc_hd__a22o_1 _5591_ (.A1(net11),
    .A2(_2345_),
    .B1(_2369_),
    .B2(net4),
    .X(_2408_));
 sky130_fd_sc_hd__and2_1 _5592_ (.A(_1649_),
    .B(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__o22a_2 _5593_ (.A1(_2406_),
    .A2(_2407_),
    .B1(_2409_),
    .B2(_1641_),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(\cu.reg_file.reg_mem[3] ),
    .A1(_2410_),
    .S(_2351_),
    .X(_2411_));
 sky130_fd_sc_hd__clkbuf_1 _5595_ (.A(_2411_),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_1 _5596_ (.A1(net128),
    .A2(_2236_),
    .B1(_2247_),
    .B2(net136),
    .X(_2412_));
 sky130_fd_sc_hd__a21o_1 _5597_ (.A1(net96),
    .A2(_2194_),
    .B1(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__or2_1 _5598_ (.A(net88),
    .B(_1330_),
    .X(_2414_));
 sky130_fd_sc_hd__a22o_1 _5599_ (.A1(net104),
    .A2(_2205_),
    .B1(_2414_),
    .B2(_1401_),
    .X(_2415_));
 sky130_fd_sc_hd__a221o_1 _5600_ (.A1(net112),
    .A2(_2147_),
    .B1(_2225_),
    .B2(net120),
    .C1(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__o22a_1 _5601_ (.A1(net80),
    .A2(_1633_),
    .B1(_2413_),
    .B2(_2416_),
    .X(_2417_));
 sky130_fd_sc_hd__a22o_1 _5602_ (.A1(\ih.t.timer_max[28] ),
    .A2(_2146_),
    .B1(_2204_),
    .B2(\ih.t.timer_max[20] ),
    .X(_2418_));
 sky130_fd_sc_hd__a221o_1 _5603_ (.A1(\ih.t.timer_max[12] ),
    .A2(_2193_),
    .B1(_2314_),
    .B2(\ih.t.timer_max[4] ),
    .C1(_2418_),
    .X(_2419_));
 sky130_fd_sc_hd__and2b_1 _5604_ (.A_N(_1400_),
    .B(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__a221o_1 _5605_ (.A1(\ih.t.timer_max[20] ),
    .A2(_2150_),
    .B1(_2319_),
    .B2(\ih.t.timer_max[4] ),
    .C1(_1661_),
    .X(_2421_));
 sky130_fd_sc_hd__o21a_1 _5606_ (.A1(_1666_),
    .A2(_2420_),
    .B1(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__a22o_1 _5607_ (.A1(\mc.cl.next_data[4] ),
    .A2(_2313_),
    .B1(net142),
    .B2(_2422_),
    .X(_2423_));
 sky130_fd_sc_hd__a221o_1 _5608_ (.A1(\ih.gpio_interrupt_mask[4] ),
    .A2(_2326_),
    .B1(_2423_),
    .B2(_2125_),
    .C1(_2327_),
    .X(_2424_));
 sky130_fd_sc_hd__o211a_1 _5609_ (.A1(_2169_),
    .A2(_2417_),
    .B1(_2424_),
    .C1(_2136_),
    .X(_2425_));
 sky130_fd_sc_hd__a31o_1 _5610_ (.A1(net72),
    .A2(_1648_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2426_));
 sky130_fd_sc_hd__a22o_1 _5611_ (.A1(net12),
    .A2(_2345_),
    .B1(_2369_),
    .B2(net5),
    .X(_2427_));
 sky130_fd_sc_hd__and2_1 _5612_ (.A(_1649_),
    .B(_2427_),
    .X(_2428_));
 sky130_fd_sc_hd__o22a_2 _5613_ (.A1(_2425_),
    .A2(_2426_),
    .B1(_2428_),
    .B2(_1641_),
    .X(_2429_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(\cu.reg_file.reg_mem[4] ),
    .A1(_2429_),
    .S(_2351_),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_1 _5615_ (.A(_2430_),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_1 _5616_ (.A1(net129),
    .A2(_2236_),
    .B1(_2247_),
    .B2(net137),
    .X(_2431_));
 sky130_fd_sc_hd__a21o_1 _5617_ (.A1(net97),
    .A2(_2194_),
    .B1(_2431_),
    .X(_2432_));
 sky130_fd_sc_hd__or2_1 _5618_ (.A(net89),
    .B(_1330_),
    .X(_2433_));
 sky130_fd_sc_hd__a22o_1 _5619_ (.A1(net105),
    .A2(_2205_),
    .B1(_2433_),
    .B2(_1401_),
    .X(_2434_));
 sky130_fd_sc_hd__a221o_1 _5620_ (.A1(net113),
    .A2(_2147_),
    .B1(_2225_),
    .B2(net121),
    .C1(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__o22a_1 _5621_ (.A1(net81),
    .A2(_1633_),
    .B1(_2432_),
    .B2(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__a22o_1 _5622_ (.A1(\ih.t.timer_max[29] ),
    .A2(_2146_),
    .B1(_2204_),
    .B2(\ih.t.timer_max[21] ),
    .X(_2437_));
 sky130_fd_sc_hd__a221o_1 _5623_ (.A1(\ih.t.timer_max[13] ),
    .A2(_2193_),
    .B1(_2314_),
    .B2(\ih.t.timer_max[5] ),
    .C1(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__and2b_1 _5624_ (.A_N(_1400_),
    .B(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__a221o_1 _5625_ (.A1(\ih.t.timer_max[21] ),
    .A2(_2150_),
    .B1(_2319_),
    .B2(\ih.t.timer_max[5] ),
    .C1(_1661_),
    .X(_2440_));
 sky130_fd_sc_hd__o21a_1 _5626_ (.A1(_1666_),
    .A2(_2439_),
    .B1(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__a22o_1 _5627_ (.A1(\mc.cl.next_data[5] ),
    .A2(_2313_),
    .B1(net142),
    .B2(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__a221o_1 _5628_ (.A1(\ih.gpio_interrupt_mask[5] ),
    .A2(_2326_),
    .B1(_2442_),
    .B2(_2125_),
    .C1(_2327_),
    .X(_2443_));
 sky130_fd_sc_hd__o211a_1 _5629_ (.A1(_2169_),
    .A2(_2436_),
    .B1(_2443_),
    .C1(_2136_),
    .X(_2444_));
 sky130_fd_sc_hd__a31o_1 _5630_ (.A1(net73),
    .A2(_1648_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2445_));
 sky130_fd_sc_hd__a22o_1 _5631_ (.A1(net13),
    .A2(_2345_),
    .B1(_2369_),
    .B2(net6),
    .X(_2446_));
 sky130_fd_sc_hd__and2_1 _5632_ (.A(_1649_),
    .B(_2446_),
    .X(_2447_));
 sky130_fd_sc_hd__o22a_4 _5633_ (.A1(_2444_),
    .A2(_2445_),
    .B1(_2447_),
    .B2(_1641_),
    .X(_2448_));
 sky130_fd_sc_hd__mux2_1 _5634_ (.A0(\cu.reg_file.reg_mem[5] ),
    .A1(_2448_),
    .S(_2351_),
    .X(_2449_));
 sky130_fd_sc_hd__clkbuf_1 _5635_ (.A(_2449_),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_1 _5636_ (.A1(net130),
    .A2(_2236_),
    .B1(_2247_),
    .B2(net138),
    .X(_2450_));
 sky130_fd_sc_hd__a21o_1 _5637_ (.A1(net98),
    .A2(_2194_),
    .B1(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__or2_1 _5638_ (.A(net90),
    .B(_1330_),
    .X(_2452_));
 sky130_fd_sc_hd__a22o_1 _5639_ (.A1(net106),
    .A2(_2204_),
    .B1(_2452_),
    .B2(_1401_),
    .X(_2453_));
 sky130_fd_sc_hd__a221o_1 _5640_ (.A1(net114),
    .A2(_2147_),
    .B1(_2225_),
    .B2(net122),
    .C1(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__o22a_1 _5641_ (.A1(net82),
    .A2(_1633_),
    .B1(_2451_),
    .B2(_2454_),
    .X(_2455_));
 sky130_fd_sc_hd__a22o_1 _5642_ (.A1(\ih.t.timer_max[30] ),
    .A2(_2146_),
    .B1(_2149_),
    .B2(\ih.t.timer_max[22] ),
    .X(_2456_));
 sky130_fd_sc_hd__a221o_1 _5643_ (.A1(\ih.t.timer_max[14] ),
    .A2(_2193_),
    .B1(_2314_),
    .B2(\ih.t.timer_max[6] ),
    .C1(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__and2b_1 _5644_ (.A_N(_1400_),
    .B(_2457_),
    .X(_2458_));
 sky130_fd_sc_hd__a221o_1 _5645_ (.A1(\ih.t.timer_max[22] ),
    .A2(_2150_),
    .B1(_2319_),
    .B2(\ih.t.timer_max[6] ),
    .C1(_1660_),
    .X(_2459_));
 sky130_fd_sc_hd__o21a_1 _5646_ (.A1(_1665_),
    .A2(_2458_),
    .B1(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__a22o_1 _5647_ (.A1(\mc.cl.next_data[6] ),
    .A2(_2313_),
    .B1(net142),
    .B2(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__a221o_1 _5648_ (.A1(\ih.gpio_interrupt_mask[6] ),
    .A2(_2326_),
    .B1(_2461_),
    .B2(_2125_),
    .C1(_2327_),
    .X(_2462_));
 sky130_fd_sc_hd__o211a_1 _5649_ (.A1(_2169_),
    .A2(_2455_),
    .B1(_2462_),
    .C1(_2136_),
    .X(_2463_));
 sky130_fd_sc_hd__a31o_1 _5650_ (.A1(net74),
    .A2(_1648_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2464_));
 sky130_fd_sc_hd__a22o_1 _5651_ (.A1(net14),
    .A2(_2345_),
    .B1(_2369_),
    .B2(net7),
    .X(_2465_));
 sky130_fd_sc_hd__and2_1 _5652_ (.A(_1649_),
    .B(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__o22a_4 _5653_ (.A1(_2463_),
    .A2(_2464_),
    .B1(_2466_),
    .B2(_1641_),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(\cu.reg_file.reg_mem[6] ),
    .A1(_2467_),
    .S(_1739_),
    .X(_2468_));
 sky130_fd_sc_hd__clkbuf_1 _5655_ (.A(_2468_),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_1 _5656_ (.A1(net131),
    .A2(_2235_),
    .B1(_2246_),
    .B2(net139),
    .X(_2469_));
 sky130_fd_sc_hd__a21o_1 _5657_ (.A1(net99),
    .A2(_2193_),
    .B1(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__or2_1 _5658_ (.A(net91),
    .B(_1329_),
    .X(_2471_));
 sky130_fd_sc_hd__a22o_1 _5659_ (.A1(net107),
    .A2(_2204_),
    .B1(_2471_),
    .B2(_1401_),
    .X(_2472_));
 sky130_fd_sc_hd__a221o_1 _5660_ (.A1(net115),
    .A2(_2146_),
    .B1(_2225_),
    .B2(net123),
    .C1(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__o22a_1 _5661_ (.A1(net83),
    .A2(_1633_),
    .B1(_2470_),
    .B2(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__a22o_1 _5662_ (.A1(\ih.t.timer_max[31] ),
    .A2(_2145_),
    .B1(_2192_),
    .B2(\ih.t.timer_max[15] ),
    .X(_2475_));
 sky130_fd_sc_hd__a221o_1 _5663_ (.A1(\ih.t.timer_max[23] ),
    .A2(_2204_),
    .B1(_2314_),
    .B2(\ih.t.timer_max[7] ),
    .C1(_2475_),
    .X(_2476_));
 sky130_fd_sc_hd__and2b_1 _5664_ (.A_N(_1400_),
    .B(_2476_),
    .X(_2477_));
 sky130_fd_sc_hd__a221o_1 _5665_ (.A1(\ih.t.timer_max[23] ),
    .A2(_2150_),
    .B1(_2319_),
    .B2(\ih.t.timer_max[7] ),
    .C1(_1660_),
    .X(_2478_));
 sky130_fd_sc_hd__o21a_1 _5666_ (.A1(_1665_),
    .A2(_2477_),
    .B1(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__a22o_1 _5667_ (.A1(\mc.cl.next_data[7] ),
    .A2(_2313_),
    .B1(net142),
    .B2(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__a221o_1 _5668_ (.A1(\ih.gpio_interrupt_mask[7] ),
    .A2(_2326_),
    .B1(_2480_),
    .B2(_2125_),
    .C1(_2327_),
    .X(_2481_));
 sky130_fd_sc_hd__o211a_1 _5669_ (.A1(_2169_),
    .A2(_2474_),
    .B1(_2481_),
    .C1(_2136_),
    .X(_2482_));
 sky130_fd_sc_hd__a31o_1 _5670_ (.A1(net75),
    .A2(_1648_),
    .A3(_2137_),
    .B1(_2274_),
    .X(_2483_));
 sky130_fd_sc_hd__a22o_1 _5671_ (.A1(net15),
    .A2(_2345_),
    .B1(_2369_),
    .B2(net8),
    .X(_2484_));
 sky130_fd_sc_hd__and2_1 _5672_ (.A(_1649_),
    .B(_2484_),
    .X(_2485_));
 sky130_fd_sc_hd__o22a_4 _5673_ (.A1(_2482_),
    .A2(_2483_),
    .B1(_2485_),
    .B2(_1641_),
    .X(_2486_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(\cu.reg_file.reg_mem[7] ),
    .A1(_2486_),
    .S(_1739_),
    .X(_2487_));
 sky130_fd_sc_hd__clkbuf_1 _5675_ (.A(_2487_),
    .X(_0205_));
 sky130_fd_sc_hd__nor2_2 _5676_ (.A(_1641_),
    .B(_2344_),
    .Y(_2488_));
 sky130_fd_sc_hd__a22oi_1 _5677_ (.A1(\ih.t.timer_max[24] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[8] ),
    .Y(_2489_));
 sky130_fd_sc_hd__or3_2 _5678_ (.A(_1489_),
    .B(_1631_),
    .C(_1661_),
    .X(_2490_));
 sky130_fd_sc_hd__o2bb2a_1 _5679_ (.A1_N(\mc.cl.next_data[8] ),
    .A2_N(_2359_),
    .B1(_2489_),
    .B2(_2490_),
    .X(_2491_));
 sky130_fd_sc_hd__a2bb2o_1 _5680_ (.A1_N(_2491_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[8] ),
    .B2(_2111_),
    .X(_2492_));
 sky130_fd_sc_hd__a31o_1 _5681_ (.A1(net16),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2492_),
    .X(_0206_));
 sky130_fd_sc_hd__a22oi_1 _5682_ (.A1(\ih.t.timer_max[25] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[9] ),
    .Y(_2493_));
 sky130_fd_sc_hd__o2bb2a_1 _5683_ (.A1_N(\mc.cl.next_data[9] ),
    .A2_N(_2359_),
    .B1(_2490_),
    .B2(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__a2bb2o_1 _5684_ (.A1_N(_2494_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[9] ),
    .B2(_1646_),
    .X(_2495_));
 sky130_fd_sc_hd__a31o_1 _5685_ (.A1(net17),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2495_),
    .X(_0207_));
 sky130_fd_sc_hd__a22oi_1 _5686_ (.A1(\ih.t.timer_max[26] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[10] ),
    .Y(_2496_));
 sky130_fd_sc_hd__o2bb2a_1 _5687_ (.A1_N(\mc.cl.next_data[10] ),
    .A2_N(_2359_),
    .B1(_2490_),
    .B2(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__a2bb2o_1 _5688_ (.A1_N(_2497_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[10] ),
    .B2(_1646_),
    .X(_2498_));
 sky130_fd_sc_hd__a31o_1 _5689_ (.A1(net3),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2498_),
    .X(_0208_));
 sky130_fd_sc_hd__a22oi_1 _5690_ (.A1(\ih.t.timer_max[27] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[11] ),
    .Y(_2499_));
 sky130_fd_sc_hd__o2bb2a_1 _5691_ (.A1_N(\mc.cl.next_data[11] ),
    .A2_N(_2359_),
    .B1(_2490_),
    .B2(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__a2bb2o_1 _5692_ (.A1_N(_2500_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[11] ),
    .B2(_1646_),
    .X(_2501_));
 sky130_fd_sc_hd__a31o_1 _5693_ (.A1(net4),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2501_),
    .X(_0209_));
 sky130_fd_sc_hd__a22oi_1 _5694_ (.A1(\ih.t.timer_max[28] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[12] ),
    .Y(_2502_));
 sky130_fd_sc_hd__o2bb2a_1 _5695_ (.A1_N(\mc.cl.next_data[12] ),
    .A2_N(_2359_),
    .B1(_2490_),
    .B2(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__a2bb2o_1 _5696_ (.A1_N(_2503_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[12] ),
    .B2(_1646_),
    .X(_2504_));
 sky130_fd_sc_hd__a31o_1 _5697_ (.A1(net5),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2504_),
    .X(_0210_));
 sky130_fd_sc_hd__a22oi_1 _5698_ (.A1(\ih.t.timer_max[29] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[13] ),
    .Y(_2505_));
 sky130_fd_sc_hd__o2bb2a_1 _5699_ (.A1_N(\mc.cl.next_data[13] ),
    .A2_N(_2359_),
    .B1(_2490_),
    .B2(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__a2bb2o_1 _5700_ (.A1_N(_2506_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[13] ),
    .B2(_1646_),
    .X(_2507_));
 sky130_fd_sc_hd__a31o_1 _5701_ (.A1(net6),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2507_),
    .X(_0211_));
 sky130_fd_sc_hd__a22oi_1 _5702_ (.A1(\ih.t.timer_max[30] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[14] ),
    .Y(_2508_));
 sky130_fd_sc_hd__o2bb2a_1 _5703_ (.A1_N(\mc.cl.next_data[14] ),
    .A2_N(_2359_),
    .B1(_2490_),
    .B2(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__a2bb2o_1 _5704_ (.A1_N(_2509_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[14] ),
    .B2(_1646_),
    .X(_2510_));
 sky130_fd_sc_hd__a31o_1 _5705_ (.A1(net7),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2510_),
    .X(_0212_));
 sky130_fd_sc_hd__a22oi_1 _5706_ (.A1(\ih.t.timer_max[31] ),
    .A2(_2151_),
    .B1(_2320_),
    .B2(\ih.t.timer_max[15] ),
    .Y(_2511_));
 sky130_fd_sc_hd__o2bb2a_1 _5707_ (.A1_N(\mc.cl.next_data[15] ),
    .A2_N(_2359_),
    .B1(_2490_),
    .B2(_2511_),
    .X(_2512_));
 sky130_fd_sc_hd__a2bb2o_1 _5708_ (.A1_N(_2512_),
    .A2_N(_1643_),
    .B1(\cu.reg_file.reg_mem[15] ),
    .B2(_1646_),
    .X(_2513_));
 sky130_fd_sc_hd__a31o_1 _5709_ (.A1(net8),
    .A2(_1650_),
    .A3(_2488_),
    .B1(_2513_),
    .X(_0213_));
 sky130_fd_sc_hd__nor2_1 _5710_ (.A(_2708_),
    .B(_1653_),
    .Y(_2514_));
 sky130_fd_sc_hd__and2b_1 _5711_ (.A_N(net190),
    .B(\mc.cl.cmp_o ),
    .X(_2515_));
 sky130_fd_sc_hd__a31o_1 _5712_ (.A1(net190),
    .A2(_2707_),
    .A3(_2514_),
    .B1(_2515_),
    .X(_0214_));
 sky130_fd_sc_hd__and3_1 _5713_ (.A(_1328_),
    .B(_1354_),
    .C(_2274_),
    .X(_2516_));
 sky130_fd_sc_hd__mux2_1 _5714_ (.A0(\ih.input_handler_enable ),
    .A1(_0618_),
    .S(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__clkbuf_1 _5715_ (.A(_2517_),
    .X(_0215_));
 sky130_fd_sc_hd__buf_2 _5716_ (.A(\mc.count ),
    .X(_2518_));
 sky130_fd_sc_hd__nor2_4 _5717_ (.A(_2518_),
    .B(_2351_),
    .Y(_2519_));
 sky130_fd_sc_hd__nor2_1 _5718_ (.A(_2351_),
    .B(_2514_),
    .Y(_2520_));
 sky130_fd_sc_hd__a22o_1 _5719_ (.A1(_2514_),
    .A2(_2519_),
    .B1(_2520_),
    .B2(_2518_),
    .X(_0216_));
 sky130_fd_sc_hd__nor2_1 _5720_ (.A(net1),
    .B(\ih.interrupt_source[3] ),
    .Y(_2521_));
 sky130_fd_sc_hd__a2111oi_1 _5721_ (.A1(net1),
    .A2(net198),
    .B1(_2872_),
    .C1(_2870_),
    .D1(_2521_),
    .Y(_0217_));
 sky130_fd_sc_hd__a22o_1 _5722_ (.A1(_2869_),
    .A2(_2870_),
    .B1(_2873_),
    .B2(net205),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _5723_ (.A(_2518_),
    .B(\mc.cl.next_data[0] ),
    .C(_2111_),
    .X(_2522_));
 sky130_fd_sc_hd__a21o_1 _5724_ (.A1(net18),
    .A2(_2519_),
    .B1(_2522_),
    .X(_0219_));
 sky130_fd_sc_hd__and3_1 _5725_ (.A(_2518_),
    .B(\mc.cl.next_data[1] ),
    .C(_2111_),
    .X(_2523_));
 sky130_fd_sc_hd__a21o_1 _5726_ (.A1(net19),
    .A2(_2519_),
    .B1(_2523_),
    .X(_0220_));
 sky130_fd_sc_hd__and3_1 _5727_ (.A(_2518_),
    .B(\mc.cl.next_data[2] ),
    .C(_2111_),
    .X(_2524_));
 sky130_fd_sc_hd__a21o_1 _5728_ (.A1(net20),
    .A2(_2519_),
    .B1(_2524_),
    .X(_0221_));
 sky130_fd_sc_hd__and3_1 _5729_ (.A(_2518_),
    .B(\mc.cl.next_data[3] ),
    .C(_2111_),
    .X(_2525_));
 sky130_fd_sc_hd__a21o_1 _5730_ (.A1(net21),
    .A2(_2519_),
    .B1(_2525_),
    .X(_0222_));
 sky130_fd_sc_hd__and3_1 _5731_ (.A(_2518_),
    .B(\mc.cl.next_data[4] ),
    .C(_2111_),
    .X(_2526_));
 sky130_fd_sc_hd__a21o_1 _5732_ (.A1(net22),
    .A2(_2519_),
    .B1(_2526_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _5733_ (.A(_2518_),
    .B(\mc.cl.next_data[5] ),
    .C(_2111_),
    .X(_2527_));
 sky130_fd_sc_hd__a21o_1 _5734_ (.A1(net23),
    .A2(_2519_),
    .B1(_2527_),
    .X(_0224_));
 sky130_fd_sc_hd__and3_1 _5735_ (.A(_2518_),
    .B(\mc.cl.next_data[6] ),
    .C(_2111_),
    .X(_2528_));
 sky130_fd_sc_hd__a21o_1 _5736_ (.A1(net24),
    .A2(_2519_),
    .B1(_2528_),
    .X(_0225_));
 sky130_fd_sc_hd__and3_1 _5737_ (.A(_2518_),
    .B(\mc.cl.next_data[7] ),
    .C(_2111_),
    .X(_2529_));
 sky130_fd_sc_hd__a21o_1 _5738_ (.A1(net25),
    .A2(_2519_),
    .B1(_2529_),
    .X(_0226_));
 sky130_fd_sc_hd__inv_2 _5739_ (.A(\cu.reg_file.reg_sp[1] ),
    .Y(_2530_));
 sky130_fd_sc_hd__mux2_1 _5740_ (.A0(_2530_),
    .A1(_1050_),
    .S(_2116_),
    .X(_2531_));
 sky130_fd_sc_hd__or4b_2 _5741_ (.A(_1007_),
    .B(_0981_),
    .C(_0989_),
    .D_N(_0994_),
    .X(_2532_));
 sky130_fd_sc_hd__or2_1 _5742_ (.A(_0296_),
    .B(_0469_),
    .X(_2533_));
 sky130_fd_sc_hd__clkbuf_2 _5743_ (.A(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__buf_2 _5744_ (.A(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__buf_2 _5745_ (.A(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__o21ai_1 _5746_ (.A1(_0986_),
    .A2(_2532_),
    .B1(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__o31a_2 _5747_ (.A1(_0740_),
    .A2(_2116_),
    .A3(_2537_),
    .B1(_2948_),
    .X(_2538_));
 sky130_fd_sc_hd__clkbuf_4 _5748_ (.A(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(\cu.reg_file.reg_sp[1] ),
    .A1(_2531_),
    .S(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__clkbuf_1 _5750_ (.A(_2540_),
    .X(_0227_));
 sky130_fd_sc_hd__nand2_1 _5751_ (.A(\cu.reg_file.reg_sp[2] ),
    .B(_2534_),
    .Y(_2541_));
 sky130_fd_sc_hd__or2_1 _5752_ (.A(\cu.reg_file.reg_sp[2] ),
    .B(_2534_),
    .X(_2542_));
 sky130_fd_sc_hd__and2_1 _5753_ (.A(_2541_),
    .B(_2542_),
    .X(_2543_));
 sky130_fd_sc_hd__xnor2_1 _5754_ (.A(_2530_),
    .B(_2543_),
    .Y(_2544_));
 sky130_fd_sc_hd__clkbuf_4 _5755_ (.A(_2115_),
    .X(_2545_));
 sky130_fd_sc_hd__mux2_1 _5756_ (.A0(_1073_),
    .A1(_2544_),
    .S(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__mux2_1 _5757_ (.A0(\cu.reg_file.reg_sp[2] ),
    .A1(_2546_),
    .S(_2539_),
    .X(_2547_));
 sky130_fd_sc_hd__clkbuf_1 _5758_ (.A(_2547_),
    .X(_0228_));
 sky130_fd_sc_hd__nor2_1 _5759_ (.A(\cu.reg_file.reg_sp[3] ),
    .B(_2534_),
    .Y(_2548_));
 sky130_fd_sc_hd__and2_1 _5760_ (.A(\cu.reg_file.reg_sp[3] ),
    .B(_2534_),
    .X(_2549_));
 sky130_fd_sc_hd__nor2_1 _5761_ (.A(_2548_),
    .B(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__a21bo_1 _5762_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_2543_),
    .B1_N(_2541_),
    .X(_2551_));
 sky130_fd_sc_hd__xor2_1 _5763_ (.A(_2550_),
    .B(_2551_),
    .X(_2552_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(_1089_),
    .A1(_2552_),
    .S(_2545_),
    .X(_2553_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(\cu.reg_file.reg_sp[3] ),
    .A1(_2553_),
    .S(_2539_),
    .X(_2554_));
 sky130_fd_sc_hd__clkbuf_1 _5766_ (.A(_2554_),
    .X(_0229_));
 sky130_fd_sc_hd__nor2_1 _5767_ (.A(\cu.reg_file.reg_sp[4] ),
    .B(_2534_),
    .Y(_2555_));
 sky130_fd_sc_hd__and2_1 _5768_ (.A(\cu.reg_file.reg_sp[4] ),
    .B(_2534_),
    .X(_2556_));
 sky130_fd_sc_hd__nor2_1 _5769_ (.A(_2555_),
    .B(_2556_),
    .Y(_2557_));
 sky130_fd_sc_hd__a21o_1 _5770_ (.A1(_2550_),
    .A2(_2551_),
    .B1(_2549_),
    .X(_2558_));
 sky130_fd_sc_hd__xor2_1 _5771_ (.A(_2557_),
    .B(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(_1160_),
    .A1(_2559_),
    .S(_2545_),
    .X(_2560_));
 sky130_fd_sc_hd__mux2_1 _5773_ (.A0(\cu.reg_file.reg_sp[4] ),
    .A1(_2560_),
    .S(_2539_),
    .X(_2561_));
 sky130_fd_sc_hd__clkbuf_1 _5774_ (.A(_2561_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_1 _5775_ (.A(\cu.reg_file.reg_sp[5] ),
    .B(_2535_),
    .X(_2562_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(\cu.reg_file.reg_sp[5] ),
    .B(_2535_),
    .Y(_2563_));
 sky130_fd_sc_hd__nand2_1 _5777_ (.A(_2562_),
    .B(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__a311o_1 _5778_ (.A1(_2550_),
    .A2(_2551_),
    .A3(_2557_),
    .B1(_2556_),
    .C1(_2549_),
    .X(_2565_));
 sky130_fd_sc_hd__xnor2_1 _5779_ (.A(_2564_),
    .B(_2565_),
    .Y(_2566_));
 sky130_fd_sc_hd__mux2_1 _5780_ (.A0(_1144_),
    .A1(_2566_),
    .S(_2545_),
    .X(_2567_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(\cu.reg_file.reg_sp[5] ),
    .A1(_2567_),
    .S(_2539_),
    .X(_2568_));
 sky130_fd_sc_hd__clkbuf_1 _5782_ (.A(_2568_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _5783_ (.A(\cu.reg_file.reg_sp[6] ),
    .B(_2535_),
    .X(_2569_));
 sky130_fd_sc_hd__nand2_1 _5784_ (.A(\cu.reg_file.reg_sp[6] ),
    .B(_2535_),
    .Y(_2570_));
 sky130_fd_sc_hd__nand2_1 _5785_ (.A(_2569_),
    .B(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__a21bo_1 _5786_ (.A1(_2562_),
    .A2(_2565_),
    .B1_N(_2563_),
    .X(_2572_));
 sky130_fd_sc_hd__xnor2_1 _5787_ (.A(_2571_),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__mux2_1 _5788_ (.A0(_1126_),
    .A1(_2573_),
    .S(_2545_),
    .X(_2574_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(\cu.reg_file.reg_sp[6] ),
    .A1(_2574_),
    .S(_2539_),
    .X(_2575_));
 sky130_fd_sc_hd__clkbuf_1 _5790_ (.A(_2575_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _5791_ (.A(\cu.reg_file.reg_sp[7] ),
    .B(_2535_),
    .X(_2576_));
 sky130_fd_sc_hd__nand2_1 _5792_ (.A(\cu.reg_file.reg_sp[7] ),
    .B(_2535_),
    .Y(_2577_));
 sky130_fd_sc_hd__nand2_1 _5793_ (.A(_2576_),
    .B(_2577_),
    .Y(_2578_));
 sky130_fd_sc_hd__a21bo_1 _5794_ (.A1(_2569_),
    .A2(_2572_),
    .B1_N(_2570_),
    .X(_2579_));
 sky130_fd_sc_hd__xnor2_1 _5795_ (.A(_2578_),
    .B(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(_1110_),
    .A1(_2580_),
    .S(_2545_),
    .X(_2581_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(\cu.reg_file.reg_sp[7] ),
    .A1(_2581_),
    .S(_2539_),
    .X(_2582_));
 sky130_fd_sc_hd__clkbuf_1 _5798_ (.A(_2582_),
    .X(_0233_));
 sky130_fd_sc_hd__or2_1 _5799_ (.A(\cu.reg_file.reg_sp[8] ),
    .B(_2535_),
    .X(_2583_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(\cu.reg_file.reg_sp[8] ),
    .B(_2535_),
    .Y(_2584_));
 sky130_fd_sc_hd__nand2_1 _5801_ (.A(_2583_),
    .B(_2584_),
    .Y(_2585_));
 sky130_fd_sc_hd__a21bo_1 _5802_ (.A1(_2576_),
    .A2(_2579_),
    .B1_N(_2577_),
    .X(_2586_));
 sky130_fd_sc_hd__xnor2_1 _5803_ (.A(_2585_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__mux2_1 _5804_ (.A0(_1622_),
    .A1(_2587_),
    .S(_2545_),
    .X(_2588_));
 sky130_fd_sc_hd__mux2_1 _5805_ (.A0(\cu.reg_file.reg_sp[8] ),
    .A1(_2588_),
    .S(_2539_),
    .X(_2589_));
 sky130_fd_sc_hd__clkbuf_1 _5806_ (.A(_2589_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _5807_ (.A(\cu.reg_file.reg_sp[9] ),
    .B(_2535_),
    .X(_2590_));
 sky130_fd_sc_hd__nand2_1 _5808_ (.A(\cu.reg_file.reg_sp[9] ),
    .B(_2536_),
    .Y(_2591_));
 sky130_fd_sc_hd__nand2_1 _5809_ (.A(_2590_),
    .B(_2591_),
    .Y(_2592_));
 sky130_fd_sc_hd__a21bo_1 _5810_ (.A1(_2583_),
    .A2(_2586_),
    .B1_N(_2584_),
    .X(_2593_));
 sky130_fd_sc_hd__xnor2_1 _5811_ (.A(_2592_),
    .B(_2593_),
    .Y(_2594_));
 sky130_fd_sc_hd__mux2_1 _5812_ (.A0(_1623_),
    .A1(_2594_),
    .S(_2545_),
    .X(_2595_));
 sky130_fd_sc_hd__mux2_1 _5813_ (.A0(\cu.reg_file.reg_sp[9] ),
    .A1(_2595_),
    .S(_2539_),
    .X(_2596_));
 sky130_fd_sc_hd__clkbuf_1 _5814_ (.A(_2596_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _5815_ (.A(\cu.reg_file.reg_sp[10] ),
    .B(_2536_),
    .X(_2597_));
 sky130_fd_sc_hd__nand2_1 _5816_ (.A(\cu.reg_file.reg_sp[10] ),
    .B(_2536_),
    .Y(_2598_));
 sky130_fd_sc_hd__nand2_1 _5817_ (.A(_2597_),
    .B(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__a21bo_1 _5818_ (.A1(_2590_),
    .A2(_2593_),
    .B1_N(_2591_),
    .X(_2600_));
 sky130_fd_sc_hd__xnor2_1 _5819_ (.A(_2599_),
    .B(_2600_),
    .Y(_2601_));
 sky130_fd_sc_hd__mux2_1 _5820_ (.A0(_1226_),
    .A1(_2601_),
    .S(_2545_),
    .X(_2602_));
 sky130_fd_sc_hd__mux2_1 _5821_ (.A0(\cu.reg_file.reg_sp[10] ),
    .A1(_2602_),
    .S(_2539_),
    .X(_2603_));
 sky130_fd_sc_hd__clkbuf_1 _5822_ (.A(_2603_),
    .X(_0236_));
 sky130_fd_sc_hd__or2_1 _5823_ (.A(\cu.reg_file.reg_sp[11] ),
    .B(_2536_),
    .X(_2604_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(\cu.reg_file.reg_sp[11] ),
    .B(_2536_),
    .Y(_2605_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_2604_),
    .B(_2605_),
    .Y(_2606_));
 sky130_fd_sc_hd__a21bo_1 _5826_ (.A1(_2597_),
    .A2(_2600_),
    .B1_N(_2598_),
    .X(_2607_));
 sky130_fd_sc_hd__xnor2_1 _5827_ (.A(_2606_),
    .B(_2607_),
    .Y(_2608_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(_1222_),
    .A1(_2608_),
    .S(_2545_),
    .X(_2609_));
 sky130_fd_sc_hd__mux2_1 _5829_ (.A0(\cu.reg_file.reg_sp[11] ),
    .A1(_2609_),
    .S(_2538_),
    .X(_2610_));
 sky130_fd_sc_hd__clkbuf_1 _5830_ (.A(_2610_),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _5831_ (.A(\cu.reg_file.reg_sp[12] ),
    .B(_2536_),
    .X(_2611_));
 sky130_fd_sc_hd__nand2_1 _5832_ (.A(\cu.reg_file.reg_sp[12] ),
    .B(_2536_),
    .Y(_2612_));
 sky130_fd_sc_hd__nand2_1 _5833_ (.A(_2611_),
    .B(_2612_),
    .Y(_2613_));
 sky130_fd_sc_hd__a21bo_1 _5834_ (.A1(_2604_),
    .A2(_2607_),
    .B1_N(_2605_),
    .X(_2614_));
 sky130_fd_sc_hd__xnor2_1 _5835_ (.A(_2613_),
    .B(_2614_),
    .Y(_2615_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(_1213_),
    .A1(_2615_),
    .S(_2115_),
    .X(_2616_));
 sky130_fd_sc_hd__mux2_1 _5837_ (.A0(\cu.reg_file.reg_sp[12] ),
    .A1(_2616_),
    .S(_2538_),
    .X(_2617_));
 sky130_fd_sc_hd__clkbuf_1 _5838_ (.A(_2617_),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _5839_ (.A(\cu.reg_file.reg_sp[13] ),
    .B(_2536_),
    .X(_2618_));
 sky130_fd_sc_hd__nand2_1 _5840_ (.A(\cu.reg_file.reg_sp[13] ),
    .B(_2536_),
    .Y(_2619_));
 sky130_fd_sc_hd__nand2_1 _5841_ (.A(_2618_),
    .B(_2619_),
    .Y(_2620_));
 sky130_fd_sc_hd__a21bo_1 _5842_ (.A1(_2611_),
    .A2(_2614_),
    .B1_N(_2612_),
    .X(_2621_));
 sky130_fd_sc_hd__xnor2_1 _5843_ (.A(_2620_),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(_1209_),
    .A1(_2622_),
    .S(_2115_),
    .X(_2623_));
 sky130_fd_sc_hd__mux2_1 _5845_ (.A0(\cu.reg_file.reg_sp[13] ),
    .A1(_2623_),
    .S(_2538_),
    .X(_2624_));
 sky130_fd_sc_hd__clkbuf_1 _5846_ (.A(_2624_),
    .X(_0239_));
 sky130_fd_sc_hd__xnor2_1 _5847_ (.A(\cu.reg_file.reg_sp[14] ),
    .B(_1287_),
    .Y(_2625_));
 sky130_fd_sc_hd__a21boi_2 _5848_ (.A1(_2618_),
    .A2(_2621_),
    .B1_N(_2619_),
    .Y(_2626_));
 sky130_fd_sc_hd__xnor2_1 _5849_ (.A(_2625_),
    .B(_2626_),
    .Y(_2627_));
 sky130_fd_sc_hd__mux2_1 _5850_ (.A0(_1624_),
    .A1(_2627_),
    .S(_2115_),
    .X(_2628_));
 sky130_fd_sc_hd__mux2_1 _5851_ (.A0(\cu.reg_file.reg_sp[14] ),
    .A1(_2628_),
    .S(_2538_),
    .X(_2629_));
 sky130_fd_sc_hd__clkbuf_1 _5852_ (.A(_2629_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _5853_ (.A(\cu.reg_file.reg_sp[14] ),
    .B(_1287_),
    .X(_2630_));
 sky130_fd_sc_hd__mux2_1 _5854_ (.A0(_1589_),
    .A1(_2630_),
    .S(_2626_),
    .X(_2631_));
 sky130_fd_sc_hd__xnor2_1 _5855_ (.A(\cu.reg_file.reg_sp[15] ),
    .B(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__mux2_1 _5856_ (.A0(_1263_),
    .A1(_2632_),
    .S(_2115_),
    .X(_2633_));
 sky130_fd_sc_hd__mux2_1 _5857_ (.A0(\cu.reg_file.reg_sp[15] ),
    .A1(_2633_),
    .S(_2538_),
    .X(_2634_));
 sky130_fd_sc_hd__clkbuf_1 _5858_ (.A(_2634_),
    .X(_0241_));
 sky130_fd_sc_hd__and2b_2 _5859_ (.A_N(_2141_),
    .B(_2320_),
    .X(_2635_));
 sky130_fd_sc_hd__o21ai_4 _5860_ (.A1(_1667_),
    .A2(_2194_),
    .B1(_2635_),
    .Y(_2636_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(_2144_),
    .A1(\ih.t.timer_max[8] ),
    .S(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_1 _5862_ (.A(_2637_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5863_ (.A0(_2155_),
    .A1(\ih.t.timer_max[9] ),
    .S(_2636_),
    .X(_2638_));
 sky130_fd_sc_hd__clkbuf_1 _5864_ (.A(_2638_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5865_ (.A0(_2157_),
    .A1(\ih.t.timer_max[10] ),
    .S(_2636_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _5866_ (.A(_2639_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5867_ (.A0(_2159_),
    .A1(\ih.t.timer_max[11] ),
    .S(_2636_),
    .X(_2640_));
 sky130_fd_sc_hd__clkbuf_1 _5868_ (.A(_2640_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5869_ (.A0(_2161_),
    .A1(\ih.t.timer_max[12] ),
    .S(_2636_),
    .X(_2641_));
 sky130_fd_sc_hd__clkbuf_1 _5870_ (.A(_2641_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5871_ (.A0(_2163_),
    .A1(\ih.t.timer_max[13] ),
    .S(_2636_),
    .X(_2642_));
 sky130_fd_sc_hd__clkbuf_1 _5872_ (.A(_2642_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5873_ (.A0(_2165_),
    .A1(\ih.t.timer_max[14] ),
    .S(_2636_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _5874_ (.A(_2643_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5875_ (.A0(_2167_),
    .A1(\ih.t.timer_max[15] ),
    .S(_2636_),
    .X(_2644_));
 sky130_fd_sc_hd__clkbuf_1 _5876_ (.A(_2644_),
    .X(_0249_));
 sky130_fd_sc_hd__o21ai_4 _5877_ (.A1(_1667_),
    .A2(_2180_),
    .B1(_2635_),
    .Y(_2645_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(_2022_),
    .A1(\ih.t.timer_max[0] ),
    .S(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__clkbuf_1 _5879_ (.A(_2646_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(_1051_),
    .A1(\ih.t.timer_max[1] ),
    .S(_2645_),
    .X(_2647_));
 sky130_fd_sc_hd__clkbuf_1 _5881_ (.A(_2647_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(_1074_),
    .A1(\ih.t.timer_max[2] ),
    .S(_2645_),
    .X(_2648_));
 sky130_fd_sc_hd__clkbuf_1 _5883_ (.A(_2648_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5884_ (.A0(_1187_),
    .A1(\ih.t.timer_max[3] ),
    .S(_2645_),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_1 _5885_ (.A(_2649_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5886_ (.A0(_1189_),
    .A1(\ih.t.timer_max[4] ),
    .S(_2645_),
    .X(_2650_));
 sky130_fd_sc_hd__clkbuf_1 _5887_ (.A(_2650_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(_1191_),
    .A1(\ih.t.timer_max[5] ),
    .S(_2645_),
    .X(_2651_));
 sky130_fd_sc_hd__clkbuf_1 _5889_ (.A(_2651_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5890_ (.A0(_1193_),
    .A1(\ih.t.timer_max[6] ),
    .S(_2645_),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _5891_ (.A(_2652_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5892_ (.A0(_1260_),
    .A1(\ih.t.timer_max[7] ),
    .S(_2645_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_1 _5893_ (.A(_2653_),
    .X(_0257_));
 sky130_fd_sc_hd__o21a_2 _5894_ (.A1(_1667_),
    .A2(_2205_),
    .B1(_2152_),
    .X(_2654_));
 sky130_fd_sc_hd__mux2_1 _5895_ (.A0(\ih.t.timer_max[16] ),
    .A1(_0618_),
    .S(_2654_),
    .X(_2655_));
 sky130_fd_sc_hd__clkbuf_1 _5896_ (.A(_2655_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5897_ (.A0(\ih.t.timer_max[17] ),
    .A1(_1051_),
    .S(_2654_),
    .X(_2656_));
 sky130_fd_sc_hd__clkbuf_1 _5898_ (.A(_2656_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5899_ (.A0(\ih.t.timer_max[18] ),
    .A1(_1074_),
    .S(_2654_),
    .X(_2657_));
 sky130_fd_sc_hd__clkbuf_1 _5900_ (.A(_2657_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5901_ (.A0(\ih.t.timer_max[19] ),
    .A1(_1187_),
    .S(_2654_),
    .X(_2658_));
 sky130_fd_sc_hd__clkbuf_1 _5902_ (.A(_2658_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5903_ (.A0(\ih.t.timer_max[20] ),
    .A1(_1189_),
    .S(_2654_),
    .X(_2659_));
 sky130_fd_sc_hd__clkbuf_1 _5904_ (.A(_2659_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5905_ (.A0(\ih.t.timer_max[21] ),
    .A1(_1191_),
    .S(_2654_),
    .X(_2660_));
 sky130_fd_sc_hd__clkbuf_1 _5906_ (.A(_2660_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5907_ (.A0(\ih.t.timer_max[22] ),
    .A1(_1193_),
    .S(_2654_),
    .X(_2661_));
 sky130_fd_sc_hd__clkbuf_1 _5908_ (.A(_2661_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5909_ (.A0(\ih.t.timer_max[23] ),
    .A1(_1260_),
    .S(_2654_),
    .X(_2662_));
 sky130_fd_sc_hd__clkbuf_1 _5910_ (.A(_2662_),
    .X(_0265_));
 sky130_fd_sc_hd__inv_2 _5911_ (.A(\cu.ir.idx[0] ),
    .Y(_2663_));
 sky130_fd_sc_hd__o21a_1 _5912_ (.A1(_2663_),
    .A2(_1644_),
    .B1(_1484_),
    .X(_2664_));
 sky130_fd_sc_hd__a21o_1 _5913_ (.A1(_2947_),
    .A2(_1482_),
    .B1(_2664_),
    .X(_2665_));
 sky130_fd_sc_hd__a22o_1 _5914_ (.A1(_2351_),
    .A2(_2664_),
    .B1(_2665_),
    .B2(net225),
    .X(_0266_));
 sky130_fd_sc_hd__nor2_4 _5915_ (.A(_2663_),
    .B(\cu.ir.idx[1] ),
    .Y(_2666_));
 sky130_fd_sc_hd__a32o_1 _5916_ (.A1(_1484_),
    .A2(_2351_),
    .A3(_2666_),
    .B1(_2665_),
    .B2(net234),
    .X(_0267_));
 sky130_fd_sc_hd__o21ai_1 _5917_ (.A1(_1780_),
    .A2(_2532_),
    .B1(net203),
    .Y(_2667_));
 sky130_fd_sc_hd__o21ai_1 _5918_ (.A1(net204),
    .A2(_2667_),
    .B1(_1781_),
    .Y(_0268_));
 sky130_fd_sc_hd__nor2_4 _5919_ (.A(\cu.ir.idx[0] ),
    .B(\cu.ir.idx[1] ),
    .Y(_2668_));
 sky130_fd_sc_hd__mux2_1 _5920_ (.A0(_2923_),
    .A1(_2350_),
    .S(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__clkbuf_1 _5921_ (.A(_2669_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5922_ (.A0(_2900_),
    .A1(_2372_),
    .S(_2668_),
    .X(_2670_));
 sky130_fd_sc_hd__clkbuf_1 _5923_ (.A(_2670_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5924_ (.A0(_2899_),
    .A1(_2391_),
    .S(_2668_),
    .X(_2671_));
 sky130_fd_sc_hd__clkbuf_1 _5925_ (.A(_2671_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(_2893_),
    .A1(_2410_),
    .S(_2668_),
    .X(_2672_));
 sky130_fd_sc_hd__clkbuf_1 _5927_ (.A(_2672_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5928_ (.A0(_0359_),
    .A1(_2429_),
    .S(_2668_),
    .X(_2673_));
 sky130_fd_sc_hd__clkbuf_1 _5929_ (.A(_2673_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5930_ (.A0(_2936_),
    .A1(_2448_),
    .S(_2668_),
    .X(_2674_));
 sky130_fd_sc_hd__clkbuf_1 _5931_ (.A(_2674_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5932_ (.A0(_2875_),
    .A1(_2467_),
    .S(_2668_),
    .X(_2675_));
 sky130_fd_sc_hd__clkbuf_1 _5933_ (.A(_2675_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5934_ (.A0(_2876_),
    .A1(_2486_),
    .S(_2668_),
    .X(_2676_));
 sky130_fd_sc_hd__clkbuf_1 _5935_ (.A(_2676_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5936_ (.A0(_0343_),
    .A1(_2350_),
    .S(_2666_),
    .X(_2677_));
 sky130_fd_sc_hd__clkbuf_1 _5937_ (.A(_2677_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5938_ (.A0(_0340_),
    .A1(_2372_),
    .S(_2666_),
    .X(_2678_));
 sky130_fd_sc_hd__clkbuf_1 _5939_ (.A(_2678_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5940_ (.A0(_0341_),
    .A1(_2391_),
    .S(_2666_),
    .X(_2679_));
 sky130_fd_sc_hd__clkbuf_1 _5941_ (.A(_2679_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5942_ (.A0(\cu.id.cb_opcode_y[0] ),
    .A1(_2410_),
    .S(_2666_),
    .X(_2680_));
 sky130_fd_sc_hd__clkbuf_1 _5943_ (.A(_2680_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(_0374_),
    .A1(_2429_),
    .S(_2666_),
    .X(_2681_));
 sky130_fd_sc_hd__clkbuf_1 _5945_ (.A(_2681_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5946_ (.A0(_0373_),
    .A1(_2448_),
    .S(_2666_),
    .X(_2682_));
 sky130_fd_sc_hd__clkbuf_1 _5947_ (.A(_2682_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5948_ (.A0(_0387_),
    .A1(_2467_),
    .S(_2666_),
    .X(_2683_));
 sky130_fd_sc_hd__clkbuf_1 _5949_ (.A(_2683_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _5950_ (.A0(_1233_),
    .A1(_2486_),
    .S(_2666_),
    .X(_2684_));
 sky130_fd_sc_hd__clkbuf_1 _5951_ (.A(_2684_),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _5952_ (.A(_2663_),
    .B(\cu.ir.idx[1] ),
    .X(_2685_));
 sky130_fd_sc_hd__clkbuf_4 _5953_ (.A(_2685_),
    .X(_2686_));
 sky130_fd_sc_hd__mux2_1 _5954_ (.A0(\cu.id.imm_i[8] ),
    .A1(_2350_),
    .S(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__clkbuf_1 _5955_ (.A(_2687_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _5956_ (.A0(\cu.id.imm_i[9] ),
    .A1(_2372_),
    .S(_2686_),
    .X(_2688_));
 sky130_fd_sc_hd__clkbuf_1 _5957_ (.A(_2688_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _5958_ (.A0(\cu.id.imm_i[10] ),
    .A1(_2391_),
    .S(_2686_),
    .X(_2689_));
 sky130_fd_sc_hd__clkbuf_1 _5959_ (.A(_2689_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _5960_ (.A0(\cu.id.imm_i[11] ),
    .A1(_2410_),
    .S(_2686_),
    .X(_2690_));
 sky130_fd_sc_hd__clkbuf_1 _5961_ (.A(_2690_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _5962_ (.A0(\cu.id.imm_i[12] ),
    .A1(_2429_),
    .S(_2686_),
    .X(_2691_));
 sky130_fd_sc_hd__clkbuf_1 _5963_ (.A(_2691_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _5964_ (.A0(\cu.id.imm_i[13] ),
    .A1(_2448_),
    .S(_2686_),
    .X(_2692_));
 sky130_fd_sc_hd__clkbuf_1 _5965_ (.A(_2692_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _5966_ (.A0(\cu.id.imm_i[14] ),
    .A1(_2467_),
    .S(_2686_),
    .X(_2693_));
 sky130_fd_sc_hd__clkbuf_1 _5967_ (.A(_2693_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _5968_ (.A0(\cu.id.imm_i[15] ),
    .A1(_2486_),
    .S(_2686_),
    .X(_2694_));
 sky130_fd_sc_hd__clkbuf_1 _5969_ (.A(_2694_),
    .X(_0292_));
 sky130_fd_sc_hd__dfrtp_4 _5970_ (.CLK(clknet_leaf_36_clk),
    .D(_0007_),
    .RESET_B(net160),
    .Q(\alu.Cin ));
 sky130_fd_sc_hd__dfrtp_1 _5971_ (.CLK(clknet_leaf_36_clk),
    .D(_0008_),
    .RESET_B(net160),
    .Q(\cu.alu_f[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5972_ (.CLK(clknet_leaf_36_clk),
    .D(_0009_),
    .RESET_B(net161),
    .Q(\cu.alu_f[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5973_ (.CLK(clknet_leaf_33_clk),
    .D(_0010_),
    .RESET_B(net164),
    .Q(\cu.alu_f[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5974_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0011_),
    .RESET_B(net161),
    .Q(\cu.alu_f[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5975_ (.CLK(clknet_leaf_33_clk),
    .D(_0012_),
    .RESET_B(net163),
    .Q(\cu.alu_f[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5976_ (.CLK(clknet_leaf_36_clk),
    .D(_0013_),
    .RESET_B(net161),
    .Q(\cu.alu_f[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5977_ (.CLK(clknet_leaf_33_clk),
    .D(_0014_),
    .RESET_B(net163),
    .Q(\cu.alu_f[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5978_ (.CLK(clknet_leaf_30_clk),
    .D(_0016_),
    .RESET_B(net188),
    .Q(\cu.pc.pc_o[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5979_ (.CLK(clknet_leaf_30_clk),
    .D(_0017_),
    .RESET_B(net187),
    .Q(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5980_ (.CLK(clknet_leaf_30_clk),
    .D(_0018_),
    .RESET_B(net187),
    .Q(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5981_ (.CLK(clknet_leaf_28_clk),
    .D(_0019_),
    .RESET_B(net187),
    .Q(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5982_ (.CLK(clknet_leaf_28_clk),
    .D(_0020_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__dfrtp_4 _5983_ (.CLK(clknet_leaf_28_clk),
    .D(_0021_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__dfrtp_4 _5984_ (.CLK(clknet_leaf_29_clk),
    .D(_0022_),
    .RESET_B(net188),
    .Q(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _5985_ (.CLK(clknet_leaf_28_clk),
    .D(_0023_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _5986_ (.CLK(clknet_leaf_28_clk),
    .D(_0024_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _5987_ (.CLK(clknet_leaf_28_clk),
    .D(_0025_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5988_ (.CLK(clknet_leaf_29_clk),
    .D(_0026_),
    .RESET_B(net188),
    .Q(\cu.pc.pc_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _5989_ (.CLK(clknet_leaf_29_clk),
    .D(_0027_),
    .RESET_B(net188),
    .Q(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__dfstp_2 _5990_ (.CLK(clknet_leaf_34_clk),
    .D(_0028_),
    .SET_B(net163),
    .Q(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _5991_ (.CLK(clknet_leaf_34_clk),
    .D(_0029_),
    .RESET_B(net163),
    .Q(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _5992_ (.CLK(clknet_leaf_34_clk),
    .D(_0030_),
    .RESET_B(net163),
    .Q(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__dfrtp_4 _5993_ (.CLK(clknet_leaf_29_clk),
    .D(_0031_),
    .RESET_B(net188),
    .Q(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _5994_ (.CLK(clknet_leaf_2_clk),
    .D(_0032_),
    .RESET_B(net155),
    .Q(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5995_ (.CLK(clknet_leaf_2_clk),
    .D(_0033_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5996_ (.CLK(clknet_leaf_2_clk),
    .D(_0034_),
    .RESET_B(net155),
    .Q(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5997_ (.CLK(clknet_leaf_2_clk),
    .D(_0035_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5998_ (.CLK(clknet_leaf_2_clk),
    .D(_0036_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_a[4] ));
 sky130_fd_sc_hd__dfrtp_4 _5999_ (.CLK(clknet_leaf_2_clk),
    .D(_0037_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_a[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6000_ (.CLK(clknet_leaf_4_clk),
    .D(_0038_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_a[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6001_ (.CLK(clknet_leaf_3_clk),
    .D(_0039_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6002_ (.CLK(clknet_leaf_20_clk),
    .D(_0040_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6003_ (.CLK(clknet_leaf_5_clk),
    .D(_0041_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6004_ (.CLK(clknet_leaf_20_clk),
    .D(_0042_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6005_ (.CLK(clknet_leaf_31_clk),
    .D(_0043_),
    .RESET_B(net183),
    .Q(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6006_ (.CLK(clknet_leaf_31_clk),
    .D(_0044_),
    .RESET_B(net183),
    .Q(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6007_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0045_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6008_ (.CLK(clknet_leaf_5_clk),
    .D(_0046_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6009_ (.CLK(clknet_leaf_31_clk),
    .D(_0047_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6010_ (.CLK(clknet_leaf_7_clk),
    .D(_0048_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6011_ (.CLK(clknet_leaf_5_clk),
    .D(_0049_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6012_ (.CLK(clknet_leaf_6_clk),
    .D(_0050_),
    .RESET_B(net171),
    .Q(\cu.reg_file.reg_c[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6013_ (.CLK(clknet_leaf_6_clk),
    .D(_0051_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_c[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6014_ (.CLK(clknet_leaf_6_clk),
    .D(_0052_),
    .RESET_B(net171),
    .Q(\cu.reg_file.reg_c[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6015_ (.CLK(clknet_leaf_7_clk),
    .D(_0053_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_c[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6016_ (.CLK(clknet_leaf_7_clk),
    .D(_0054_),
    .RESET_B(net171),
    .Q(\cu.reg_file.reg_c[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6017_ (.CLK(clknet_leaf_7_clk),
    .D(_0055_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6018_ (.CLK(clknet_leaf_31_clk),
    .D(_0056_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6019_ (.CLK(clknet_leaf_6_clk),
    .D(_0057_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6020_ (.CLK(clknet_leaf_20_clk),
    .D(_0058_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6021_ (.CLK(clknet_leaf_31_clk),
    .D(_0059_),
    .RESET_B(net183),
    .Q(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6022_ (.CLK(clknet_leaf_31_clk),
    .D(_0060_),
    .RESET_B(net183),
    .Q(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6023_ (.CLK(clknet_leaf_31_clk),
    .D(_0061_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6024_ (.CLK(clknet_leaf_5_clk),
    .D(_0062_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6025_ (.CLK(clknet_leaf_31_clk),
    .D(_0063_),
    .RESET_B(net185),
    .Q(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6026_ (.CLK(clknet_leaf_9_clk),
    .D(_0064_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_e[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6027_ (.CLK(clknet_leaf_2_clk),
    .D(_0065_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6028_ (.CLK(clknet_leaf_2_clk),
    .D(_0066_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6029_ (.CLK(clknet_leaf_2_clk),
    .D(_0067_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6030_ (.CLK(clknet_leaf_5_clk),
    .D(_0068_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_e[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6031_ (.CLK(clknet_leaf_2_clk),
    .D(_0069_),
    .RESET_B(net155),
    .Q(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6032_ (.CLK(clknet_leaf_4_clk),
    .D(_0070_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_e[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6033_ (.CLK(clknet_leaf_4_clk),
    .D(_0071_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_e[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6034_ (.CLK(clknet_leaf_33_clk),
    .D(_0072_),
    .RESET_B(net163),
    .Q(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6035_ (.CLK(clknet_leaf_34_clk),
    .D(_0073_),
    .RESET_B(net163),
    .Q(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6036_ (.CLK(clknet_leaf_33_clk),
    .D(_0074_),
    .RESET_B(net163),
    .Q(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6037_ (.CLK(clknet_leaf_33_clk),
    .D(_0075_),
    .RESET_B(net163),
    .Q(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6038_ (.CLK(clknet_leaf_33_clk),
    .D(_0076_),
    .RESET_B(net164),
    .Q(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6039_ (.CLK(clknet_leaf_33_clk),
    .D(_0077_),
    .RESET_B(net163),
    .Q(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6040_ (.CLK(clknet_leaf_33_clk),
    .D(_0078_),
    .RESET_B(net164),
    .Q(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6041_ (.CLK(clknet_leaf_34_clk),
    .D(_0079_),
    .RESET_B(net164),
    .Q(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6042_ (.CLK(clknet_leaf_40_clk),
    .D(_0080_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6043_ (.CLK(clknet_leaf_4_clk),
    .D(_0081_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6044_ (.CLK(clknet_leaf_5_clk),
    .D(_0082_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_l[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6045_ (.CLK(clknet_leaf_6_clk),
    .D(_0083_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_l[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6046_ (.CLK(clknet_leaf_6_clk),
    .D(_0084_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_l[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6047_ (.CLK(clknet_leaf_7_clk),
    .D(_0085_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_l[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6048_ (.CLK(clknet_leaf_6_clk),
    .D(_0086_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_l[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6049_ (.CLK(clknet_leaf_6_clk),
    .D(_0087_),
    .RESET_B(net170),
    .Q(\cu.reg_file.reg_l[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6050_ (.CLK(clknet_leaf_22_clk),
    .D(_0088_),
    .RESET_B(net190),
    .Q(\mc.cl.next_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6051_ (.CLK(clknet_leaf_22_clk),
    .D(_0089_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6052_ (.CLK(clknet_leaf_22_clk),
    .D(_0090_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6053_ (.CLK(clknet_leaf_22_clk),
    .D(_0091_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6054_ (.CLK(clknet_leaf_22_clk),
    .D(_0092_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6055_ (.CLK(clknet_leaf_24_clk),
    .D(_0093_),
    .RESET_B(net191),
    .Q(\mc.cl.next_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6056_ (.CLK(clknet_leaf_22_clk),
    .D(_0094_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6057_ (.CLK(clknet_leaf_22_clk),
    .D(_0095_),
    .RESET_B(net190),
    .Q(\mc.cl.next_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6058_ (.CLK(clknet_leaf_25_clk),
    .D(\mc.cc.enable ),
    .RESET_B(net194),
    .Q(\mc.cc.enable_edge_detector.prev_data ));
 sky130_fd_sc_hd__dfrtp_4 _6059_ (.CLK(clknet_leaf_4_clk),
    .D(_0096_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_sp[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6060_ (.CLK(clknet_leaf_25_clk),
    .D(\mc.rw.next_state[0] ),
    .RESET_B(net194),
    .Q(\mc.rw.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6061_ (.CLK(clknet_leaf_25_clk),
    .D(\mc.rw.next_state[1] ),
    .RESET_B(net194),
    .Q(\mc.rw.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6062_ (.CLK(clknet_leaf_25_clk),
    .D(\mc.rw.next_state[2] ),
    .RESET_B(net194),
    .Q(\mc.rw.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6063_ (.CLK(clknet_leaf_25_clk),
    .D(net211),
    .RESET_B(net194),
    .Q(\mc.cc.count[0] ));
 sky130_fd_sc_hd__dfstp_1 _6064_ (.CLK(clknet_leaf_26_clk),
    .D(_0098_),
    .SET_B(net194),
    .Q(\mc.cc.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6065_ (.CLK(clknet_leaf_26_clk),
    .D(net224),
    .RESET_B(net194),
    .Q(\mc.cc.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6066_ (.CLK(clknet_leaf_26_clk),
    .D(_0100_),
    .RESET_B(net195),
    .Q(\mc.cc.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6067_ (.CLK(clknet_leaf_19_clk),
    .D(_0101_),
    .RESET_B(net180),
    .Q(\ih.gpio_interrupt_mask[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6068_ (.CLK(clknet_leaf_16_clk),
    .D(_0102_),
    .RESET_B(net174),
    .Q(\ih.gpio_interrupt_mask[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6069_ (.CLK(clknet_leaf_12_clk),
    .D(_0103_),
    .RESET_B(net174),
    .Q(\ih.gpio_interrupt_mask[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6070_ (.CLK(clknet_leaf_12_clk),
    .D(_0104_),
    .RESET_B(net168),
    .Q(\ih.gpio_interrupt_mask[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6071_ (.CLK(clknet_leaf_12_clk),
    .D(_0105_),
    .RESET_B(net174),
    .Q(\ih.gpio_interrupt_mask[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6072_ (.CLK(clknet_leaf_16_clk),
    .D(_0106_),
    .RESET_B(net174),
    .Q(\ih.gpio_interrupt_mask[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6073_ (.CLK(clknet_leaf_19_clk),
    .D(_0107_),
    .RESET_B(net180),
    .Q(\ih.gpio_interrupt_mask[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6074_ (.CLK(clknet_leaf_16_clk),
    .D(_0108_),
    .RESET_B(net180),
    .Q(\ih.gpio_interrupt_mask[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6075_ (.CLK(clknet_leaf_18_clk),
    .D(_0109_),
    .RESET_B(net180),
    .Q(\ih.t.enable ));
 sky130_fd_sc_hd__dfrtp_2 _6076_ (.CLK(clknet_leaf_23_clk),
    .D(_0110_),
    .RESET_B(net191),
    .Q(\ih.t.timer_max[24] ));
 sky130_fd_sc_hd__dfrtp_4 _6077_ (.CLK(clknet_leaf_23_clk),
    .D(_0111_),
    .RESET_B(net191),
    .Q(\ih.t.timer_max[25] ));
 sky130_fd_sc_hd__dfrtp_2 _6078_ (.CLK(clknet_leaf_23_clk),
    .D(_0112_),
    .RESET_B(net191),
    .Q(\ih.t.timer_max[26] ));
 sky130_fd_sc_hd__dfrtp_2 _6079_ (.CLK(clknet_leaf_23_clk),
    .D(_0113_),
    .RESET_B(net192),
    .Q(\ih.t.timer_max[27] ));
 sky130_fd_sc_hd__dfrtp_4 _6080_ (.CLK(clknet_leaf_23_clk),
    .D(_0114_),
    .RESET_B(net192),
    .Q(\ih.t.timer_max[28] ));
 sky130_fd_sc_hd__dfrtp_2 _6081_ (.CLK(clknet_leaf_23_clk),
    .D(_0115_),
    .RESET_B(net193),
    .Q(\ih.t.timer_max[29] ));
 sky130_fd_sc_hd__dfrtp_2 _6082_ (.CLK(clknet_leaf_23_clk),
    .D(_0116_),
    .RESET_B(net191),
    .Q(\ih.t.timer_max[30] ));
 sky130_fd_sc_hd__dfrtp_2 _6083_ (.CLK(clknet_leaf_23_clk),
    .D(_0117_),
    .RESET_B(net191),
    .Q(\ih.t.timer_max[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6084_ (.CLK(clknet_leaf_19_clk),
    .D(_0118_),
    .RESET_B(net180),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _6085_ (.CLK(clknet_leaf_12_clk),
    .D(_0119_),
    .RESET_B(net174),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _6086_ (.CLK(clknet_leaf_13_clk),
    .D(_0120_),
    .RESET_B(net173),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_4 _6087_ (.CLK(clknet_leaf_8_clk),
    .D(_0121_),
    .RESET_B(net168),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_4 _6088_ (.CLK(clknet_leaf_24_clk),
    .D(_0122_),
    .RESET_B(net190),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_4 _6089_ (.CLK(clknet_leaf_12_clk),
    .D(_0123_),
    .RESET_B(net168),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_4 _6090_ (.CLK(clknet_leaf_7_clk),
    .D(_0124_),
    .RESET_B(net171),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_4 _6091_ (.CLK(clknet_leaf_21_clk),
    .D(_0125_),
    .RESET_B(net183),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _6092_ (.CLK(clknet_leaf_24_clk),
    .D(_0126_),
    .RESET_B(net192),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _6093_ (.CLK(clknet_leaf_13_clk),
    .D(_0127_),
    .RESET_B(net173),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_4 _6094_ (.CLK(clknet_leaf_28_clk),
    .D(_0128_),
    .RESET_B(net186),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _6095_ (.CLK(clknet_leaf_10_clk),
    .D(_0129_),
    .RESET_B(net166),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_4 _6096_ (.CLK(clknet_leaf_10_clk),
    .D(_0130_),
    .RESET_B(net166),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_2 _6097_ (.CLK(clknet_leaf_27_clk),
    .D(_0131_),
    .RESET_B(net195),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_4 _6098_ (.CLK(clknet_leaf_9_clk),
    .D(_0132_),
    .RESET_B(net165),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_2 _6099_ (.CLK(clknet_leaf_9_clk),
    .D(_0133_),
    .RESET_B(net165),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_4 _6100_ (.CLK(clknet_leaf_21_clk),
    .D(_0134_),
    .RESET_B(net182),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_4 _6101_ (.CLK(clknet_leaf_28_clk),
    .D(_0135_),
    .RESET_B(net186),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_2 _6102_ (.CLK(clknet_leaf_13_clk),
    .D(_0136_),
    .RESET_B(net173),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_4 _6103_ (.CLK(clknet_leaf_31_clk),
    .D(_0137_),
    .RESET_B(net183),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_2 _6104_ (.CLK(clknet_leaf_9_clk),
    .D(_0138_),
    .RESET_B(net166),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_4 _6105_ (.CLK(clknet_leaf_9_clk),
    .D(_0139_),
    .RESET_B(net165),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_4 _6106_ (.CLK(clknet_leaf_28_clk),
    .D(_0140_),
    .RESET_B(net186),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_2 _6107_ (.CLK(clknet_leaf_27_clk),
    .D(_0141_),
    .RESET_B(net195),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_4 _6108_ (.CLK(clknet_leaf_28_clk),
    .D(_0142_),
    .RESET_B(net195),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _6109_ (.CLK(clknet_leaf_28_clk),
    .D(_0143_),
    .RESET_B(net186),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _6110_ (.CLK(clknet_leaf_11_clk),
    .D(_0144_),
    .RESET_B(net167),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _6111_ (.CLK(clknet_leaf_31_clk),
    .D(_0145_),
    .RESET_B(net183),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _6112_ (.CLK(clknet_leaf_13_clk),
    .D(_0146_),
    .RESET_B(net173),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_2 _6113_ (.CLK(clknet_leaf_28_clk),
    .D(_0147_),
    .RESET_B(net186),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_4 _6114_ (.CLK(clknet_leaf_27_clk),
    .D(_0148_),
    .RESET_B(net195),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 _6115_ (.CLK(clknet_leaf_28_clk),
    .D(_0149_),
    .RESET_B(net187),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 _6116_ (.CLK(clknet_leaf_24_clk),
    .D(_0150_),
    .RESET_B(net192),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _6117_ (.CLK(clknet_leaf_13_clk),
    .D(_0151_),
    .RESET_B(net173),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_4 _6118_ (.CLK(clknet_leaf_11_clk),
    .D(_0152_),
    .RESET_B(net167),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_2 _6119_ (.CLK(clknet_leaf_10_clk),
    .D(_0153_),
    .RESET_B(net167),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_4 _6120_ (.CLK(clknet_leaf_13_clk),
    .D(_0154_),
    .RESET_B(net173),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_4 _6121_ (.CLK(clknet_leaf_21_clk),
    .D(_0155_),
    .RESET_B(net184),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_4 _6122_ (.CLK(clknet_leaf_11_clk),
    .D(_0156_),
    .RESET_B(net167),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_1 _6123_ (.CLK(clknet_leaf_16_clk),
    .D(_0157_),
    .RESET_B(net174),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_1 _6124_ (.CLK(clknet_leaf_23_clk),
    .D(_0158_),
    .RESET_B(net192),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _6125_ (.CLK(clknet_leaf_13_clk),
    .D(_0159_),
    .RESET_B(net173),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_4 _6126_ (.CLK(clknet_leaf_11_clk),
    .D(_0160_),
    .RESET_B(net167),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 _6127_ (.CLK(clknet_leaf_10_clk),
    .D(_0161_),
    .RESET_B(net167),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_4 _6128_ (.CLK(clknet_leaf_22_clk),
    .D(_0162_),
    .RESET_B(net190),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 _6129_ (.CLK(clknet_leaf_21_clk),
    .D(_0163_),
    .RESET_B(net182),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_4 _6130_ (.CLK(clknet_leaf_20_clk),
    .D(_0164_),
    .RESET_B(net172),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_4 _6131_ (.CLK(clknet_leaf_24_clk),
    .D(_0165_),
    .RESET_B(net192),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 _6132_ (.CLK(clknet_leaf_27_clk),
    .D(_0166_),
    .RESET_B(net195),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_1 _6133_ (.CLK(clknet_leaf_13_clk),
    .D(_0167_),
    .RESET_B(net173),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_2 _6134_ (.CLK(clknet_leaf_10_clk),
    .D(_0168_),
    .RESET_B(net166),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_4 _6135_ (.CLK(clknet_leaf_9_clk),
    .D(_0169_),
    .RESET_B(net165),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_4 _6136_ (.CLK(clknet_leaf_9_clk),
    .D(_0170_),
    .RESET_B(net165),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_2 _6137_ (.CLK(clknet_leaf_10_clk),
    .D(_0171_),
    .RESET_B(net166),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_4 _6138_ (.CLK(clknet_leaf_28_clk),
    .D(_0172_),
    .RESET_B(net187),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_4 _6139_ (.CLK(clknet_leaf_20_clk),
    .D(_0173_),
    .RESET_B(net182),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_2 _6140_ (.CLK(clknet_leaf_24_clk),
    .D(_0174_),
    .RESET_B(net192),
    .Q(net132));
 sky130_fd_sc_hd__dfrtp_4 _6141_ (.CLK(clknet_leaf_24_clk),
    .D(_0175_),
    .RESET_B(net192),
    .Q(net133));
 sky130_fd_sc_hd__dfrtp_1 _6142_ (.CLK(clknet_leaf_13_clk),
    .D(_0176_),
    .RESET_B(net173),
    .Q(net134));
 sky130_fd_sc_hd__dfrtp_1 _6143_ (.CLK(clknet_leaf_12_clk),
    .D(_0177_),
    .RESET_B(net168),
    .Q(net135));
 sky130_fd_sc_hd__dfrtp_4 _6144_ (.CLK(clknet_leaf_9_clk),
    .D(_0178_),
    .RESET_B(net165),
    .Q(net136));
 sky130_fd_sc_hd__dfrtp_2 _6145_ (.CLK(clknet_leaf_10_clk),
    .D(_0179_),
    .RESET_B(net166),
    .Q(net137));
 sky130_fd_sc_hd__dfrtp_2 _6146_ (.CLK(clknet_leaf_11_clk),
    .D(_0180_),
    .RESET_B(net167),
    .Q(net138));
 sky130_fd_sc_hd__dfrtp_4 _6147_ (.CLK(clknet_leaf_31_clk),
    .D(_0181_),
    .RESET_B(net183),
    .Q(net139));
 sky130_fd_sc_hd__dfrtp_4 _6148_ (.CLK(clknet_leaf_20_clk),
    .D(_0182_),
    .RESET_B(net182),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_4 _6149_ (.CLK(clknet_leaf_8_clk),
    .D(_0183_),
    .RESET_B(net172),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_4 _6150_ (.CLK(clknet_leaf_12_clk),
    .D(_0184_),
    .RESET_B(net174),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_4 _6151_ (.CLK(clknet_leaf_11_clk),
    .D(_0185_),
    .RESET_B(net168),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_4 _6152_ (.CLK(clknet_leaf_12_clk),
    .D(_0186_),
    .RESET_B(net177),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_4 _6153_ (.CLK(clknet_leaf_15_clk),
    .D(_0187_),
    .RESET_B(net177),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_4 _6154_ (.CLK(clknet_leaf_13_clk),
    .D(_0188_),
    .RESET_B(net173),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_2 _6155_ (.CLK(clknet_leaf_11_clk),
    .D(_0189_),
    .RESET_B(net168),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _6156_ (.CLK(clknet_leaf_19_clk),
    .D(_0190_),
    .RESET_B(net180),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_4 _6157_ (.CLK(clknet_leaf_20_clk),
    .D(_0191_),
    .RESET_B(net172),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_4 _6158_ (.CLK(clknet_leaf_20_clk),
    .D(_0192_),
    .RESET_B(net172),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_4 _6159_ (.CLK(clknet_leaf_20_clk),
    .D(_0193_),
    .RESET_B(net172),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_4 _6160_ (.CLK(clknet_leaf_20_clk),
    .D(_0194_),
    .RESET_B(net172),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _6161_ (.CLK(clknet_leaf_10_clk),
    .D(_0195_),
    .RESET_B(net167),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_4 _6162_ (.CLK(clknet_leaf_10_clk),
    .D(_0196_),
    .RESET_B(net166),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_2 _6163_ (.CLK(clknet_leaf_10_clk),
    .D(_0197_),
    .RESET_B(net166),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _6164_ (.CLK(clknet_leaf_41_clk),
    .D(_0198_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_mem[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6165_ (.CLK(clknet_leaf_0_clk),
    .D(_0199_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_mem[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6166_ (.CLK(clknet_leaf_3_clk),
    .D(_0200_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_mem[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6167_ (.CLK(clknet_leaf_3_clk),
    .D(_0201_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6168_ (.CLK(clknet_leaf_3_clk),
    .D(_0202_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6169_ (.CLK(clknet_leaf_3_clk),
    .D(_0203_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_mem[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6170_ (.CLK(clknet_leaf_40_clk),
    .D(_0204_),
    .RESET_B(net164),
    .Q(\cu.reg_file.reg_mem[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6171_ (.CLK(clknet_leaf_38_clk),
    .D(_0205_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_mem[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6172_ (.CLK(clknet_leaf_21_clk),
    .D(_0206_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[8] ));
 sky130_fd_sc_hd__dfrtp_2 _6173_ (.CLK(clknet_leaf_21_clk),
    .D(_0207_),
    .RESET_B(net184),
    .Q(\cu.reg_file.reg_mem[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6174_ (.CLK(clknet_leaf_21_clk),
    .D(_0208_),
    .RESET_B(net184),
    .Q(\cu.reg_file.reg_mem[10] ));
 sky130_fd_sc_hd__dfrtp_2 _6175_ (.CLK(clknet_leaf_20_clk),
    .D(_0209_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__dfrtp_2 _6176_ (.CLK(clknet_leaf_21_clk),
    .D(_0210_),
    .RESET_B(net184),
    .Q(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6177_ (.CLK(clknet_leaf_21_clk),
    .D(_0211_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6178_ (.CLK(clknet_leaf_21_clk),
    .D(_0212_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[14] ));
 sky130_fd_sc_hd__dfrtp_4 _6179_ (.CLK(clknet_leaf_21_clk),
    .D(_0213_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6180_ (.CLK(clknet_leaf_36_clk),
    .D(_0000_),
    .RESET_B(net161),
    .Q(\ih.interrupt_source[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6181_ (.CLK(clknet_leaf_25_clk),
    .D(_0214_),
    .Q(\mc.cl.cmp_o ));
 sky130_fd_sc_hd__dfrtp_1 _6182_ (.CLK(clknet_leaf_7_clk),
    .D(_0215_),
    .RESET_B(net172),
    .Q(\ih.input_handler_enable ));
 sky130_fd_sc_hd__dfrtp_4 _6183_ (.CLK(clknet_leaf_22_clk),
    .D(_0216_),
    .RESET_B(net190),
    .Q(\mc.count ));
 sky130_fd_sc_hd__dfrtp_1 _6184_ (.CLK(clknet_leaf_35_clk),
    .D(net199),
    .RESET_B(net162),
    .Q(\ih.interrupt_source[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6185_ (.CLK(clknet_leaf_35_clk),
    .D(_0218_),
    .RESET_B(net162),
    .Q(\ih.interrupt_source[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6186_ (.CLK(clknet_leaf_22_clk),
    .D(_0219_),
    .RESET_B(net190),
    .Q(\mc.cl.next_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6187_ (.CLK(clknet_leaf_22_clk),
    .D(_0220_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6188_ (.CLK(clknet_leaf_22_clk),
    .D(_0221_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6189_ (.CLK(clknet_leaf_22_clk),
    .D(_0222_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6190_ (.CLK(clknet_leaf_22_clk),
    .D(_0223_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6191_ (.CLK(clknet_leaf_22_clk),
    .D(_0224_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6192_ (.CLK(clknet_leaf_22_clk),
    .D(_0225_),
    .RESET_B(net190),
    .Q(\mc.cl.next_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6193_ (.CLK(clknet_leaf_22_clk),
    .D(_0226_),
    .RESET_B(net196),
    .Q(\mc.cl.next_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6194_ (.CLK(clknet_leaf_35_clk),
    .D(net1),
    .RESET_B(net162),
    .Q(\ih.ip_ed.prev_data ));
 sky130_fd_sc_hd__dfrtp_1 _6195_ (.CLK(clknet_leaf_7_clk),
    .D(net2),
    .RESET_B(net171),
    .Q(\ih.ih.ih.prev_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6196_ (.CLK(clknet_leaf_10_clk),
    .D(net9),
    .RESET_B(net167),
    .Q(\ih.ih.ih.prev_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6197_ (.CLK(clknet_leaf_11_clk),
    .D(net10),
    .RESET_B(net168),
    .Q(\ih.ih.ih.prev_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6198_ (.CLK(clknet_leaf_11_clk),
    .D(net11),
    .RESET_B(net168),
    .Q(\ih.ih.ih.prev_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6199_ (.CLK(clknet_leaf_11_clk),
    .D(net12),
    .RESET_B(net168),
    .Q(\ih.ih.ih.prev_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6200_ (.CLK(clknet_leaf_9_clk),
    .D(net13),
    .RESET_B(net169),
    .Q(\ih.ih.ih.prev_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6201_ (.CLK(clknet_leaf_12_clk),
    .D(net14),
    .RESET_B(net169),
    .Q(\ih.ih.ih.prev_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6202_ (.CLK(clknet_leaf_7_clk),
    .D(net15),
    .RESET_B(net172),
    .Q(\ih.ih.ih.prev_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6203_ (.CLK(clknet_leaf_7_clk),
    .D(net16),
    .RESET_B(net172),
    .Q(\ih.ih.ih.prev_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6204_ (.CLK(clknet_leaf_8_clk),
    .D(net17),
    .RESET_B(net169),
    .Q(\ih.ih.ih.prev_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6205_ (.CLK(clknet_leaf_9_clk),
    .D(net3),
    .RESET_B(net169),
    .Q(\ih.ih.ih.prev_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6206_ (.CLK(clknet_leaf_10_clk),
    .D(net4),
    .RESET_B(net167),
    .Q(\ih.ih.ih.prev_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6207_ (.CLK(clknet_leaf_12_clk),
    .D(net5),
    .RESET_B(net169),
    .Q(\ih.ih.ih.prev_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6208_ (.CLK(clknet_leaf_8_clk),
    .D(net6),
    .RESET_B(net169),
    .Q(\ih.ih.ih.prev_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6209_ (.CLK(clknet_leaf_9_clk),
    .D(net7),
    .RESET_B(net169),
    .Q(\ih.ih.ih.prev_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6210_ (.CLK(clknet_leaf_9_clk),
    .D(net8),
    .RESET_B(net166),
    .Q(\ih.ih.ih.prev_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6211_ (.CLK(clknet_leaf_7_clk),
    .D(\ih.ih.int_f.data_in ),
    .RESET_B(net181),
    .Q(\ih.ih.int_f.prev_data ));
 sky130_fd_sc_hd__dfrtp_4 _6212_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[0] ),
    .RESET_B(net176),
    .Q(\ih.t.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6213_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[1] ),
    .RESET_B(net176),
    .Q(\ih.t.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6214_ (.CLK(clknet_leaf_13_clk),
    .D(\ih.t.next_count[2] ),
    .RESET_B(net176),
    .Q(\ih.t.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6215_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[3] ),
    .RESET_B(net176),
    .Q(\ih.t.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6216_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[4] ),
    .RESET_B(net176),
    .Q(\ih.t.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6217_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[5] ),
    .RESET_B(net176),
    .Q(\ih.t.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6218_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[6] ),
    .RESET_B(net176),
    .Q(\ih.t.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6219_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[7] ),
    .RESET_B(net176),
    .Q(\ih.t.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6220_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[8] ),
    .RESET_B(net176),
    .Q(\ih.t.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6221_ (.CLK(clknet_leaf_14_clk),
    .D(\ih.t.next_count[9] ),
    .RESET_B(net175),
    .Q(\ih.t.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6222_ (.CLK(clknet_leaf_15_clk),
    .D(net216),
    .RESET_B(net175),
    .Q(\ih.t.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6223_ (.CLK(clknet_leaf_15_clk),
    .D(\ih.t.next_count[11] ),
    .RESET_B(net175),
    .Q(\ih.t.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6224_ (.CLK(clknet_leaf_15_clk),
    .D(\ih.t.next_count[12] ),
    .RESET_B(net175),
    .Q(\ih.t.count[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6225_ (.CLK(clknet_leaf_15_clk),
    .D(\ih.t.next_count[13] ),
    .RESET_B(net175),
    .Q(\ih.t.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6226_ (.CLK(clknet_leaf_15_clk),
    .D(\ih.t.next_count[14] ),
    .RESET_B(net177),
    .Q(\ih.t.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6227_ (.CLK(clknet_leaf_17_clk),
    .D(\ih.t.next_count[15] ),
    .RESET_B(net178),
    .Q(\ih.t.count[15] ));
 sky130_fd_sc_hd__dfrtp_2 _6228_ (.CLK(clknet_leaf_17_clk),
    .D(\ih.t.next_count[16] ),
    .RESET_B(net178),
    .Q(\ih.t.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _6229_ (.CLK(clknet_leaf_17_clk),
    .D(\ih.t.next_count[17] ),
    .RESET_B(net178),
    .Q(\ih.t.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6230_ (.CLK(clknet_leaf_17_clk),
    .D(\ih.t.next_count[18] ),
    .RESET_B(net178),
    .Q(\ih.t.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6231_ (.CLK(clknet_leaf_17_clk),
    .D(net214),
    .RESET_B(net179),
    .Q(\ih.t.count[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6232_ (.CLK(clknet_leaf_17_clk),
    .D(\ih.t.next_count[20] ),
    .RESET_B(net179),
    .Q(\ih.t.count[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6233_ (.CLK(clknet_leaf_17_clk),
    .D(\ih.t.next_count[21] ),
    .RESET_B(net179),
    .Q(\ih.t.count[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6234_ (.CLK(clknet_leaf_17_clk),
    .D(\ih.t.next_count[22] ),
    .RESET_B(net179),
    .Q(\ih.t.count[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6235_ (.CLK(clknet_leaf_23_clk),
    .D(\ih.t.next_count[23] ),
    .RESET_B(net179),
    .Q(\ih.t.count[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6236_ (.CLK(clknet_leaf_24_clk),
    .D(\ih.t.next_count[24] ),
    .RESET_B(net192),
    .Q(\ih.t.count[24] ));
 sky130_fd_sc_hd__dfrtp_2 _6237_ (.CLK(clknet_leaf_24_clk),
    .D(\ih.t.next_count[25] ),
    .RESET_B(net193),
    .Q(\ih.t.count[25] ));
 sky130_fd_sc_hd__dfrtp_1 _6238_ (.CLK(clknet_leaf_24_clk),
    .D(\ih.t.next_count[26] ),
    .RESET_B(net193),
    .Q(\ih.t.count[26] ));
 sky130_fd_sc_hd__dfrtp_1 _6239_ (.CLK(clknet_leaf_25_clk),
    .D(\ih.t.next_count[27] ),
    .RESET_B(net193),
    .Q(\ih.t.count[27] ));
 sky130_fd_sc_hd__dfrtp_2 _6240_ (.CLK(clknet_leaf_25_clk),
    .D(\ih.t.next_count[28] ),
    .RESET_B(net194),
    .Q(\ih.t.count[28] ));
 sky130_fd_sc_hd__dfrtp_1 _6241_ (.CLK(clknet_leaf_26_clk),
    .D(\ih.t.next_count[29] ),
    .RESET_B(net194),
    .Q(\ih.t.count[29] ));
 sky130_fd_sc_hd__dfrtp_1 _6242_ (.CLK(clknet_leaf_26_clk),
    .D(\ih.t.next_count[30] ),
    .RESET_B(net194),
    .Q(\ih.t.count[30] ));
 sky130_fd_sc_hd__dfrtp_1 _6243_ (.CLK(clknet_leaf_25_clk),
    .D(\ih.t.next_count[31] ),
    .RESET_B(net195),
    .Q(\ih.t.count[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6244_ (.CLK(clknet_leaf_37_clk),
    .D(_0015_),
    .RESET_B(net160),
    .Q(\cu.id.interrupt_requested ));
 sky130_fd_sc_hd__dfrtp_4 _6245_ (.CLK(clknet_leaf_3_clk),
    .D(_0227_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6246_ (.CLK(clknet_leaf_3_clk),
    .D(_0228_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6247_ (.CLK(clknet_leaf_1_clk),
    .D(_0229_),
    .RESET_B(net152),
    .Q(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6248_ (.CLK(clknet_leaf_42_clk),
    .D(_0230_),
    .RESET_B(net152),
    .Q(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6249_ (.CLK(clknet_leaf_1_clk),
    .D(_0231_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6250_ (.CLK(clknet_leaf_1_clk),
    .D(_0232_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6251_ (.CLK(clknet_leaf_1_clk),
    .D(_0233_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__dfstp_2 _6252_ (.CLK(clknet_leaf_1_clk),
    .D(_0234_),
    .SET_B(net155),
    .Q(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__dfstp_2 _6253_ (.CLK(clknet_leaf_2_clk),
    .D(_0235_),
    .SET_B(net155),
    .Q(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__dfstp_2 _6254_ (.CLK(clknet_leaf_2_clk),
    .D(_0236_),
    .SET_B(net155),
    .Q(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__dfstp_2 _6255_ (.CLK(clknet_leaf_2_clk),
    .D(_0237_),
    .SET_B(net154),
    .Q(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__dfstp_2 _6256_ (.CLK(clknet_leaf_2_clk),
    .D(_0238_),
    .SET_B(net156),
    .Q(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__dfstp_2 _6257_ (.CLK(clknet_leaf_3_clk),
    .D(_0239_),
    .SET_B(net156),
    .Q(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__dfstp_2 _6258_ (.CLK(clknet_leaf_4_clk),
    .D(_0240_),
    .SET_B(net157),
    .Q(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__dfstp_2 _6259_ (.CLK(clknet_leaf_4_clk),
    .D(_0241_),
    .SET_B(net157),
    .Q(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__dfstp_2 _6260_ (.CLK(clknet_leaf_23_clk),
    .D(_0242_),
    .SET_B(net191),
    .Q(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__dfstp_2 _6261_ (.CLK(clknet_leaf_23_clk),
    .D(_0243_),
    .SET_B(net193),
    .Q(\ih.t.timer_max[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6262_ (.CLK(clknet_leaf_23_clk),
    .D(_0244_),
    .RESET_B(net193),
    .Q(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6263_ (.CLK(clknet_leaf_23_clk),
    .D(_0245_),
    .RESET_B(net191),
    .Q(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6264_ (.CLK(clknet_leaf_23_clk),
    .D(_0246_),
    .RESET_B(net192),
    .Q(\ih.t.timer_max[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6265_ (.CLK(clknet_leaf_18_clk),
    .D(_0247_),
    .RESET_B(net193),
    .Q(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__dfstp_1 _6266_ (.CLK(clknet_leaf_23_clk),
    .D(_0248_),
    .SET_B(net191),
    .Q(\ih.t.timer_max[14] ));
 sky130_fd_sc_hd__dfstp_1 _6267_ (.CLK(clknet_leaf_23_clk),
    .D(_0249_),
    .SET_B(net191),
    .Q(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6268_ (.CLK(clknet_leaf_13_clk),
    .D(_0250_),
    .RESET_B(net174),
    .Q(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6269_ (.CLK(clknet_leaf_15_clk),
    .D(_0251_),
    .RESET_B(net175),
    .Q(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6270_ (.CLK(clknet_leaf_13_clk),
    .D(_0252_),
    .RESET_B(net174),
    .Q(\ih.t.timer_max[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6271_ (.CLK(clknet_leaf_15_clk),
    .D(_0253_),
    .RESET_B(net175),
    .Q(\ih.t.timer_max[3] ));
 sky130_fd_sc_hd__dfstp_1 _6272_ (.CLK(clknet_leaf_15_clk),
    .D(_0254_),
    .SET_B(net175),
    .Q(\ih.t.timer_max[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6273_ (.CLK(clknet_leaf_15_clk),
    .D(_0255_),
    .RESET_B(net175),
    .Q(\ih.t.timer_max[5] ));
 sky130_fd_sc_hd__dfstp_1 _6274_ (.CLK(clknet_leaf_15_clk),
    .D(_0256_),
    .SET_B(net177),
    .Q(\ih.t.timer_max[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6275_ (.CLK(clknet_leaf_15_clk),
    .D(_0257_),
    .RESET_B(net175),
    .Q(\ih.t.timer_max[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6276_ (.CLK(clknet_leaf_16_clk),
    .D(_0258_),
    .RESET_B(net180),
    .Q(\ih.t.timer_max[16] ));
 sky130_fd_sc_hd__dfrtp_2 _6277_ (.CLK(clknet_leaf_16_clk),
    .D(_0259_),
    .RESET_B(net178),
    .Q(\ih.t.timer_max[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6278_ (.CLK(clknet_leaf_16_clk),
    .D(_0260_),
    .RESET_B(net178),
    .Q(\ih.t.timer_max[18] ));
 sky130_fd_sc_hd__dfrtp_2 _6279_ (.CLK(clknet_leaf_16_clk),
    .D(_0261_),
    .RESET_B(net178),
    .Q(\ih.t.timer_max[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6280_ (.CLK(clknet_leaf_16_clk),
    .D(_0262_),
    .RESET_B(net178),
    .Q(\ih.t.timer_max[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6281_ (.CLK(clknet_leaf_17_clk),
    .D(_0263_),
    .RESET_B(net178),
    .Q(\ih.t.timer_max[21] ));
 sky130_fd_sc_hd__dfrtp_4 _6282_ (.CLK(clknet_leaf_16_clk),
    .D(_0264_),
    .RESET_B(net180),
    .Q(\ih.t.timer_max[22] ));
 sky130_fd_sc_hd__dfrtp_2 _6283_ (.CLK(clknet_leaf_16_clk),
    .D(_0265_),
    .RESET_B(net178),
    .Q(\ih.t.timer_max[23] ));
 sky130_fd_sc_hd__dfrtp_2 _6284_ (.CLK(clknet_leaf_36_clk),
    .D(_0266_),
    .RESET_B(net161),
    .Q(\cu.ir.idx[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6285_ (.CLK(clknet_leaf_38_clk),
    .D(_0267_),
    .RESET_B(net161),
    .Q(\cu.ir.idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6286_ (.CLK(clknet_leaf_37_clk),
    .D(_0268_),
    .RESET_B(net160),
    .Q(\cu.id.can_be_interrupted ));
 sky130_fd_sc_hd__dfrtp_4 _6287_ (.CLK(clknet_leaf_42_clk),
    .D(_0269_),
    .RESET_B(net152),
    .Q(\cu.id.opcode[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6288_ (.CLK(clknet_leaf_42_clk),
    .D(_0270_),
    .RESET_B(net152),
    .Q(\cu.id.opcode[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6289_ (.CLK(clknet_leaf_42_clk),
    .D(_0271_),
    .RESET_B(net153),
    .Q(\cu.id.opcode[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6290_ (.CLK(clknet_leaf_42_clk),
    .D(_0272_),
    .RESET_B(net152),
    .Q(\cu.id.alu_opcode[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6291_ (.CLK(clknet_leaf_42_clk),
    .D(_0273_),
    .RESET_B(net152),
    .Q(\cu.id.alu_opcode[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6292_ (.CLK(clknet_leaf_42_clk),
    .D(_0274_),
    .RESET_B(net152),
    .Q(\cu.id.alu_opcode[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6293_ (.CLK(clknet_leaf_42_clk),
    .D(_0275_),
    .RESET_B(net153),
    .Q(\cu.id.opcode[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6294_ (.CLK(clknet_leaf_42_clk),
    .D(_0276_),
    .RESET_B(net153),
    .Q(\cu.id.opcode[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6295_ (.CLK(clknet_leaf_0_clk),
    .D(_0277_),
    .RESET_B(net152),
    .Q(\cu.id.cb_opcode_z[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6296_ (.CLK(clknet_leaf_0_clk),
    .D(_0278_),
    .RESET_B(net152),
    .Q(\cu.id.cb_opcode_z[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6297_ (.CLK(clknet_leaf_41_clk),
    .D(_0279_),
    .RESET_B(net159),
    .Q(\cu.id.cb_opcode_z[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6298_ (.CLK(clknet_leaf_42_clk),
    .D(_0280_),
    .RESET_B(net152),
    .Q(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6299_ (.CLK(clknet_leaf_42_clk),
    .D(_0281_),
    .RESET_B(net153),
    .Q(\cu.id.cb_opcode_y[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6300_ (.CLK(clknet_leaf_38_clk),
    .D(_0282_),
    .RESET_B(net162),
    .Q(\cu.id.cb_opcode_y[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6301_ (.CLK(clknet_leaf_38_clk),
    .D(_0283_),
    .RESET_B(net160),
    .Q(\cu.id.cb_opcode_x[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6302_ (.CLK(clknet_leaf_36_clk),
    .D(_0284_),
    .RESET_B(net161),
    .Q(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6303_ (.CLK(clknet_leaf_7_clk),
    .D(_0285_),
    .RESET_B(net170),
    .Q(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6304_ (.CLK(clknet_leaf_9_clk),
    .D(_0286_),
    .RESET_B(net165),
    .Q(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6305_ (.CLK(clknet_leaf_9_clk),
    .D(_0287_),
    .RESET_B(net165),
    .Q(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6306_ (.CLK(clknet_leaf_9_clk),
    .D(_0288_),
    .RESET_B(net165),
    .Q(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6307_ (.CLK(clknet_leaf_7_clk),
    .D(_0289_),
    .RESET_B(net165),
    .Q(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6308_ (.CLK(clknet_leaf_31_clk),
    .D(_0290_),
    .RESET_B(net183),
    .Q(\cu.id.imm_i[13] ));
 sky130_fd_sc_hd__dfrtp_4 _6309_ (.CLK(clknet_leaf_20_clk),
    .D(_0291_),
    .RESET_B(net182),
    .Q(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__dfrtp_4 _6310_ (.CLK(clknet_leaf_31_clk),
    .D(_0292_),
    .RESET_B(net183),
    .Q(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6311_ (.CLK(clknet_leaf_37_clk),
    .D(_0004_),
    .RESET_B(net160),
    .Q(\cu.id.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6312_ (.CLK(clknet_leaf_37_clk),
    .D(_0005_),
    .RESET_B(net160),
    .Q(\cu.id.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6313_ (.CLK(clknet_leaf_37_clk),
    .D(_0006_),
    .RESET_B(net160),
    .Q(\cu.id.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6314_ (.CLK(clknet_leaf_37_clk),
    .D(net201),
    .RESET_B(net161),
    .Q(\cu.id.is_halted ));
 sky130_fd_sc_hd__dfrtp_4 _6315_ (.CLK(clknet_leaf_37_clk),
    .D(_0003_),
    .RESET_B(net160),
    .Q(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__dfrtp_1 _6316_ (.CLK(clknet_leaf_37_clk),
    .D(_0002_),
    .RESET_B(net160),
    .Q(\cu.id.is_interrupted ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(net159),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net159),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net159),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net159),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(net197),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 fanout162 (.A(net197),
    .X(net162));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net197),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net169),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(net181),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_2 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(net181),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net177),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 fanout177 (.A(net181),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_2 fanout181 (.A(net197),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net184),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 fanout185 (.A(net196),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net196),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net196),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(net196),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(net26),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\ih.ip_ed.prev_data ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\ih.t.count[30] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\cu.alu_f[5] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\cu.alu_f[3] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\mc.cc.count[0] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0097_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\cu.alu_f[4] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\ih.t.count[19] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\ih.t.next_count[19] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\ih.t.count[10] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\ih.t.next_count[10] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0217_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\ih.t.count[16] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\ih.t.count[13] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\ih.t.count[22] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\ih.t.count[4] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\ih.t.count[28] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\ih.t.count[25] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\mc.cc.count[3] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0099_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\cu.ir.idx[0] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\ih.t.count[9] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\cu.id.interrupt_requested ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\ih.t.count[7] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\mc.cc.count[1] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\ih.t.count[6] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\ih.t.count[21] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\ih.t.count[27] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\ih.t.count[24] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\ih.ih.ih.prev_data[11] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\cu.ir.idx[1] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\ih.t.count[15] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\cu.id.is_halted ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0001_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\ih.interrupt_source[1] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\cu.id.can_be_interrupted ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\cu.id.is_interrupted ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\ih.interrupt_source[2] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\cu.id.is_halted ),
    .X(net206));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(interrupt_gpio_in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(keypad_input[2]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(keypad_input[3]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(keypad_input[4]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(keypad_input[5]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(keypad_input[6]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(keypad_input[7]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(keypad_input[8]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(keypad_input[9]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(memory_data_in[0]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(memory_data_in[1]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(keypad_input[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(memory_data_in[2]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(memory_data_in[3]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(memory_data_in[4]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(memory_data_in[5]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(memory_data_in[6]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(memory_data_in[7]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(nrst),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(programmable_gpio_in[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(programmable_gpio_in[1]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(programmable_gpio_in[2]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(keypad_input[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(programmable_gpio_in[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(programmable_gpio_in[4]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(programmable_gpio_in[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(programmable_gpio_in[6]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(programmable_gpio_in[7]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input4 (.A(keypad_input[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(keypad_input[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(keypad_input[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(keypad_input[14]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(keypad_input[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(keypad_input[1]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 max_cap1 (.A(_2324_),
    .X(net237));
 sky130_fd_sc_hd__buf_1 max_cap140 (.A(_2873_),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_16 max_cap141 (.A(_2181_),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap142 (.A(net237),
    .X(net142));
 sky130_fd_sc_hd__buf_2 max_cap143 (.A(_0509_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 max_cap144 (.A(net238),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 max_cap146 (.A(net240),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 max_cap147 (.A(_0468_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 max_cap148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 max_cap149 (.A(net241),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 max_cap151 (.A(net243),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 max_cap3 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 max_cap5 (.A(_0335_),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(ss3[0]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(ss3[1]));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net102),
    .X(ss3[2]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(ss3[3]));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(ss3[4]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(ss3[5]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(ss3[6]));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(ss3[7]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(ss4[0]));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(ss4[1]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(ss4[2]));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(ss4[3]));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(ss4[4]));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net113),
    .X(ss4[5]));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(ss4[6]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(ss4[7]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(ss5[0]));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net117),
    .X(ss5[1]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(ss5[2]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(ss5[3]));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net120),
    .X(ss5[4]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(ss5[5]));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net122),
    .X(ss5[6]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(ss5[7]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(ss6[0]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(ss6[1]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(ss6[2]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(ss6[3]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(ss6[4]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(ss6[5]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(ss6[6]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(ss6[7]));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net132),
    .X(ss7[0]));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net133),
    .X(ss7[1]));
 sky130_fd_sc_hd__clkbuf_4 output134 (.A(net134),
    .X(ss7[2]));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net135),
    .X(ss7[3]));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net136),
    .X(ss7[4]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(ss7[5]));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net138),
    .X(ss7[6]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(ss7[7]));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net35),
    .X(memory_address_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(memory_address_out[10]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(memory_address_out[11]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(memory_address_out[12]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(memory_address_out[13]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(memory_address_out[14]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(memory_address_out[15]));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .X(memory_address_out[1]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(memory_address_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net44),
    .X(memory_address_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output45 (.A(net45),
    .X(memory_address_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(memory_address_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net47),
    .X(memory_address_out[6]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(memory_address_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net49),
    .X(memory_address_out[8]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(memory_address_out[9]));
 sky130_fd_sc_hd__clkbuf_4 output51 (.A(net51),
    .X(memory_data_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(memory_data_out[1]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(memory_data_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(memory_data_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .X(memory_data_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output56 (.A(net56),
    .X(memory_data_out[5]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(memory_data_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(memory_data_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output59 (.A(net59),
    .X(memory_wr));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(programmable_gpio_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(programmable_gpio_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(programmable_gpio_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(programmable_gpio_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(programmable_gpio_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(programmable_gpio_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(programmable_gpio_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(programmable_gpio_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(programmable_gpio_wr[0]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(programmable_gpio_wr[1]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(programmable_gpio_wr[2]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(programmable_gpio_wr[3]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(programmable_gpio_wr[4]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(programmable_gpio_wr[5]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(programmable_gpio_wr[6]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(programmable_gpio_wr[7]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(ss0[0]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(ss0[1]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(ss0[2]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(ss0[3]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(ss0[4]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(ss0[5]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(ss0[6]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(ss0[7]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(ss1[0]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(ss1[1]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(ss1[2]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net87),
    .X(ss1[3]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(ss1[4]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(ss1[5]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(ss1[6]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(ss1[7]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(ss2[0]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(ss2[1]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(ss2[2]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net95),
    .X(ss2[3]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(ss2[4]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(ss2[5]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(ss2[6]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(ss2[7]));
 sky130_fd_sc_hd__buf_1 wire145 (.A(_0985_),
    .X(net145));
 sky130_fd_sc_hd__buf_1 wire150 (.A(net242),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2 (.A(_1280_),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 wire4 (.A(_0481_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 wire6 (.A(_0448_),
    .X(net242));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7 (.A(_2895_),
    .X(net243));
endmodule

