* NGSPICE file created from z23.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt z23 clk interrupt_gpio_in keypad_input[0] keypad_input[10] keypad_input[11]
+ keypad_input[12] keypad_input[13] keypad_input[14] keypad_input[15] keypad_input[1]
+ keypad_input[2] keypad_input[3] keypad_input[4] keypad_input[5] keypad_input[6]
+ keypad_input[7] keypad_input[8] keypad_input[9] memory_address_out[0] memory_address_out[10]
+ memory_address_out[11] memory_address_out[12] memory_address_out[13] memory_address_out[14]
+ memory_address_out[15] memory_address_out[1] memory_address_out[2] memory_address_out[3]
+ memory_address_out[4] memory_address_out[5] memory_address_out[6] memory_address_out[7]
+ memory_address_out[8] memory_address_out[9] memory_data_in[0] memory_data_in[1]
+ memory_data_in[2] memory_data_in[3] memory_data_in[4] memory_data_in[5] memory_data_in[6]
+ memory_data_in[7] memory_data_out[0] memory_data_out[1] memory_data_out[2] memory_data_out[3]
+ memory_data_out[4] memory_data_out[5] memory_data_out[6] memory_data_out[7] memory_wr
+ nrst programmable_gpio_in[0] programmable_gpio_in[1] programmable_gpio_in[2] programmable_gpio_in[3]
+ programmable_gpio_in[4] programmable_gpio_in[5] programmable_gpio_in[6] programmable_gpio_in[7]
+ programmable_gpio_out[0] programmable_gpio_out[1] programmable_gpio_out[2] programmable_gpio_out[3]
+ programmable_gpio_out[4] programmable_gpio_out[5] programmable_gpio_out[6] programmable_gpio_out[7]
+ programmable_gpio_wr[0] programmable_gpio_wr[1] programmable_gpio_wr[2] programmable_gpio_wr[3]
+ programmable_gpio_wr[4] programmable_gpio_wr[5] programmable_gpio_wr[6] programmable_gpio_wr[7]
+ ss0[0] ss0[1] ss0[2] ss0[3] ss0[4] ss0[5] ss0[6] ss0[7] ss1[0] ss1[1] ss1[2] ss1[3]
+ ss1[4] ss1[5] ss1[6] ss1[7] ss2[0] ss2[1] ss2[2] ss2[3] ss2[4] ss2[5] ss2[6] ss2[7]
+ ss3[0] ss3[1] ss3[2] ss3[3] ss3[4] ss3[5] ss3[6] ss3[7] ss4[0] ss4[1] ss4[2] ss4[3]
+ ss4[4] ss4[5] ss4[6] ss4[7] ss5[0] ss5[1] ss5[2] ss5[3] ss5[4] ss5[5] ss5[6] ss5[7]
+ ss6[0] ss6[1] ss6[2] ss6[3] ss6[4] ss6[5] ss6[6] ss6[7] ss7[0] ss7[1] ss7[2] ss7[3]
+ ss7[4] ss7[5] ss7[6] ss7[7] vccd1 vssd1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5417__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3155_ cu.id.alu_opcode\[0\] vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__clkbuf_4
X_3086_ _2752_ _2822_ ih.t.count\[9\] vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5968__A1 _2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _0588_ _1059_ _0606_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5727_ _2518_ mc.cl.next_data\[2\] _2111_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__and3_1
XANTENNA__5485__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5658_ net91 _1329_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__or2_1
X_4609_ _1652_ mc.cc.count\[3\] mc.cc.enable_edge_detector.prev_data vssd1 vssd1 vccd1
+ vccd1 _1653_ sky130_fd_sc_hd__or3b_2
X_5589_ _2169_ _2398_ _2405_ _2136_ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4829__B cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5350__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output56_A net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4960_ _1799_ _1942_ _1948_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4891_ _2920_ cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3911_ _0973_ _0329_ _0379_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__nor3_1
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5512_ net67 _1638_ _2279_ net66 vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3594__D1 _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3820__B_N _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3773_ cu.reg_file.reg_a\[5\] _0625_ _0628_ cu.reg_file.reg_mem\[13\] _0848_ vssd1
+ vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5886__A0 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5443_ _2139_ _2247_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__nand2_1
X_5374_ _2230_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_4325_ cu.reg_file.reg_sp\[3\] _0993_ _1344_ cu.id.cb_opcode_y\[0\] _1324_ vssd1
+ vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__a221o_1
X_4256_ _1323_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5260__S _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3207_ _2897_ _2932_ _2935_ _2937_ _2943_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__o2111a_1
X_4187_ _1234_ _1182_ _1023_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__o21a_1
X_3138_ cu.id.opcode\[6\] vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__clkbuf_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _2756_ _2806_ ih.t.count\[15\] vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5565__C1 _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5580__A2 _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3591__A1 cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3591__B2 cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5345__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3654__A _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5090_ cu.reg_file.reg_d\[4\] _2047_ _2039_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__mux2_1
X_4110_ _1013_ _1182_ _1023_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4041_ _0607_ _1114_ _0632_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__o21a_1
XANTENNA__5080__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5992_ clknet_leaf_34_clk _0030_ net163 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4943_ _1932_ _1933_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4874_ cu.pc.pc_o\[5\] _1870_ _1815_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__mux2_1
XANTENNA__5020__A1 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3825_ _0737_ _0752_ _0898_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a31o_1
XANTENNA__3031__B1 ih.t.timer_max\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3756_ cu.reg_file.reg_mem\[15\] _0640_ _0830_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5970__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3582__A1 cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3582__B2 cu.reg_file.reg_a\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5426_ _2022_ net69 _2260_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__mux2_1
X_3687_ _0762_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__inv_2
X_5357_ _2220_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
X_5288_ _1369_ _2179_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__and2_4
X_4308_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__clkbuf_4
X_4239_ _0343_ _1295_ _1298_ _1299_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__a221o_1
XANTENNA__4826__C cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4842__B cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3458__B _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5011__A1 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3573__B2 cu.reg_file.reg_e\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap5 _0335_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5002__A1 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4590_ _1415_ _1630_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__or3_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3610_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[3\] vssd1 vssd1 vccd1 vccd1 _0686_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3541_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6260_ clknet_leaf_23_clk _0242_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[8\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__5688__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3472_ _0371_ _0376_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__or2_1
X_6191_ clknet_leaf_22_clk _0224_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5211_ _0619_ ih.gpio_interrupt_mask\[0\] _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__mux2_1
X_5142_ _2081_ cu.reg_file.reg_h\[6\] _2069_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__mux2_1
XANTENNA__4927__B _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5073_ _2034_ _1792_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__nor2_8
X_4024_ _1032_ _1095_ _1097_ _0770_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5975_ clknet_leaf_33_clk _0012_ net163 vssd1 vssd1 vccd1 vccd1 cu.alu_f\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4926_ _2920_ _1521_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__or2_1
X_4857_ _1853_ _1854_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3278__B _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3808_ cu.reg_file.reg_b\[2\] _0426_ _0429_ cu.reg_file.reg_d\[2\] vssd1 vssd1 vccd1
+ vccd1 _0884_ sky130_fd_sc_hd__a22o_1
XANTENNA__5493__B _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4752__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4788_ _2953_ _0339_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__nor2_2
X_3739_ _0813_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__nand2_1
X_5409_ _1075_ net134 _2248_ vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4268__C1 _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4853__A _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3794__B2 cu.reg_file.reg_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3794__A1 cu.reg_file.reg_a\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5535__A2 _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5299__A1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4763__A _1739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5578__B _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2972_ net10 vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5760_ cu.reg_file.reg_sp\[3\] _2534_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4711_ ih.t.count\[25\] ih.t.count\[26\] _1723_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__and3_1
X_5691_ mc.cl.next_data\[11\] _2359_ _2490_ _2499_ vssd1 vssd1 vccd1 vccd1 _2500_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3785__A1 cu.id.imm_i\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4642_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] ih.t.count\[3\] vssd1 vssd1
+ vccd1 vccd1 _1680_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _2702_ _1052_ _1623_ _2697_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__a22o_1
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6312_ clknet_leaf_37_clk _0005_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3524_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__inv_2
X_6243_ clknet_leaf_25_clk ih.t.next_count\[31\] net195 vssd1 vssd1 vccd1 vccd1 ih.t.count\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4938__A cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3455_ _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__buf_2
X_6174_ clknet_leaf_21_clk _0208_ net184 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_3386_ _0455_ _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5125_ _2070_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__clkbuf_1
X_5056_ cu.reg_file.reg_c\[0\] _2022_ _2025_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5462__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4007_ _1076_ _1077_ _1080_ _0517_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__o31a_1
XFILLER_0_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5958_ cu.id.imm_i\[10\] _2391_ _2686_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__mux2_1
X_4909_ _1900_ _1901_ _1798_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3776__A1 cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3776__B2 cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4973__A0 cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5889_ _2651_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold30 ih.t.count\[7\] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6020__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4583__A _1561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4716__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3519__B2 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output86_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3662__A _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5141__A0 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4477__B _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6108__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _0308_ _0315_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__nor2_1
XANTENNA__5692__B2 _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3171_ cu.id.opcode\[7\] cu.id.opcode\[6\] vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__and2b_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3207__B1 _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5812_ _1623_ _2594_ _2545_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5743_ _2533_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__3758__A1 cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3758__B2 cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2955_ mc.rw.state\[2\] _2695_ mc.rw.state\[0\] vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5674_ cu.reg_file.reg_mem\[7\] _2486_ _1739_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__mux2_1
XANTENNA__4707__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4625_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4556_ _1296_ _1607_ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__a21o_1
X_3507_ _0321_ _0322_ _0328_ _0334_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__or4_4
XANTENNA__5263__S _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4487_ cu.reg_file.reg_h\[3\] _1316_ _1312_ cu.reg_file.reg_b\[3\] _1543_ vssd1 vssd1
+ vccd1 vccd1 _1544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5132__A0 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6226_ clknet_leaf_15_clk ih.t.next_count\[14\] net177 vssd1 vssd1 vccd1 vccd1 ih.t.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3438_ _0384_ _0392_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__nand2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ clknet_leaf_20_clk _0191_ net172 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4486__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3369_ cu.id.cb_opcode_y\[0\] _0361_ _0444_ _0343_ _0322_ vssd1 vssd1 vccd1 vccd1
+ _0445_ sky130_fd_sc_hd__a221o_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _2059_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5435__A1 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6088_ clknet_leaf_24_clk _0122_ net190 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_4
X_5039_ _2013_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3945__C_N _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3749__B2 cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5371__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 memory_address_out[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__4578__A _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[7] sky130_fd_sc_hd__clkbuf_4
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 memory_data_out[2] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 ss2[5] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 ss1[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5674__A1 _2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5426__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output124_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5348__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5362__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4165__A1 _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4410_ cu.pc.pc_o\[7\] _1322_ _1315_ cu.reg_file.reg_e\[7\] _1470_ vssd1 vssd1 vccd1
+ vccd1 _1471_ sky130_fd_sc_hd__a221o_1
X_5390_ _1075_ net126 _2237_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4341_ _1382_ _1398_ _1399_ _1405_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__a31o_2
XANTENNA__5083__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3912__A1 _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4272_ cu.reg_file.reg_c\[1\] _1281_ _1338_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4468__A2 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6011_ clknet_leaf_5_clk _0049_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3223_ _2902_ _2884_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__and2_1
XANTENNA__5417__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ _2888_ _2889_ _2890_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3085_ ih.t.count\[9\] _2752_ _2822_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout155_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3987_ _1060_ _0588_ _0599_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__and3_1
X_5726_ net19 _2519_ _2523_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5657_ net99 _2193_ _2469_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__a21o_1
X_4608_ mc.cc.count\[2\] mc.cc.count\[1\] mc.cc.count\[0\] vssd1 vssd1 vccd1 vccd1
+ _1652_ sky130_fd_sc_hd__or3_1
X_5588_ ih.gpio_interrupt_mask\[3\] _2326_ _2404_ _2125_ _2327_ vssd1 vssd1 vccd1
+ vccd1 _2405_ sky130_fd_sc_hd__a221o_1
X_4539_ _1296_ _1591_ _1592_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__a21o_1
XANTENNA__5105__A0 cu.reg_file.reg_e\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5656__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5656__B2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6209_ clknet_leaf_9_clk net7 net169 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5895__A1 _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output49_A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4890_ _2920_ cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__nor2_1
X_3910_ _0526_ net145 vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__nand2_4
XANTENNA__4490__B _1545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5078__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3841_ _0401_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4386__A1 cu.reg_file.reg_c\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3772_ cu.pc.pc_o\[13\] _0740_ _0846_ _0847_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__a211o_1
X_5511_ net64 _2277_ _2179_ net65 vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5335__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4138__A1 _0916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5442_ _2271_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
X_5373_ _1188_ net119 _2226_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__mux2_1
XANTENNA__4649__C _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4324_ cu.reg_file.reg_l\[3\] _1317_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4255_ _1268_ _1302_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__nand2_2
X_3206_ _2940_ _2942_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__nor2_1
X_4186_ _1127_ _1236_ _1238_ _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__a31o_2
X_3137_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[0\] cu.id.alu_opcode\[3\] vssd1 vssd1
+ vccd1 vccd1 _2874_ sky130_fd_sc_hd__and3_2
XFILLER_0_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3068_ ih.t.timer_max\[15\] _2755_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5709_ net8 _1650_ _2488_ _2513_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5326__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5877__A1 _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4591__A _1455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4368__A1 cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4368__B2 _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4540__A1 cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4040_ _0610_ _1111_ _1112_ _1113_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5991_ clknet_leaf_34_clk _0029_ net163 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_4942_ _1918_ _1923_ _1919_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4873_ _1862_ _1869_ _1809_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5556__B1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3824_ _0892_ _0895_ _0898_ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3755_ cu.reg_file.reg_b\[7\] _0426_ _0429_ cu.reg_file.reg_d\[7\] vssd1 vssd1 vccd1
+ vccd1 _0831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3686_ _0694_ _0701_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5425_ _2139_ _2180_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5356_ _1190_ net112 _2215_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5271__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4307_ _1306_ _1362_ _1367_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__o21a_2
X_5287_ _1329_ _1354_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__nor2_2
XANTENNA__3580__A cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4238_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4169_ _0829_ _0838_ _1060_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4522__B2 cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4522__A1 cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4586__A _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5538__B1 _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4210__B1 _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5356__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3540_ _0518_ _0568_ _0571_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__or4b_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5210_ _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__clkbuf_4
X_3471_ _0399_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nor2_2
X_6190_ clknet_leaf_22_clk _0223_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5141_ _1624_ _1126_ _2066_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5072_ _1790_ _0348_ _0351_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__or3_2
XFILLER_0_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4023_ _0918_ _1096_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5974_ clknet_2_1__leaf_clk _0011_ net161 vssd1 vssd1 vccd1 vccd1 cu.alu_f\[4\] sky130_fd_sc_hd__dfrtp_1
X_4925_ _1521_ _1907_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4856_ _1841_ _1844_ _1842_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3807_ cu.reg_file.reg_sp\[10\] _0636_ _0748_ cu.reg_file.reg_h\[2\] vssd1 vssd1
+ vccd1 vccd1 _0883_ sky130_fd_sc_hd__a22o_1
XANTENNA__5266__S _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4787_ _0343_ _1299_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3738_ _0801_ _0812_ _0798_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3669_ cu.pc.pc_o\[8\] _0740_ _0742_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5408_ _2250_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4504__A1 cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4504__B2 cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5339_ _1190_ net104 _2206_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__mux2_1
XANTENNA__4853__B cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6297__RESET_B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire145 _0985_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_1
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5940__A0 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3932__B _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3379__B _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2971_ net4 vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4710_ net222 _1723_ _1725_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[25\] sky130_fd_sc_hd__a21oi_1
X_5690_ ih.t.timer_max\[27\] _2151_ _2320_ ih.t.timer_max\[11\] vssd1 vssd1 vccd1
+ vccd1 _2499_ sky130_fd_sc_hd__a22oi_1
X_4641_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] ih.t.count\[3\] vssd1 vssd1
+ vccd1 vccd1 _1679_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5086__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4572_ _0516_ _1230_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__nor2_8
XFILLER_0_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6311_ clknet_leaf_37_clk _0004_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3523_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__buf_2
X_6242_ clknet_leaf_26_clk ih.t.next_count\[30\] net194 vssd1 vssd1 vccd1 vccd1 ih.t.count\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3454_ _0519_ _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__or2_1
XANTENNA__4938__B _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4498__B1 _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6173_ clknet_leaf_21_clk _0207_ net184 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_3385_ _2896_ _0324_ _2912_ _0346_ _2949_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5124_ _2067_ cu.reg_file.reg_h\[0\] _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout185_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5055_ _2002_ _2024_ _2951_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__o21a_4
XANTENNA__4954__A _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4006_ _0817_ _1078_ _1079_ _0810_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _2688_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4908_ _1900_ _1901_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__or2_1
XANTENNA__3776__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5888_ _1191_ ih.t.timer_max\[5\] _2645_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4839_ cu.pc.pc_o\[3\] _1826_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold20 ih.t.count\[16\] vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 mc.cc.count\[1\] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5634__S _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output79_A net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__A1 _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3170_ cu.id.alu_opcode\[0\] cu.id.alu_opcode\[3\] cu.id.alu_opcode\[1\] vssd1 vssd1
+ vccd1 vccd1 _2907_ sky130_fd_sc_hd__and3b_1
XANTENNA__4774__A _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5811_ _2592_ _2593_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5742_ _0296_ _0469_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__or2_1
XANTENNA__3758__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2954_ mc.rw.state\[1\] vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5673_ _2482_ _2483_ _2485_ _1641_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__o22a_4
XFILLER_0_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4624_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4555_ cu.id.imm_i\[15\] _1294_ _1297_ cu.pc.pc_o\[15\] _1489_ vssd1 vssd1 vccd1
+ vccd1 _1608_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4949__A cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3506_ _0341_ _0443_ _0336_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__a21o_1
X_4486_ cu.pc.pc_o\[11\] _1321_ _1314_ cu.reg_file.reg_d\[3\] _1542_ vssd1 vssd1 vccd1
+ vccd1 _1543_ sky130_fd_sc_hd__a221o_1
X_6225_ clknet_leaf_15_clk ih.t.next_count\[13\] net175 vssd1 vssd1 vccd1 vccd1 ih.t.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_3437_ alu.Cin _0512_ _0510_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__a21o_1
XANTENNA__5132__A1 _1089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6156_ clknet_leaf_19_clk _0190_ net180 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _0442_ _0437_ _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__a21o_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ cu.reg_file.reg_e\[2\] _1074_ _2056_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__mux2_1
X_6087_ clknet_leaf_8_clk _0121_ net168 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_4
X_3299_ _0373_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__nand2_1
X_5038_ cu.reg_file.reg_b\[3\] _2012_ _2006_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3749__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5371__A1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 memory_address_out[2] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 ss0[0] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 memory_data_out[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5123__A1 _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 ss1[3] sky130_fd_sc_hd__clkbuf_4
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 ss2[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5584__A_N _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3437__A1 alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5362__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ _1400_ _1403_ _1404_ _1371_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4271_ cu.reg_file.reg_e\[1\] _1283_ _1285_ cu.reg_file.reg_l\[1\] _1337_ vssd1 vssd1
+ vccd1 vccd1 _1338_ sky130_fd_sc_hd__a221o_1
X_6010_ clknet_leaf_7_clk _0048_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3222_ _2892_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__inv_2
X_3153_ cu.id.alu_opcode\[3\] cu.id.alu_opcode\[1\] vssd1 vssd1 vccd1 vccd1 _2890_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3084_ ih.t.timer_max\[9\] _2751_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__nand2_1
XANTENNA__3428__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4009__A _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3986_ _0575_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__clkbuf_4
X_5725_ _2518_ mc.cl.next_data\[1\] _2111_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3600__A1 cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5656_ net131 _2235_ _2246_ net139 vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__a22o_1
X_4607_ mc.rw.state\[2\] mc.rw.state\[1\] mc.rw.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _1651_ sky130_fd_sc_hd__nor3_1
XFILLER_0_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5587_ mc.cl.next_data\[3\] _2313_ net142 _2403_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4398__B _1455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4538_ cu.id.imm_i\[14\] _1295_ _1298_ cu.pc.pc_o\[14\] _1489_ vssd1 vssd1 vccd1
+ vccd1 _1592_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4469_ cu.reg_file.reg_sp\[10\] _0992_ _1344_ cu.id.imm_i\[10\] _1324_ vssd1 vssd1
+ vccd1 vccd1 _1527_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5105__A1 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6208_ clknet_leaf_8_clk net6 net169 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4864__B1 cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6139_ clknet_leaf_20_clk _0173_ net182 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_4
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5041__A0 cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4304__C1 _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3840_ _0774_ _0775_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__and2_2
XANTENNA__5032__A0 cu.reg_file.reg_b\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5583__A1 ih.t.timer_max\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3771_ cu.reg_file.reg_b\[5\] _0743_ _0624_ cu.reg_file.reg_sp\[13\] vssd1 vssd1
+ vccd1 vccd1 _0847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5510_ net68 _1648_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5441_ _2022_ net74 _2270_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5372_ _2229_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__clkbuf_1
X_4323_ cu.id.cb_opcode_y\[0\] _1295_ _1298_ cu.pc.pc_o\[3\] _1305_ vssd1 vssd1 vccd1
+ vccd1 _1388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3649__B2 cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3649__A1 cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4254_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__buf_2
X_3205_ _2902_ _2936_ _2885_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__and4_1
X_4185_ _0387_ _1234_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3136_ _2745_ _2869_ _2871_ net140 net202 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a32o_1
X_3067_ ih.t.count\[16\] _2804_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__xnor2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4074__A1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4173__S _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5574__A1 _2391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5708_ _2512_ _1643_ cu.reg_file.reg_mem\[15\] _1646_ vssd1 vssd1 vccd1 vccd1 _2513_
+ sky130_fd_sc_hd__a2bb2o_1
X_3969_ _0611_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5326__A1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5639_ net106 _2204_ _2452_ _1401_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4837__A0 cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4591__B _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3812__B2 cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3812__A1 cu.reg_file.reg_b\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5014__A0 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4368__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5565__B2 ih.t.timer_max\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3000__B net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4540__A2 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3951__A _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output61_A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ clknet_leaf_34_clk _0028_ net163 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[12\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__5089__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4941_ _2920_ cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3803__B2 cu.reg_file.reg_sp\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4872_ _1867_ _1868_ _1799_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__mux2_1
XANTENNA__5005__A0 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5556__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3823_ _0747_ _0751_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3754_ cu.reg_file.reg_sp\[15\] _0636_ _0748_ cu.reg_file.reg_h\[7\] vssd1 vssd1
+ vccd1 vccd1 _0830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3685_ _0758_ _0760_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__nand2_1
XANTENNA__3845__B _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5424_ _2259_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5355_ _2219_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4306_ _1348_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__inv_2
X_5286_ _2178_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4237_ _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3580__B _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4168_ _1144_ _1160_ _1237_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3119_ _2797_ _2799_ _2800_ _2856_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__or4_1
X_4099_ _0948_ _0959_ _0773_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4867__A _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4522__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3797__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4210__A1 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3470_ _0296_ _0528_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__or2_2
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5140_ _2080_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_1
X_5071_ _2033_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5474__A0 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4022_ _0768_ _0772_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5973_ clknet_leaf_33_clk _0010_ net164 vssd1 vssd1 vccd1 vccd1 cu.alu_f\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4924_ _1916_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5529__A1 _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4855_ _1851_ _1852_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4786_ _1299_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3806_ cu.id.imm_i\[10\] _0739_ _0881_ _0653_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__a22o_2
X_3737_ _0801_ _0812_ _0798_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__or3_1
X_3668_ cu.reg_file.reg_b\[0\] _0743_ _0624_ cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1
+ vccd1 _0744_ sky130_fd_sc_hd__a22o_1
X_5407_ _1052_ net133 _2248_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__mux2_1
XANTENNA__5701__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3599_ cu.reg_file.reg_l\[4\] _0621_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__a21o_1
X_5338_ _2210_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__clkbuf_1
X_5269_ _1642_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5217__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5940__A1 _2391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4259__A1 cu.reg_file.reg_e\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5920__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4259__B2 cu.reg_file.reg_l\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2970_ net9 vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__inv_2
XANTENNA__4431__A1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5367__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4640_ _1678_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3676__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4195__B1 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4571_ _2702_ _0619_ _1622_ _2697_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__a22o_1
X_6310_ clknet_leaf_31_clk _0292_ net183 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__6202__D net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5989__RESET_B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3522_ _0440_ _0589_ _0591_ _0593_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__o41a_4
X_6241_ clknet_leaf_26_clk ih.t.next_count\[29\] net194 vssd1 vssd1 vccd1 vccd1 ih.t.count\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3453_ _0400_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__or2_1
X_6172_ clknet_leaf_21_clk _0206_ net182 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4498__B2 cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4498__A1 cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3384_ _0345_ _0450_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__or3b_2
X_5123_ _2066_ _2068_ _2951_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__a21bo_4
X_5054_ _2004_ _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__nor2_1
XANTENNA__4954__B cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4005_ _0817_ _0808_ _0776_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5956_ cu.id.imm_i\[9\] _2372_ _2686_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5887_ _2650_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
X_4907_ _1885_ _1888_ _1886_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4838_ _1837_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5277__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4769_ _1300_ _1644_ _1268_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__o21a_1
XANTENNA__5922__A1 _2372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold32 ih.t.count\[6\] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 ih.t.count\[30\] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 ih.t.count\[13\] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5438__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__C _1598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4880__A _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3496__A alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3943__B _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4120__A _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3662__C _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4774__B _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5810_ _2583_ _2586_ _2584_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5741_ _1007_ _0981_ _0989_ _0994_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__or4b_2
XANTENNA__4404__B2 cu.reg_file.reg_l\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5672_ _1649_ _2484_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4623_ _0315_ _1658_ _1659_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__or3b_4
X_4554_ cu.reg_file.reg_b\[7\] net144 _1284_ cu.reg_file.reg_h\[7\] _1606_ vssd1 vssd1
+ vccd1 vccd1 _1607_ sky130_fd_sc_hd__a221o_1
XANTENNA__3391__A1 _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3505_ cu.reg_file.reg_l\[2\] _0422_ _0577_ _0579_ _0580_ vssd1 vssd1 vccd1 vccd1
+ _0581_ sky130_fd_sc_hd__a2111o_1
XANTENNA__4668__C _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6224_ clknet_leaf_15_clk ih.t.next_count\[12\] net175 vssd1 vssd1 vccd1 vccd1 ih.t.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4485_ cu.reg_file.reg_sp\[11\] _0992_ _1343_ cu.id.imm_i\[11\] _1324_ vssd1 vssd1
+ vccd1 vccd1 _1542_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _0395_ _0400_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6155_ clknet_leaf_11_clk _0189_ net168 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _0328_ _0334_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__or2_1
XANTENNA__4965__A _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6086_ clknet_leaf_13_clk _0120_ net173 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _2058_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
X_5037_ _1187_ _1222_ _2002_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__mux2_1
X_3298_ cu.id.cb_opcode_y\[1\] vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5939_ _2678_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4205__A _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 memory_address_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 memory_data_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[6] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 ss0[1] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 ss2[7] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 ss1[4] sky130_fd_sc_hd__clkbuf_4
XANTENNA__4594__B _1372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3003__B net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4115__A _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output91_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4270_ cu.reg_file.reg_a\[1\] _1276_ _1287_ cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1
+ vccd1 _1337_ sky130_fd_sc_hd__a22o_1
X_3221_ _2925_ _2932_ _2904_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__o21ai_1
X_3152_ cu.id.opcode\[0\] cu.id.opcode\[2\] cu.id.opcode\[1\] vssd1 vssd1 vccd1 vccd1
+ _2889_ sky130_fd_sc_hd__and3_1
X_3083_ ih.t.count\[10\] _2820_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3428__A2 _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3985_ _0603_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__inv_2
X_5724_ net18 _2519_ _2522_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3600__A2 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5655_ _2468_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606_ _1649_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5586_ _1666_ _2401_ _2402_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4537_ cu.reg_file.reg_b\[6\] _1281_ _1285_ cu.reg_file.reg_h\[6\] _1590_ vssd1 vssd1
+ vccd1 vccd1 _1591_ sky130_fd_sc_hd__a221o_1
X_4468_ _1521_ _1485_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__o21a_1
X_6207_ clknet_leaf_12_clk net5 net169 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3419_ net147 _0473_ _0479_ _0463_ _0458_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__o2111a_4
X_4399_ _1455_ _1459_ _1460_ _1371_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__a22o_1
X_6138_ clknet_leaf_28_clk _0172_ net187 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4864__A1 cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6069_ clknet_leaf_12_clk _0103_ net174 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6039__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5813__A0 cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4589__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3355__A1 cu.reg_file.reg_c\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3355__B2 cu.reg_file.reg_e\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5501__C1 _1660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3014__A ih.t.timer_max\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5804__A0 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4771__C _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3770_ cu.reg_file.reg_d\[5\] _0488_ _0741_ cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1
+ vccd1 _0846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5375__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5440_ _2139_ _2236_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5371_ _1075_ net118 _2226_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6210__D net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4322_ _1271_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4253_ _1319_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nor2_2
X_3204_ cu.id.opcode\[2\] cu.id.opcode\[1\] _2875_ _2876_ vssd1 vssd1 vccd1 vccd1
+ _2941_ sky130_fd_sc_hd__and4bb_2
X_4184_ _0701_ _1245_ _1253_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__a21o_1
X_3135_ net1 _2872_ _2870_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__nor3_1
X_3066_ ih.t.timer_max\[16\] _2756_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__xor2_1
XANTENNA__6132__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5271__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout160_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3968_ _0599_ _0603_ _0606_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ mc.cl.next_data\[15\] _2359_ _2490_ _2511_ vssd1 vssd1 vccd1 vccd1 _2512_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_9_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3585__B2 cu.reg_file.reg_l\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5285__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3899_ _0359_ _0973_ _0364_ _0974_ _0296_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5638_ net90 _1330_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5569_ _2169_ _2379_ _2386_ _2136_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3888__A2 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3812__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3567__A1_N _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5014__A1 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3951__B _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output54_A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4940_ _1929_ _1930_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__nor2_1
XANTENNA__3803__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4871_ _1144_ _1862_ _1795_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__mux2_1
XANTENNA__5005__A1 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6205__D net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3822_ _0896_ _0897_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__nand2_2
XANTENNA__5556__A2 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ cu.id.imm_i\[15\] _0739_ _0828_ _0653_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3684_ _0714_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5423_ net68 _2085_ _2258_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__mux2_1
XANTENNA__4516__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5354_ _1188_ net111 _2215_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _2701_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5285_ net83 _1260_ _2170_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__mux2_1
XANTENNA__4819__A1 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6313__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4236_ _2946_ _1303_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4167_ _0617_ _1050_ _1073_ _1089_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__or4_1
X_3118_ _2802_ _2803_ _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__or3_1
XANTENNA__5244__A1 _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4098_ _0916_ _0946_ _1171_ _1032_ _0918_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__o221a_1
X_3049_ _2761_ _2785_ ih.t.count\[23\] vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4867__B cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4586__C _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3797__B2 cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3797__A1 cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5538__A2 _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4123__A _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5070_ cu.reg_file.reg_c\[7\] _1260_ _2025_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__mux2_1
XANTENNA__5474__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4021_ _1093_ _1094_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nor2_1
XANTENNA__3485__B1 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ clknet_leaf_36_clk _0009_ net161 vssd1 vssd1 vccd1 vccd1 cu.alu_f\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4923_ cu.pc.pc_o\[9\] _1915_ _1815_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__mux2_1
XANTENNA__3788__A1 cu.reg_file.reg_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4732__S _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4017__B _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4854_ _0374_ cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__nand2_1
X_4785_ net200 _1787_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__nor2_1
X_3805_ cu.reg_file.reg_a\[2\] _0625_ _0628_ cu.reg_file.reg_mem\[10\] _0880_ vssd1
+ vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3736_ _0802_ _0804_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__or3_2
XFILLER_0_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4752__A3 _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3667_ _0464_ _0480_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__and2_2
X_5406_ _2249_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5701__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3598_ cu.reg_file.reg_c\[4\] _0485_ _0489_ cu.reg_file.reg_e\[4\] vssd1 vssd1 vccd1
+ vccd1 _0674_ sky130_fd_sc_hd__a22o_1
X_5337_ _1188_ net103 _2206_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__mux2_1
XANTENNA__4179__S _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5268_ _2168_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5799__A cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4219_ _1286_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__buf_2
X_5199_ net210 _2708_ _2119_ mc.cc.enable_edge_detector.prev_data vssd1 vssd1 vccd1
+ vccd1 _0097_ sky130_fd_sc_hd__a22o_1
XANTENNA__5311__B _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4976__B1 cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5153__A0 cu.reg_file.reg_l\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4118__A _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5392__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4195__B2 _1027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4195__A1 _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4570_ _0824_ _0819_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__and2_4
X_3521_ _0293_ _0596_ _0440_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_3_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5144__A0 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6240_ clknet_leaf_25_clk ih.t.next_count\[28\] net194 vssd1 vssd1 vccd1 vccd1 ih.t.count\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_3452_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__buf_2
X_3383_ _2889_ _0301_ _2933_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or3_1
X_6171_ clknet_leaf_38_clk _0205_ net161 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5122_ _0352_ _1792_ _1790_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__or3b_1
X_5053_ _0350_ _0358_ _0366_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__or3_1
X_4004_ _0808_ _0810_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5955_ _2687_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__clkbuf_1
X_5886_ _1189_ ih.t.timer_max\[4\] _2645_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4906_ _1898_ _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__or2_1
X_4837_ cu.pc.pc_o\[2\] _1836_ _1815_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4768_ net206 _1775_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4699_ _1717_ _1718_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[21\] sky130_fd_sc_hd__nor2_1
XANTENNA__5293__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3719_ _0788_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5135__A0 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5686__B2 ih.t.timer_max\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 ih.t.count\[22\] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5438__A1 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 cu.alu_f\[5\] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 ih.t.count\[21\] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5610__A1 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4880__B cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4401__A _1455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5126__A0 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5677__B2 ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3017__A ih.t.timer_max\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__A1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5232__A _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5601__A1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5740_ _2530_ _1050_ _2116_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__mux2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5671_ net15 _2345_ _2369_ net8 vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__a22o_1
X_4622_ _1653_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4553_ cu.reg_file.reg_d\[7\] _1282_ _1286_ cu.reg_file.reg_sp\[15\] vssd1 vssd1
+ vccd1 vccd1 _1606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4484_ cu.pc.pc_o\[11\] _1485_ _1540_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__o21a_1
X_3504_ cu.reg_file.reg_mem\[2\] _0418_ _0419_ cu.reg_file.reg_h\[2\] vssd1 vssd1
+ vccd1 vccd1 _0580_ sky130_fd_sc_hd__a22o_1
X_6223_ clknet_leaf_15_clk ih.t.next_count\[11\] net175 vssd1 vssd1 vccd1 vccd1 ih.t.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3435_ alu.Cin _0510_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6154_ clknet_leaf_13_clk _0188_ net173 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4340__A1 _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3366_ _0321_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
XANTENNA__4965__B cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6085_ clknet_leaf_12_clk _0119_ net174 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout190_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ cu.id.cb_opcode_y\[2\] vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__buf_4
X_5105_ cu.reg_file.reg_e\[1\] _1051_ _2056_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__mux2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _2011_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_1
X_5938_ _0340_ _2372_ _2666_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__mux2_1
XANTENNA__3603__B1 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5869_ _2161_ ih.t.timer_max\[12\] _2636_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__mux2_1
XANTENNA__5356__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5659__B2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5659__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 memory_address_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 memory_data_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 ss1[5] sky130_fd_sc_hd__clkbuf_4
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 ss0[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5052__A _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4891__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5926__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output84_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3220_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3151_ _2875_ _2876_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__nor2_2
X_3082_ ih.t.timer_max\[10\] _2752_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6208__D net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4306__A _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3984_ _0370_ _1052_ _1058_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5723_ _2518_ mc.cl.next_data\[0\] _2111_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5654_ cu.reg_file.reg_mem\[6\] _2467_ _1739_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__mux2_1
X_4605_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__buf_2
X_5585_ ih.t.timer_max\[19\] _2150_ _2319_ ih.t.timer_max\[3\] _1661_ vssd1 vssd1
+ vccd1 vccd1 _2402_ sky130_fd_sc_hd__a221o_1
XANTENNA__5973__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4536_ cu.reg_file.reg_d\[6\] _1283_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4467_ _1296_ _1523_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__a21o_1
X_4398_ _1441_ _1455_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__nor2_1
X_6206_ clknet_leaf_10_clk net4 net167 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3418_ _0482_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__and2_2
X_6137_ clknet_leaf_10_clk _0171_ net166 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_2
X_3349_ _0405_ _0412_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__or2b_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ clknet_leaf_16_clk _0102_ net174 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5019_ _1998_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output122_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3291__A1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3965__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5370_ _2228_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4543__B2 cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4543__A1 cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4321_ cu.reg_file.reg_c\[3\] _1281_ _1385_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4796__A _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4252_ _0295_ _2914_ _0320_ _1310_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__or4_1
XANTENNA__5404__B _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3203_ _2938_ _2939_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4183_ _0701_ _1252_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3134_ _2745_ _2869_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__or2b_1
X_3065_ ih.t.count\[17\] _2757_ _2801_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout153_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3967_ _0599_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__nor2_1
X_5706_ ih.t.timer_max\[31\] _2151_ _2320_ ih.t.timer_max\[15\] vssd1 vssd1 vccd1
+ vccd1 _2511_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4782__A1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3898_ _0520_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5637_ net98 _2194_ _2450_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5568_ ih.gpio_interrupt_mask\[2\] _2326_ _2385_ _2125_ _2327_ vssd1 vssd1 vccd1
+ vccd1 _2386_ sky130_fd_sc_hd__a221o_1
X_4519_ _1296_ _1572_ _1573_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__a21o_1
X_5499_ _2180_ _2193_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__or2_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5330__A _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output47_A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__A0 cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _1865_ _1866_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3821_ _0895_ _0892_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__or2b_1
XANTENNA__5386__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3752_ cu.reg_file.reg_a\[7\] _0625_ _0628_ cu.reg_file.reg_mem\[15\] _0827_ vssd1
+ vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _0715_ _0711_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5422_ _1306_ _2257_ _2137_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__and3_1
XANTENNA__4516__A1 cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4516__B2 cu.reg_file.reg_sp\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5353_ _2218_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
X_4304_ _2701_ _1354_ _1353_ _1369_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4819__A2 _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5284_ _2177_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4235_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__inv_2
XANTENNA__5492__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4166_ _1175_ _1200_ _1232_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__a31o_1
X_3117_ _2805_ _2807_ _2808_ _2854_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4097_ _0945_ _0946_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__xor2_1
X_3048_ ih.t.count\[23\] _2761_ _2785_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4999_ _1984_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4691__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6023__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3797__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5934__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4020_ _0801_ _0812_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4682__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5564__A_N _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5971_ clknet_leaf_36_clk _0008_ net160 vssd1 vssd1 vccd1 vccd1 cu.alu_f\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4922_ _1909_ _1914_ _1809_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__mux2_1
X_4853_ _0374_ cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3804_ cu.pc.pc_o\[10\] _0740_ _0878_ _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__a211o_1
X_4784_ _1000_ _1786_ cu.id.is_halted vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3735_ _0805_ _0808_ _0810_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__or3_2
X_5405_ _0619_ net132 _2248_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__mux2_1
X_3666_ cu.reg_file.reg_d\[0\] _0488_ _0741_ cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1
+ vccd1 _0742_ sky130_fd_sc_hd__a22o_1
X_3597_ _0374_ _0672_ _0294_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__mux2_1
X_5336_ _2209_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__clkbuf_1
X_5267_ ih.t.timer_max\[31\] _2167_ _2153_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__mux2_1
X_4218_ _0295_ _0469_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__nor2_4
XANTENNA__4673__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5198_ mc.cc.count\[3\] _1652_ _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__o21ba_1
X_4149_ _0941_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__nand2_1
XANTENNA__4976__A1 cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5153__A1 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4664__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3467__A1 cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3957__B _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5392__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4195__A2 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3520_ _0594_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__nand2_1
X_3451_ _0521_ _0524_ _0525_ _0526_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__and4b_1
XANTENNA__5144__A1 _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3382_ net148 _0454_ _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__a21oi_4
X_6170_ clknet_leaf_40_clk _0204_ net164 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5121_ _1622_ _0617_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__mux2_1
X_5052_ _0618_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4003_ _0764_ _1064_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5954_ cu.id.imm_i\[8\] _2350_ _2686_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__mux2_1
XANTENNA__5080__A0 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5885_ _2649_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ cu.id.cb_opcode_x\[1\] cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__and2_1
X_4836_ _1828_ _1835_ _1809_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4767_ _1483_ _1632_ _1643_ _1771_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__o311a_1
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5574__S _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4698_ net230 _1714_ _1687_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__o21ai_1
X_3718_ _0664_ _0682_ _0793_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3649_ cu.reg_file.reg_sp\[7\] _0413_ _0419_ cu.reg_file.reg_h\[7\] _0724_ vssd1
+ vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__a221o_1
XANTENNA__5135__A1 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5319_ _2199_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_1
Xhold23 ih.t.count\[4\] vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlygate4sd3_1
X_6299_ clknet_leaf_42_clk _0281_ net153 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold12 cu.alu_f\[3\] vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 ih.t.count\[27\] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__A1 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4219__A _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2962__A _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5610__A2 _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3621__B2 cu.reg_file.reg_h\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3621__A1 cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4889__A cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 keypad_input[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5126__A1 _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4033__A2_N _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5062__A0 cu.reg_file.reg_c\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5601__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3612__A1 cu.reg_file.reg_h\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ net75 _1648_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3612__B2 cu.reg_file.reg_a\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4621_ _1647_ _1663_ _2706_ vssd1 vssd1 vccd1 vccd1 mc.rw.next_state\[1\] sky130_fd_sc_hd__a21o_1
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5394__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ _1382_ _1602_ _1603_ _1605_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__a31o_2
X_4483_ _1296_ _1538_ _1539_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__a21o_1
X_3503_ cu.reg_file.reg_sp\[2\] _0413_ _0415_ cu.reg_file.reg_d\[2\] _0578_ vssd1
+ vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__a221o_1
XANTENNA__5117__A1 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6222_ clknet_leaf_15_clk net216 net175 vssd1 vssd1 vccd1 vccd1 ih.t.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3434_ _0447_ net143 vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__xnor2_2
X_6153_ clknet_leaf_15_clk _0187_ net177 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ cu.reg_file.reg_l\[0\] _0422_ _0431_ _0434_ _0440_ vssd1 vssd1 vccd1 vccd1
+ _0441_ sky130_fd_sc_hd__a2111o_1
X_6084_ clknet_leaf_19_clk _0118_ net180 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5104_ _2057_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
X_3296_ cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ cu.reg_file.reg_b\[2\] _2010_ _2006_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5937_ _2677_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3603__A1 cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3603__B2 cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5868_ _2640_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5356__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4819_ _0343_ _1299_ _1818_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__a21oi_1
X_5799_ cu.reg_file.reg_sp\[8\] _2535_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 memory_address_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 memory_address_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 memory_data_out[6] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[0] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 ss0[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__4619__A0 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4891__B cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__A0 cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4555__C1 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5942__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5504__D1 _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4858__A0 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4248__B_N _1311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3150_ _2883_ _2884_ _2885_ _2886_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__and4_2
X_3081_ ih.t.count\[11\] _2753_ _2817_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__and3_1
XANTENNA__5283__A0 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5586__A1 _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3983_ cu.alu_f\[1\] _1023_ _1056_ _1057_ _1027_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o221a_1
X_5722_ _2869_ _2870_ _2873_ net205 vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__a22o_1
XANTENNA__3597__A0 _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5653_ _2463_ _2464_ _2466_ _1641_ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__o22a_4
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5584_ _1400_ _2400_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__and2b_1
X_4604_ _1485_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4535_ cu.reg_file.reg_sp\[14\] _1286_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4466_ cu.id.imm_i\[10\] _1294_ _1297_ _1521_ _1489_ vssd1 vssd1 vccd1 vccd1 _1524_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4397_ _2701_ _1441_ _1353_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__a21o_1
XANTENNA__5510__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6205_ clknet_leaf_9_clk net3 net169 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3417_ _0458_ _0486_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nor2_1
XANTENNA__4695__C _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6136_ clknet_leaf_9_clk _0170_ net165 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3348_ _0408_ _0407_ _0293_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__a21o_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6067_ clknet_leaf_19_clk _0101_ net180 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3279_ _0340_ _0341_ _0343_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5299__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5018_ cu.reg_file.reg_a\[6\] _1997_ _1985_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5577__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5501__A1 ih.t.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4304__A2 _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3815__A1 cu.reg_file.reg_a\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output115_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5017__A0 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5002__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4240__A1 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4018__A1_N _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5740__A1 _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4320_ cu.reg_file.reg_e\[3\] _1283_ _1285_ cu.reg_file.reg_l\[3\] _1384_ vssd1 vssd1
+ vccd1 vccd1 _1385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4251_ _1318_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__inv_2
X_3202_ _2899_ cu.id.opcode\[1\] _2875_ _2876_ vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3205__B _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4182_ _1248_ _1251_ _0588_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__mux2_1
X_3133_ _2870_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__inv_2
XANTENNA__4059__B2 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3064_ _2757_ _2801_ ih.t.count\[17\] vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3806__A1 cu.id.imm_i\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5008__A0 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5559__B2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ _0447_ _0588_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5705_ net7 _1650_ _2488_ _2510_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__a31o_1
XANTENNA__4782__A2 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5636_ net130 _2236_ _2247_ net138 vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__a22o_1
X_3897_ _2885_ _2886_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5567_ mc.cl.next_data\[2\] _2359_ net237 _2384_ vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5498_ ih.t.timer_max\[0\] _2314_ _2317_ _1400_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__o2bb2a_1
X_4518_ cu.id.imm_i\[13\] _1294_ _1297_ cu.pc.pc_o\[13\] _1488_ vssd1 vssd1 vccd1
+ vccd1 _1573_ sky130_fd_sc_hd__a221o_1
X_4449_ cu.reg_file.reg_sp\[9\] _0993_ _1344_ cu.id.imm_i\[9\] _1324_ vssd1 vssd1
+ vccd1 vccd1 _1508_ sky130_fd_sc_hd__a221o_1
X_6119_ clknet_leaf_10_clk _0153_ net167 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4470__A1 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2970__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4222__A1 cu.reg_file.reg_c\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5722__A1 _2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5486__A0 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5240__B _1372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3976__A _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _0892_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__or2b_1
X_3751_ cu.pc.pc_o\[15\] _0740_ _0825_ _0826_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3682_ _0511_ _0712_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5421_ _1329_ _1372_ _1369_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__and3_1
XANTENNA__4516__A2 _1282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4600__A _1632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5352_ _1075_ net110 _2215_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__mux2_1
X_4303_ _1368_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5283_ net82 _1193_ _2170_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4234_ _1300_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4165_ _0387_ _1234_ _0824_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__a21oi_1
X_3116_ _2810_ _2811_ _2853_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__or3_1
XANTENNA__5431__A _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4096_ _0546_ _0733_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__xor2_1
X_3047_ ih.t.timer_max\[22\] _2760_ ih.t.timer_max\[23\] vssd1 vssd1 vccd1 vccd1 _2785_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4998_ _2951_ _0367_ _0352_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3949_ _1023_ _1024_ alu.Cin _1021_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4507__A2 _1545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5619_ net105 _2205_ _2433_ _1401_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__a22o_1
XANTENNA__5704__B2 _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4140__B1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5640__B1 _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5950__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4434__A1 cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4434__B2 cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5970_ clknet_leaf_36_clk _0007_ net160 vssd1 vssd1 vccd1 vccd1 alu.Cin sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4921_ _1912_ _1913_ _1798_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__mux2_1
X_4852_ cu.pc.pc_o\[4\] _1838_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3803_ cu.reg_file.reg_b\[2\] _0743_ _0624_ cu.reg_file.reg_sp\[10\] vssd1 vssd1
+ vccd1 vccd1 _0879_ sky130_fd_sc_hd__a22o_1
XANTENNA__5934__A1 _2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4783_ _0986_ _0989_ _0994_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3734_ _0763_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3665_ _0464_ _0482_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__and2_2
X_5404_ net141 _2247_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__nand2_8
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3596_ ih.interrupt_source\[3\] ih.interrupt_source\[2\] vssd1 vssd1 vccd1 vccd1
+ _0672_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5335_ _1075_ net102 _2206_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5266_ _1110_ _1263_ _1666_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4217_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__buf_2
X_5197_ mc.cc.count\[0\] _2708_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__or2_2
X_4148_ _0939_ _0940_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__or2_1
X_4079_ _1060_ _0600_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4189__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5684__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6244__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5916__A1 _1484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3450_ _2925_ _2901_ _2912_ _2897_ _2935_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__o221a_1
X_3381_ cu.id.starting_int_service _0382_ _0456_ _2896_ vssd1 vssd1 vccd1 vccd1 _0457_
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ _2065_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__buf_4
X_5051_ _2021_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4002_ _0761_ _0764_ _0772_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__and3b_1
XANTENNA__5974__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4407__A1 cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4407__B2 cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5953_ _2685_ vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5080__A1 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5884_ _1187_ ih.t.timer_max\[3\] _2645_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__mux2_1
X_4904_ _2920_ cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5907__A1 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4835_ _1833_ _1834_ _1799_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__mux2_1
X_4766_ _1303_ _1772_ _1773_ _1765_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3717_ _0652_ _0663_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__and2b_1
X_4697_ ih.t.count\[21\] _1714_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3648_ cu.reg_file.reg_d\[7\] _0415_ _0432_ cu.reg_file.reg_b\[7\] vssd1 vssd1 vccd1
+ vccd1 _0724_ sky130_fd_sc_hd__a22o_1
X_3579_ cu.id.cb_opcode_y\[2\] _0654_ _0294_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__mux2_1
X_5318_ _1188_ net95 _2195_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__mux2_1
Xhold13 mc.cc.count\[0\] vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlygate4sd3_1
X_6298_ clknet_leaf_42_clk _0280_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_y\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold24 ih.t.count\[28\] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 ih.t.count\[24\] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ ih.t.timer_max\[25\] _2155_ _2153_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__mux2_1
XANTENNA__4934__S _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2962__B _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5005__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5062__A1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3612__A2 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4620_ _1651_ _1662_ _2699_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4573__B1 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4551_ _1402_ _1598_ _1604_ _1371_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4482_ cu.id.imm_i\[11\] _1294_ _1297_ cu.pc.pc_o\[11\] _1489_ vssd1 vssd1 vccd1
+ vccd1 _1539_ sky130_fd_sc_hd__a221o_1
X_3502_ cu.reg_file.reg_b\[2\] _0432_ _0433_ cu.reg_file.reg_a\[2\] vssd1 vssd1 vccd1
+ vccd1 _0578_ sky130_fd_sc_hd__a22o_1
X_6221_ clknet_leaf_14_clk ih.t.next_count\[9\] net175 vssd1 vssd1 vccd1 vccd1 ih.t.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3433_ _0491_ _0497_ _0506_ _0508_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__o31ai_2
X_6152_ clknet_leaf_12_clk _0186_ net177 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5103_ cu.reg_file.reg_e\[0\] _2022_ _2056_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__mux2_1
X_3364_ _0293_ _0362_ _0438_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or4_4
X_6083_ clknet_leaf_23_clk _0117_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _2950_ _0361_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__nand2_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _1074_ _1226_ _2002_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5936_ _0343_ _2350_ _2666_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__mux2_1
X_5867_ _2159_ ih.t.timer_max\[11\] _2636_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__mux2_1
X_4818_ _0343_ _1299_ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5798_ _2582_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4749_ _1739_ _1757_ _1483_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__a21oi_1
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 memory_address_out[10] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 memory_data_out[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 memory_address_out[6] sky130_fd_sc_hd__clkbuf_4
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__3134__A _2745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2973__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3358__A1 cu.reg_file.reg_b\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3358__B2 cu.reg_file.reg_a\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3309__A _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5504__C1 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5524__A _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3080_ _2753_ _2817_ ih.t.count\[11\] vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5283__A1 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3982_ _0298_ _1001_ _1002_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__o21ai_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4794__A0 _0617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5721_ net1 net198 _2872_ _2870_ _2521_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4603__A _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5652_ _1649_ _2465_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__and2_1
X_5583_ ih.t.timer_max\[11\] _2193_ _2314_ ih.t.timer_max\[3\] _2399_ vssd1 vssd1
+ vccd1 vccd1 _2400_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4603_ _1646_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__buf_2
XFILLER_0_60_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4534_ _1580_ _1582_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5434__A _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4465_ cu.reg_file.reg_b\[2\] net238 _1284_ cu.reg_file.reg_h\[2\] _1522_ vssd1 vssd1
+ vccd1 vccd1 _1523_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5510__A2 _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4396_ _1419_ _1436_ _1456_ _1445_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__nand4_1
X_6204_ clknet_leaf_8_clk net17 net169 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3416_ net147 _0473_ net146 _0463_ _0458_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__o2111a_4
X_6135_ clknet_leaf_9_clk _0169_ net165 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_4
XANTENNA__3521__A1 _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3347_ _0417_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ clknet_leaf_26_clk _0100_ net195 vssd1 vssd1 vccd1 vccd1 mc.cc.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _2883_ _2936_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__or2_1
X_5017_ _1193_ _1624_ _0368_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__mux2_1
XANTENNA__4482__C1 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5577__A2 _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5919_ cu.ir.idx\[0\] cu.ir.idx\[1\] vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__nor2_4
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3760__A1 cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5017__A1 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output108_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3751__A1 cu.pc.pc_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4250_ _2893_ _2901_ _2923_ _2936_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__or4b_4
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4700__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3201_ cu.id.alu_opcode\[0\] _2894_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__or2b_1
X_4181_ _1249_ _1250_ _0599_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__mux2_1
XANTENNA__3503__A1 cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3132_ ih.ih.int_f.prev_data ih.ih.int_f.data_in ih.input_handler_enable vssd1 vssd1
+ vccd1 vccd1 _2870_ sky130_fd_sc_hd__and3b_4
X_3063_ ih.t.timer_max\[16\] _2756_ ih.t.timer_max\[17\] vssd1 vssd1 vccd1 vccd1 _2801_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5008__A1 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5559__A2 _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3824__A2_N _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _0710_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5704_ _2509_ _1643_ cu.reg_file.reg_mem\[14\] _1646_ vssd1 vssd1 vccd1 vccd1 _2510_
+ sky130_fd_sc_hd__a2bb2o_1
X_3896_ _2935_ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5635_ _2449_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5566_ _1666_ _2382_ _2383_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5497_ _2315_ _2316_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__nor2_1
X_4517_ cu.reg_file.reg_b\[5\] net144 _1284_ cu.reg_file.reg_h\[5\] _1571_ vssd1 vssd1
+ vccd1 vccd1 _1572_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3742__A1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4448_ cu.reg_file.reg_h\[1\] _1316_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__and2_1
XANTENNA__5495__A1 ih.t.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5495__B2 ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4379_ _1404_ _1417_ _1434_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__a21bo_1
X_6118_ clknet_leaf_11_clk _0152_ net167 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ clknet_leaf_6_clk _0087_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4470__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5722__A2 _2870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5486__A1 _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4997__A0 _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5948__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3750_ cu.reg_file.reg_b\[7\] _0743_ _0624_ cu.reg_file.reg_sp\[15\] vssd1 vssd1
+ vccd1 vccd1 _0826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3681_ _0664_ _0756_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__xnor2_1
X_5420_ _2256_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5351_ _2217_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4600__B _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5282_ _2176_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
X_4302_ _1306_ _1362_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4233_ cu.id.state\[1\] vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _1233_ _0371_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__nor2_1
X_3115_ _2813_ _2815_ _2816_ _2852_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__or4_1
XANTENNA__5431__B _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4095_ _0566_ _1110_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__xnor2_1
X_3046_ _2762_ _2782_ ih.t.count\[24\] vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4997_ _0618_ _1622_ _0368_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__mux2_1
X_3948_ _0572_ _1020_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5165__A0 cu.reg_file.reg_l\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4998__A _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3879_ _0771_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__or2b_1
X_5618_ net89 _1330_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4510__B _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5549_ net69 _1649_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__a31o_1
XANTENNA__4912__A0 cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5640__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5640__B2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4903__A0 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5008__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5631__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4434__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5631__B2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4920_ _1623_ _1909_ _1794_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__mux2_1
X_4851_ _1849_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3802_ cu.reg_file.reg_d\[2\] _0488_ _0741_ cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1
+ vccd1 _0878_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4782_ _0350_ _2948_ _1782_ net204 vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3733_ _0759_ _0783_ _0784_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3664_ _0501_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5698__B2 ih.t.timer_max\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__A1 ih.t.timer_max\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5403_ _2246_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3595_ _0576_ _0665_ _0667_ _0670_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__o2bb2a_1
X_5334_ _2208_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5265_ _2166_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4122__B2 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4216_ _1279_ _1275_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__nor2_4
X_5196_ _2117_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
X_4147_ _0951_ _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__nor2_1
XANTENNA__5622__A1 ih.t.timer_max\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4078_ _0558_ _0663_ _0822_ _0694_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a22o_1
X_3029_ ih.t.count\[31\] _2766_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5386__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5138__A0 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5689__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4361__A1 _1415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2976__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5861__A1 ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3321__C1 _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6284__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5377__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5916__A2 _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5129__A0 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3380_ _0300_ _2911_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5301__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5050_ cu.reg_file.reg_b\[7\] _2020_ _2006_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4606__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ _2663_ cu.ir.idx\[1\] vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__and2_1
X_4903_ _1622_ _1896_ _1795_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__mux2_1
XANTENNA__3615__B1 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5883_ _2648_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4834_ _1073_ _1828_ _1795_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4765_ _1747_ _1763_ _1761_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__a21boi_1
XANTENNA__5437__A _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3716_ _0733_ _0790_ _0729_ _0791_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__o2bb2a_1
X_4696_ _1716_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[20\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3647_ _0293_ _0372_ _0634_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__or3_1
X_3578_ ih.interrupt_source\[3\] ih.interrupt_source\[1\] vssd1 vssd1 vccd1 vccd1
+ _0654_ sky130_fd_sc_hd__or2_1
X_5317_ _2198_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_1
Xhold14 _0097_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dlygate4sd3_1
X_6297_ clknet_leaf_41_clk _0279_ net159 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_z\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold25 ih.t.count\[25\] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 ih.ih.ih.prev_data\[11\] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _1050_ _1623_ _1667_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__mux2_1
X_5179_ mc.cl.next_data\[12\] net22 mc.count vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5347__A _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output138_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5021__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5956__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4145__B _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4573__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4161__A _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4573__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550_ _1585_ _1598_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4481_ cu.reg_file.reg_b\[3\] net144 _1284_ cu.reg_file.reg_h\[3\] _1537_ vssd1 vssd1
+ vccd1 vccd1 _1538_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3501_ cu.reg_file.reg_c\[2\] _0427_ _0430_ cu.reg_file.reg_e\[2\] vssd1 vssd1 vccd1
+ vccd1 _0577_ sky130_fd_sc_hd__a22o_1
X_6220_ clknet_leaf_14_clk ih.t.next_count\[8\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3432_ _0343_ _2949_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4325__A1 cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4325__B2 cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6151_ clknet_leaf_11_clk _0185_ net168 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ net151 _2914_ _0318_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__or3_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5102_ _2035_ _2055_ _2951_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__o21a_4
X_6082_ clknet_leaf_23_clk _0116_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__buf_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _2009_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout169_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4336__A _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5935_ _2676_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
X_5866_ _2639_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
X_4817_ _0340_ cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5797_ cu.reg_file.reg_sp\[7\] _2581_ _2539_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__mux2_1
X_4748_ _0371_ _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__nand2_1
X_4679_ ih.t.count\[15\] _1702_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 memory_address_out[11] sky130_fd_sc_hd__buf_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 memory_address_out[7] sky130_fd_sc_hd__buf_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 memory_wr sky130_fd_sc_hd__clkbuf_4
XANTENNA__4945__S _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3625__A1_N _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3000__A_N net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__A _1309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4555__B2 cu.pc.pc_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4555__A1 cu.id.imm_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3309__B _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3818__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4156__A _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3981_ _1023_ _1054_ _1055_ cu.alu_f\[1\] vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__o2bb2a_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5720_ net1 ih.interrupt_source\[3\] vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_42_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5651_ net14 _2345_ _2369_ net7 vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__a22o_1
X_5582_ ih.t.timer_max\[27\] _2146_ _2204_ ih.t.timer_max\[19\] vssd1 vssd1 vccd1
+ vccd1 _2399_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ _1645_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4533_ _1353_ _1579_ _1583_ _1584_ _1587_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__a221o_1
XFILLER_0_13_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5434__B _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6203_ clknet_leaf_7_clk net16 net172 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4464_ cu.reg_file.reg_d\[2\] _1282_ _1286_ cu.reg_file.reg_sp\[10\] vssd1 vssd1
+ vccd1 vccd1 _1522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4395_ _1419_ _1436_ _1445_ _1456_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__a31o_1
X_3415_ cu.reg_file.reg_c\[0\] _0485_ _0489_ cu.reg_file.reg_e\[0\] _0490_ vssd1 vssd1
+ vccd1 vccd1 _0491_ sky130_fd_sc_hd__a221o_1
X_6134_ clknet_leaf_10_clk _0168_ net166 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3346_ _0414_ _0421_ _0417_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__a21oi_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ clknet_leaf_26_clk net224 net194 vssd1 vssd1 vccd1 vccd1 mc.cc.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6316__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _2892_ _0324_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5016_ _1996_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5918_ net204 _2667_ _1781_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5849_ _2625_ _2626_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4537__A1 cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4537__B2 cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3760__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2984__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output82_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3751__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3200_ _2936_ _2901_ _2898_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__or3_2
X_4180_ _0694_ _1040_ _1060_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__mux2_1
X_3131_ _2768_ _2864_ _2867_ _2868_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__or4b_4
X_3062_ ih.t.count\[18\] _2758_ _2798_ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4464__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3964_ _0570_ _0712_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5703_ mc.cl.next_data\[14\] _2359_ _2490_ _2508_ vssd1 vssd1 vccd1 vccd1 _2509_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3895_ _2893_ _2896_ _2912_ _2923_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__o22a_1
XANTENNA__4519__A1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5634_ cu.reg_file.reg_mem\[5\] _2448_ _2351_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5565_ ih.t.timer_max\[18\] _2150_ _2319_ ih.t.timer_max\[2\] _1661_ vssd1 vssd1
+ vccd1 vccd1 _2383_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5496_ ih.t.timer_max\[24\] _2146_ _2204_ ih.t.timer_max\[16\] vssd1 vssd1 vccd1
+ vccd1 _2316_ sky130_fd_sc_hd__a22o_1
X_4516_ cu.reg_file.reg_d\[5\] _1282_ _1286_ cu.reg_file.reg_sp\[13\] vssd1 vssd1
+ vccd1 vccd1 _1571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4447_ cu.id.imm_i\[9\] _1295_ _1298_ cu.pc.pc_o\[9\] _1305_ vssd1 vssd1 vccd1 vccd1
+ _1506_ sky130_fd_sc_hd__a221o_1
X_6117_ clknet_leaf_13_clk _0151_ net173 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
X_4378_ _1404_ _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__nand2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5180__A _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ _0403_ _0404_ cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__a21o_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ clknet_leaf_6_clk _0086_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3430__A1 alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3430__B2 cu.reg_file.reg_a\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2979__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4446__B1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output120_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4997__A1 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4137__C _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4749__A1 _1739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5946__A0 _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3421__A1 cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5964__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3680_ _0718_ _0755_ _0720_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5350_ _1052_ net109 _2215_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5281_ net81 _1191_ _2170_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__mux2_1
X_4301_ cu.reg_file.reg_c\[2\] _1313_ _1363_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_
+ sky130_fd_sc_hd__a211o_1
X_4232_ cu.id.state\[0\] vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__buf_2
XANTENNA__3488__A1 cu.reg_file.reg_a\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4163_ _2920_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__buf_4
X_3114_ _2818_ _2819_ _2851_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__or3_1
X_4094_ _1090_ _1164_ _1166_ _0611_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__o221a_1
X_3045_ ih.t.count\[24\] _2762_ _2782_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4996_ _1982_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3947_ _1003_ _1011_ _1020_ _1022_ _2948_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__o41a_2
XFILLER_0_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3878_ _0898_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__xnor2_1
X_5617_ net97 _2194_ _2431_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__a21o_1
XANTENNA__5165__A1 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5548_ _2169_ _2358_ _2366_ _2136_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__o211a_1
XANTENNA__4510__C _1545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5479_ _2301_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5625__C1 _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5640__A2 _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3651__B2 cu.reg_file.reg_a\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5928__A0 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4254__A _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3333__A cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output45_A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__A0 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ cu.pc.pc_o\[3\] _1848_ _1815_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4164__A _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3801_ _0875_ _0876_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__or2_1
X_4781_ net200 _1785_ net204 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__o21ba_1
X_3732_ _0806_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3663_ _0738_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5402_ _1369_ _2148_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5333_ _1052_ net101 _2206_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3594_ cu.reg_file.reg_l\[4\] _0422_ _0668_ _0669_ _0576_ vssd1 vssd1 vccd1 vccd1
+ _0670_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5264_ ih.t.timer_max\[30\] _2165_ _2153_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4122__A2 _1186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5195_ cu.reg_file.reg_sp\[0\] _2085_ _2116_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__mux2_1
X_4215_ _1282_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__buf_2
X_4146_ _0917_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5083__A0 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4077_ _0570_ _0684_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3028_ ih.t.timer_max\[30\] _2765_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3633__A1 _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5386__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4979_ _1948_ _1956_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__and2b_1
XANTENNA__3397__B1 _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5138__A1 _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5689__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3321__B1 cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5074__A0 _0617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4821__A0 _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3624__A1 cu.reg_file.reg_l\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5377__A1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5916__A3 _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5808__A cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5129__A1 _1073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5301__A1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5951_ _2684_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3615__A1 cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4902_ _1894_ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3615__B2 cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5882_ _1074_ ih.t.timer_max\[2\] _2645_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4833_ _1831_ _1832_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5718__A _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4764_ _1268_ _1747_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5437__B _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ _0566_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4695_ _1714_ _1715_ _1672_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3646_ _0652_ _0663_ _0685_ _0718_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a221o_1
XANTENNA__5453__A _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5976__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3577_ _0507_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__buf_8
X_5316_ _1075_ net94 _2195_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6296_ clknet_leaf_0_clk _0278_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_z\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5247_ _2154_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__clkbuf_1
Xhold26 mc.cc.count\[3\] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 cu.ir.idx\[1\] vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 cu.alu_f\[4\] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _2104_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
X_4129_ _0959_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__or2_1
XANTENNA__5056__A0 cu.reg_file.reg_c\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4031__B2 _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5295__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4098__A1 _0916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4098__B2 _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5047__A0 cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4270__B2 cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4270__A1 cu.reg_file.reg_a\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4558__C1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4573__A2 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3500_ _0440_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4161__B _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4480_ cu.reg_file.reg_d\[3\] _1282_ _1286_ cu.reg_file.reg_sp\[11\] vssd1 vssd1
+ vccd1 vccd1 _1537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3431_ _0504_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__inv_2
XANTENNA__4325__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6150_ clknet_leaf_12_clk _0184_ net174 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3362_ _2880_ _0437_ _0323_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _1791_ _0366_ _2037_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__and3_1
X_6081_ clknet_leaf_23_clk _0115_ net193 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3293_ _2951_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__and2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5032_ cu.reg_file.reg_b\[1\] _2008_ _2006_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__mux2_1
XANTENNA__5038__A0 cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5934_ _2876_ _2486_ _2668_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__mux2_1
X_5865_ _2157_ ih.t.timer_max\[10\] _2636_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4816_ _1299_ cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5796_ _1110_ _2580_ _2545_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__mux2_1
XANTENNA__5882__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4747_ _1754_ _1747_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4678_ _1704_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5513__B2 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5513__A1 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3629_ cu.reg_file.reg_h\[2\] _0495_ _0499_ cu.reg_file.reg_a\[2\] vssd1 vssd1 vccd1
+ vccd1 _0705_ sky130_fd_sc_hd__a22o_1
XANTENNA__5183__A _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 memory_address_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 memory_address_out[8] sky130_fd_sc_hd__clkbuf_4
X_6279_ clknet_leaf_16_clk _0261_ net178 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5277__A0 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5029__A0 cu.reg_file.reg_b\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__B _1311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4961__S _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3763__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5504__A1 _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3818__A1 cu.reg_file.reg_b\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3818__B2 cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3341__A _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5032__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3980_ _0395_ _1019_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__nor2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3995__B _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5650_ net74 _1648_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__a31o_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _1364_ _1489_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5581_ net79 _1633_ _2394_ _2397_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__o22a_1
X_4532_ _1585_ _1586_ _1356_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4900__A cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3754__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4463_ cu.pc.pc_o\[10\] vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6202_ clknet_leaf_7_clk net15 net172 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3414_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[0\] vssd1 vssd1 vccd1 vccd1 _0490_
+ sky130_fd_sc_hd__o211a_1
X_4394_ _1396_ _1455_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6133_ clknet_leaf_13_clk _0167_ net173 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
X_3345_ _0409_ _0407_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ clknet_leaf_26_clk _0098_ net194 vssd1 vssd1 vccd1 vccd1 mc.cc.count\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _0348_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__nor2_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ cu.reg_file.reg_a\[5\] _1995_ _1985_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout181_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4482__B2 cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4482__A1 cu.id.imm_i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5917_ _1780_ _2532_ net203 vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _2618_ _2621_ _2619_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__a21boi_2
X_5779_ _2564_ _2565_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5991__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3161__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6097__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3100__S ih.t.timer_max\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5816__A cu.reg_file.reg_sp\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5489__B1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3130_ ih.t.count\[30\] _2866_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__nand2_1
X_3061_ _2758_ _2798_ ih.t.count\[18\] vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4464__B2 cu.reg_file.reg_sp\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4167__A _0617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5413__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5964__A1 _2448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__A2 _1632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3963_ _0918_ _1029_ _1034_ _1037_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__o22a_1
X_5702_ ih.t.timer_max\[30\] _2151_ _2320_ ih.t.timer_max\[14\] vssd1 vssd1 vccd1
+ vccd1 _2508_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3894_ _0967_ _0969_ _0328_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__a21oi_1
X_5633_ _2444_ _2445_ _2447_ _1641_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__o22a_4
X_5564_ _1400_ _2381_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4515_ _1382_ _1564_ _1565_ _1570_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__a31o_1
X_5495_ ih.t.enable _2257_ _2192_ ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1 _2315_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4446_ _1503_ _1504_ _1296_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__o21a_1
X_4377_ _1415_ _1434_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__nor2_1
XANTENNA__4152__B1 _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6116_ clknet_leaf_24_clk _0150_ net192 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3328_ _2925_ _2890_ _2932_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__or3_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ clknet_leaf_7_clk _0085_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3259_ _0321_ _0322_ _0328_ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__nor4_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5400__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output113_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5946__A1 _2448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3421__A2 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5280_ _2175_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ cu.pc.pc_o\[2\] _1322_ _1317_ cu.reg_file.reg_l\[2\] _1365_ vssd1 vssd1 vccd1
+ vccd1 _1366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4231_ cu.pc.pc_o\[0\] vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5882__A0 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4162_ _1209_ _1213_ _1222_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__nor4_1
X_3113_ _2821_ _2823_ _2824_ _2850_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__or4_1
X_4093_ _1090_ _1164_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__nand2_1
X_3044_ ih.t.timer_max\[24\] _2761_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4625__A _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4995_ cu.pc.pc_o\[15\] _1981_ _1814_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3946_ _1012_ _0996_ _1016_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3877_ _0737_ _0752_ _0899_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5616_ net129 _2236_ _2247_ net137 vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5890__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5547_ ih.gpio_interrupt_mask\[1\] _2326_ _2365_ _2125_ _2327_ vssd1 vssd1 vccd1
+ vccd1 _2366_ sky130_fd_sc_hd__a221o_1
X_5478_ net65 _0618_ _2300_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__mux2_1
X_4429_ _1488_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__buf_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5130__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4535__A cu.reg_file.reg_sp\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5928__A1 _2429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5305__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6041__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5616__B1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__A1 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3627__C1 cu.reg_file.reg_l\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5040__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4780_ _1768_ _1784_ _0350_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__o21a_1
X_3800_ _0874_ _0871_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3731_ _0572_ _0510_ _0712_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _2950_ _2913_ _0536_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5401_ _2245_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
X_3593_ cu.reg_file.reg_mem\[4\] _0418_ _0433_ cu.reg_file.reg_a\[4\] vssd1 vssd1
+ vccd1 vccd1 _0669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5332_ _2207_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5263_ _1126_ _1624_ _1666_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__mux2_1
XANTENNA__4339__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4214_ _1279_ _1275_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__nor2b_4
X_5194_ _2115_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__inv_2
X_4145_ _1214_ _0779_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__or2_1
XANTENNA__5083__A1 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4076_ _0918_ _0766_ _1149_ _0517_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3027_ ih.t.timer_max\[28\] ih.t.timer_max\[29\] _2764_ vssd1 vssd1 vccd1 vccd1 _2765_
+ sky130_fd_sc_hd__or3_1
XANTENNA__3633__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _1233_ cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__xor2_1
XANTENNA__5186__A _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3929_ _0976_ _0980_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3434__A _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5074__A1 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5808__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5824__A cu.reg_file.reg_sp\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5035__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5837__A0 cu.reg_file.reg_sp\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5950_ _1233_ _2486_ _2666_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__mux2_1
X_4901_ cu.pc.pc_o\[7\] _1872_ cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4812__A1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4812__B2 _1484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5881_ _2647_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4832_ _0340_ cu.pc.pc_o\[1\] _1819_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4763_ _1739_ _1770_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__nand2_1
XANTENNA__4576__B1 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4694_ ih.t.count\[18\] ih.t.count\[19\] _1708_ ih.t.count\[20\] vssd1 vssd1 vccd1
+ vccd1 _1715_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3714_ _0643_ _0632_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5990__SET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3645_ _0719_ _0720_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3576_ _0576_ _0646_ _0648_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o2bb2a_4
X_5315_ _2197_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
X_6295_ clknet_leaf_0_clk _0277_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_z\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3551__B2 cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3551__A1 cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5828__A0 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5246_ ih.t.timer_max\[24\] _2144_ _2153_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold16 ih.t.count\[19\] vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 ih.t.count\[15\] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 _0099_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _1647_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__and2_1
XANTENNA__5056__A1 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4128_ _0949_ _0958_ _0779_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__a21o_1
XANTENNA__3701__B _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4059_ _0917_ _0757_ _0804_ _0776_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4813__A _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5295__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4558__B1 _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3781__A1 cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4161__C _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3781__B2 cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3430_ alu.Cin _0498_ _0499_ cu.reg_file.reg_a\[0\] _0505_ vssd1 vssd1 vccd1 vccd1
+ _0506_ sky130_fd_sc_hd__a221o_1
X_3361_ _0308_ _0315_ _0435_ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__and4bb_2
XANTENNA__4730__B1 _1644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3074__A ih.t.timer_max\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6080_ clknet_leaf_23_clk _0114_ net192 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5100_ _2054_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _2953_ _0339_ _0352_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__o211a_4
X_5031_ _1051_ _1623_ _2002_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__mux2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5933_ _2675_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__clkbuf_1
X_5864_ _2638_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
X_4815_ _1816_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5795_ _2578_ _2579_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4746_ _1483_ _1748_ _1754_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3772__A1 cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4677_ _1702_ _1703_ _1672_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__and3b_1
XANTENNA__5464__A _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3628_ cu.reg_file.reg_c\[2\] _0485_ _0489_ cu.reg_file.reg_e\[2\] _0703_ vssd1 vssd1
+ vccd1 vccd1 _0704_ sky130_fd_sc_hd__a221o_1
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 memory_address_out[13] sky130_fd_sc_hd__buf_2
X_3559_ _0295_ _2921_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__or3_1
X_6278_ clknet_leaf_16_clk _0260_ net178 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5498__A1_N ih.t.timer_max\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5277__A1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5229_ _1306_ _2137_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__and2_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3763__A1 cu.reg_file.reg_sp\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3763__B2 cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3515__A1 cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3515__B2 cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3818__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4437__B _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3341__B _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4600_ _1632_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__nor2_4
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5580_ net111 _2147_ _2225_ net119 _2396_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__a221o_1
X_4531_ _1567_ _1579_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__nand2_1
XANTENNA__4900__B cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3754__B2 cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3754__A1 cu.reg_file.reg_sp\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4462_ _1513_ _1514_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__nand2_1
X_6201_ clknet_leaf_12_clk net14 net169 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3506__A1 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3413_ _0480_ _0487_ _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__a21o_2
XFILLER_0_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4393_ _1449_ _1450_ _1454_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__o21a_2
XFILLER_0_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6132_ clknet_leaf_27_clk _0166_ net195 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_4
X_3344_ cu.reg_file.reg_mem\[0\] _0418_ _0419_ cu.reg_file.reg_h\[0\] vssd1 vssd1
+ vccd1 vccd1 _0420_ sky130_fd_sc_hd__a22o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4628__A ih.t.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6063_ clknet_leaf_25_clk net211 net194 vssd1 vssd1 vccd1 vccd1 mc.cc.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _0299_ _2953_ _0349_ _2914_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__a221o_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _1191_ _1209_ _0368_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5916_ _1484_ _2351_ _2666_ _2665_ net234 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__a32o_1
XANTENNA__5195__A0 cu.reg_file.reg_sp\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5847_ cu.reg_file.reg_sp\[14\] _1287_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5778_ _2550_ _2551_ _2557_ _2556_ _2549_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__a311o_1
XFILLER_0_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4729_ _1738_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[31\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5498__B2 _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5133__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4972__S _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4704__C _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6066__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4933__A0 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5816__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5489__B2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5489__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5832__A cu.reg_file.reg_sp\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4448__A cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output68_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3060_ ih.t.timer_max\[18\] _2757_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__nand2_1
XANTENNA__5043__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5661__A1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4464__A2 _1282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4167__B _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5413__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5701_ net6 _1650_ _2488_ _2507_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a31o_1
X_3962_ _0572_ _0510_ _0401_ _1035_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__o311a_1
XANTENNA__4767__A3 _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3893_ _2893_ _0386_ _0308_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5632_ _1649_ _2446_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4630__B _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5563_ ih.t.timer_max\[10\] _2193_ _2314_ ih.t.timer_max\[2\] _2380_ vssd1 vssd1
+ vccd1 vccd1 _2381_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4514_ _1402_ _1561_ _1569_ _1371_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__a2bb2o_1
X_5494_ _1400_ _2287_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ cu.reg_file.reg_b\[1\] _1281_ _1283_ cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1
+ vccd1 _1504_ sky130_fd_sc_hd__a22o_1
XANTENNA__5742__A _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4376_ _1419_ _1423_ _1437_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__nand3_1
X_6115_ clknet_leaf_28_clk _0149_ net187 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_4
XANTENNA__5461__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3327_ _2878_ _0402_ _2877_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__a21o_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5888__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4455__A2 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6046_ clknet_leaf_6_clk _0084_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_3258_ _0329_ _0332_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or3_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _2925_ _2901_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4391__A1 cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5652__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_output106_A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5038__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5331__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4230_ _1297_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5882__A1 ih.t.timer_max\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4161_ _0516_ _0819_ _1226_ _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__or4b_1
XANTENNA__3082__A ih.t.timer_max\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3112_ _2826_ _2827_ _2849_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__or3_1
X_4092_ _0519_ _1165_ _0614_ _0551_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__o211ai_1
XANTENNA__5634__A1 _2448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3043_ ih.t.count\[25\] _2780_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5398__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4994_ _1975_ _1980_ _1808_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__mux2_1
X_3945_ _0982_ _0997_ _0986_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__nor3b_1
X_5615_ _2430_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
X_3876_ _0887_ _0901_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5546_ mc.cl.next_data\[1\] _2359_ _2324_ _2364_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__a22o_1
X_5477_ _2299_ _2284_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5472__A _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5322__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4428_ _1269_ _1484_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__nor2_1
X_4359_ _1397_ _1395_ _1421_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__a21o_1
XANTENNA__4088__A _0617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4816__A _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6029_ clknet_leaf_2_clk _0067_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5411__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4535__B _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5366__B _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5696__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4116__B2 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5616__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5616__B2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3730_ _0759_ _0783_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__xor2_1
XANTENNA__3349__B_N _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _0645_ _0722_ _0734_ _0736_ _0730_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__a311o_1
X_5400_ _1261_ net131 _2237_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__mux2_1
X_3592_ cu.reg_file.reg_c\[4\] _0427_ _0430_ cu.reg_file.reg_e\[4\] vssd1 vssd1 vccd1
+ vccd1 _0668_ sky130_fd_sc_hd__a22o_1
X_5331_ _0619_ net100 _2206_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5262_ _2164_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4213_ net238 vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__buf_2
X_5193_ _2114_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__clkbuf_2
X_4144_ _0952_ _0955_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4075_ _0767_ _0773_ _1145_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__a31o_1
X_3026_ ih.t.timer_max\[27\] _2763_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__or2_2
XANTENNA__4355__B _1415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4977_ _1963_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3928_ _0994_ _0989_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3859_ _0898_ _0934_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__xor2_2
XFILLER_0_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4346__B2 cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4346__A1 _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5529_ _1649_ _2347_ _2348_ _1641_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3715__A _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3003__A_N net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5141__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5534__B1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5824__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5316__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5840__A cu.reg_file.reg_sp\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output50_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5880_ _1051_ ih.t.timer_max\[1\] _2645_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4900_ cu.pc.pc_o\[7\] cu.pc.pc_o\[8\] _1872_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__and3_1
XANTENNA__4812__A2 _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5448__S0 _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4831_ _1829_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4191__A _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4762_ _1301_ _1300_ _1748_ _1268_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__a31o_1
XANTENNA__5773__A0 cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4693_ ih.t.count\[19\] ih.t.count\[20\] _1711_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3713_ _0664_ _0684_ _0787_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__nand4_1
X_3644_ _0671_ _0681_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3575_ cu.reg_file.reg_l\[5\] _0422_ _0649_ _0650_ _0576_ vssd1 vssd1 vccd1 vccd1
+ _0651_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_87_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5314_ _1052_ net93 _2195_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__mux2_1
X_6294_ clknet_leaf_42_clk _0276_ net153 vssd1 vssd1 vccd1 vccd1 cu.id.opcode\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__3551__A2 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5245_ _1667_ _2147_ _2152_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__o21a_4
Xhold17 ih.t.next_count\[19\] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4500__A1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold28 cu.ir.idx\[0\] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ mc.cl.next_data\[11\] net21 mc.count vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__mux2_1
Xhold39 cu.id.is_halted vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlygate4sd3_1
X_4127_ _0916_ _0944_ _1196_ _1032_ _0918_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__o221a_1
X_4058_ _0757_ _0767_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3009_ ih.t.timer_max\[3\] _2746_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5764__A0 _1089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4319__B2 cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4319__A1 cu.reg_file.reg_a\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3445__A _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5136__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4558__B2 cu.id.imm_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4558__A1 cu.reg_file.reg_sp\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3339__B _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3781__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output98_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5046__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _2908_ _0342_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__nor2_1
XANTENNA__4730__A1 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _2007_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__clkbuf_1
X_3291_ _0350_ _0358_ _0366_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__o21a_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5932_ _2875_ _2467_ _2668_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4914__A cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5863_ _2155_ ih.t.timer_max\[9\] _2636_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _1299_ _1810_ _1815_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__mux2_1
XANTENNA__5746__B1 _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5794_ _2569_ _2572_ _2570_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__a21bo_1
X_4745_ _0296_ _0320_ _1319_ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4676_ ih.t.count\[12\] ih.t.count\[13\] _1696_ ih.t.count\[14\] vssd1 vssd1 vccd1
+ vccd1 _1703_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3772__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3627_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[2\] vssd1 vssd1 vccd1 vccd1 _0703_
+ sky130_fd_sc_hd__o211a_1
X_3558_ _0322_ _0633_ _0443_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6277_ clknet_leaf_16_clk _0259_ net178 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5480__A _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3489_ _0294_ _0372_ _0536_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__o21ai_1
X_5228_ _1415_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__nor2_4
XANTENNA__4485__B1 _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5159_ cu.reg_file.reg_l\[4\] _1189_ _2088_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__mux2_1
XANTENNA__3712__B _0733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_36_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3279__A1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output136_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4453__B _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4530_ _1567_ _1579_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ _1515_ _1516_ _1519_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__o21ai_4
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6200_ clknet_leaf_9_clk net13 net169 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3412_ net147 _0473_ _0479_ _0486_ _0483_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__o2111a_4
X_6131_ clknet_leaf_24_clk _0165_ net192 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_4
X_4392_ cu.reg_file.reg_c\[6\] _1313_ _1451_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_
+ sky130_fd_sc_hd__a211o_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _0412_ _0414_ _0405_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__nor3b_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4628__B _2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6062_ clknet_leaf_25_clk mc.rw.next_state\[2\] net194 vssd1 vssd1 vccd1 vccd1 mc.rw.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _0296_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__clkbuf_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _1994_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5915_ _2663_ cu.ir.idx\[1\] vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__nor2_4
XFILLER_0_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5846_ _2624_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ net8 vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5777_ _2562_ _2563_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__nand2_1
XANTENNA__5195__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4728_ _1672_ _1736_ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4659_ ih.t.count\[8\] _1689_ _1687_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5670__A2 _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5958__A0 cu.id.imm_i\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3984__A2 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5489__A2 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6035__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5324__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5832__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4551__A2_N _1598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3352__B _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5661__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4167__C _1073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3961_ _0781_ _0712_ _0773_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__a21oi_1
X_5700_ _2506_ _1643_ cu.reg_file.reg_mem\[13\] _1646_ vssd1 vssd1 vccd1 vccd1 _2507_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3892_ _0379_ net150 vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5631_ net13 _2345_ _2369_ net6 vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5562_ ih.t.timer_max\[26\] _2146_ _2204_ ih.t.timer_max\[18\] vssd1 vssd1 vccd1
+ vccd1 _2380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4513_ _1567_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5493_ mc.cl.cmp_o _1648_ _1631_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3246__C _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4444_ cu.reg_file.reg_sp\[9\] _1287_ _1285_ cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1
+ vccd1 _1503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4639__A _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4375_ _1419_ _1423_ _1437_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__a21o_1
XANTENNA__5123__B1_N _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3543__A _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6114_ clknet_leaf_27_clk _0148_ net195 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_4
X_3326_ _2899_ _2900_ _2894_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__a21bo_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6045_ clknet_leaf_6_clk _0083_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _2888_ _2927_ _2933_ _2934_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__and4_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ _2892_ _2894_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__nand2_4
XANTENNA__3415__A1 cu.reg_file.reg_c\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3415__B2 cu.reg_file.reg_e\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5829_ cu.reg_file.reg_sp\[11\] _2609_ _2538_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__mux2_1
XANTENNA__5409__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3351__B1 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5144__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5159__A1 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output80_A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5331__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4160_ _1032_ _1227_ _1228_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o211a_2
X_3111_ _2829_ _2831_ _2832_ _2848_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__or4_1
XANTENNA__3893__A1 _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ _0820_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__inv_2
XANTENNA__5095__A0 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3042_ ih.t.timer_max\[25\] _2762_ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__xor2_1
XANTENNA__4194__A _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3810__B _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5398__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4993_ _1978_ _1979_ _1798_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__mux2_1
X_3944_ _0531_ _1018_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3875_ _0877_ _0904_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__xnor2_1
X_5614_ cu.reg_file.reg_mem\[4\] _2429_ _2351_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5545_ _1666_ _2362_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__o21a_1
XANTENNA__5570__A1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5476_ _2225_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__inv_2
XANTENNA__5322__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4427_ cu.reg_file.reg_b\[0\] net144 _1284_ cu.reg_file.reg_h\[0\] _1486_ vssd1 vssd1
+ vccd1 vccd1 _1487_ sky130_fd_sc_hd__a221o_1
X_4358_ _1397_ _1395_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nand3_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4088__B _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4289_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5086__A0 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3309_ _0359_ _2893_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__nand2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6028_ clknet_leaf_2_clk _0066_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4816__B cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5139__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4116__A2 _1186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4521__C1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3183__A cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5077__B1 _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4824__A0 cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5616__A2 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5049__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3660_ _0731_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3591_ cu.reg_file.reg_sp\[4\] _0413_ _0419_ cu.reg_file.reg_h\[4\] _0666_ vssd1
+ vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a221o_1
X_5330_ _2205_ net141 vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__nand2_8
XFILLER_0_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5261_ ih.t.timer_max\[29\] _2163_ _2153_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4212_ _1272_ _1275_ _1276_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__nor4b_1
X_5192_ _1790_ _0352_ _2951_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__or3b_1
XANTENNA__5068__A0 cu.reg_file.reg_c\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4917__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4143_ _0516_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__nor2_4
X_4074_ _0776_ _0805_ _1147_ _0817_ _0777_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a221o_1
XANTENNA__3821__A _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3025_ ih.t.timer_max\[25\] ih.t.timer_max\[26\] _2762_ vssd1 vssd1 vccd1 vccd1 _2763_
+ sky130_fd_sc_hd__or3_1
XANTENNA__4291__B2 _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4976_ cu.pc.pc_o\[13\] _1939_ cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3927_ _1001_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__nand2_1
XANTENNA__3268__A _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3858_ _0920_ _0796_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__nand2_1
X_3789_ _0861_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__xnor2_1
X_5528_ net2 _2148_ _2344_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5459_ _2286_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4546__B _1598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4806__B1 _1807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5658__A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5534__B2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5534__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5840__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5470__A0 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5448__S1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4830_ _0341_ cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5287__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _1769_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4576__A2 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4692_ net213 _1711_ _1713_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[19\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3712_ _0644_ _0733_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3643_ _0652_ _0663_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5313_ _2196_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3574_ cu.reg_file.reg_mem\[5\] _0640_ _0433_ cu.reg_file.reg_a\[5\] vssd1 vssd1
+ vccd1 vccd1 _0650_ sky130_fd_sc_hd__a22o_1
X_6293_ clknet_leaf_42_clk _0275_ net153 vssd1 vssd1 vccd1 vccd1 cu.id.opcode\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_5244_ _1661_ _2151_ _2141_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__o21ba_1
Xhold18 ih.t.count\[10\] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 ih.t.count\[9\] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _2102_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
X_4126_ _0945_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5680__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4057_ _1121_ _1130_ _0817_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__o21a_1
X_3008_ ih.t.timer_max\[0\] ih.t.timer_max\[1\] ih.t.timer_max\[2\] vssd1 vssd1 vccd1
+ vccd1 _2746_ sky130_fd_sc_hd__or3_1
XANTENNA__5213__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4959_ _1945_ _1947_ _1798_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3775__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5516__A1 _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5417__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3339__C _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3636__A _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4730__A2 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3290_ _0359_ _2915_ _0316_ _0363_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__o2111a_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5062__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _2674_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5862_ _2637_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4813_ _1814_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5746__A1 _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5793_ _2576_ _2577_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__nand2_1
X_4744_ _0338_ _1749_ _1750_ _1752_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4675_ ih.t.count\[13\] ih.t.count\[14\] _1699_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__and3_1
X_3626_ _0694_ _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3557_ _0442_ _0437_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__nand2_1
X_6276_ clknet_leaf_16_clk _0258_ net180 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_5227_ _1636_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3488_ cu.reg_file.reg_a\[7\] _0499_ _0494_ cu.reg_file.reg_mem\[7\] _0563_ vssd1
+ vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__a221o_1
XANTENNA__4377__A _1415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4485__B2 cu.id.imm_i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4485__A1 cu.reg_file.reg_sp\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5158_ _2092_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4096__B _0733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5664__A_N _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5089_ _1189_ _1213_ _2035_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__mux2_1
X_4109_ _1168_ _1179_ _1180_ _1182_ _1023_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4840__A cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4986__S _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4173__A0 _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3576__A1_N _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4287__A _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3279__B1_N _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3279__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output129_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5520__S0 _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5728__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4460_ _1371_ _1517_ _1518_ _1511_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_68_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4896__S _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3411_ _0483_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nor2_2
X_4391_ cu.pc.pc_o\[6\] _1322_ _1315_ cu.reg_file.reg_e\[6\] _1452_ vssd1 vssd1 vccd1
+ vccd1 _1453_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6130_ clknet_leaf_20_clk _0164_ net172 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_4
X_3342_ _0407_ _0417_ _0409_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ clknet_leaf_25_clk mc.rw.next_state\[1\] net194 vssd1 vssd1 vccd1 vccd1 mc.rw.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4467__A1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _2874_ _2927_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__nor2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ cu.reg_file.reg_a\[4\] _1993_ _1985_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__mux2_1
XANTENNA__4925__A _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5914_ _2351_ _2664_ _2665_ net225 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5845_ cu.reg_file.reg_sp\[13\] _2623_ _2538_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2988_ net2 vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5776_ cu.reg_file.reg_sp\[5\] _2535_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__nand2_1
X_4727_ ih.t.count\[30\] ih.t.count\[31\] _1732_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4658_ ih.t.count\[8\] _1689_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3609_ _0664_ _0684_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__nor2_1
X_4589_ _1329_ _1401_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__nand2_4
X_6259_ clknet_leaf_4_clk _0241_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[15\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__5407__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5958__A1 _2391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4570__A _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5385__B _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6075__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6004__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4449__A1 cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4449__B2 cu.id.imm_i\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4167__D _1089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4745__A _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3960_ _0781_ _0712_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__or2_1
XANTENNA__4621__A1 _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3891_ _2883_ _0304_ _0966_ _2893_ _0301_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ net73 _1648_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5561_ net78 _1633_ _2375_ _2378_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4512_ _1566_ _1561_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__or2_1
X_5492_ net76 _1633_ _2309_ _2311_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4443_ _1382_ _1498_ _1499_ _1502_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__a31o_2
X_4374_ _1435_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6113_ clknet_leaf_28_clk _0147_ net186 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_2
X_3325_ _0395_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or2_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ clknet_leaf_5_clk _0082_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3256_ _0330_ _0331_ _2932_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a21oi_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _2901_ _2923_ _2874_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__or3b_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5828_ _1222_ _2608_ _2545_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5759_ cu.reg_file.reg_sp\[3\] _2534_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4128__B1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3453__B _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3575__D1 _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3590__A1 cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5335__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3590__B2 cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output73_A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3110_ _2834_ _2843_ _2844_ _2847_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ _1129_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5095__A1 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3041_ _2763_ _2777_ ih.t.count\[26\] vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5070__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4992_ _1263_ _1975_ _1794_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _0971_ _0986_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__or2_2
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3874_ _0856_ _0908_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5613_ _2425_ _2426_ _2428_ _1641_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__o22a_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3566__D1 _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5544_ ih.t.timer_max\[17\] _2151_ _2319_ ih.t.timer_max\[1\] _1661_ vssd1 vssd1
+ vccd1 vccd1 _2363_ sky130_fd_sc_hd__a221o_1
XANTENNA__5570__A2 _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5475_ _2298_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3581__A1 cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4426_ cu.reg_file.reg_d\[0\] _1282_ _1286_ cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1
+ vccd1 _1486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4357_ _1419_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__nand2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3704__D _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4288_ _2698_ mc.rw.state\[1\] mc.rw.state\[0\] vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__or3_1
XANTENNA__5086__A1 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3308_ _0317_ _0379_ _0383_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__or3_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _0310_ _0311_ _0312_ _0314_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__or4b_4
X_6027_ clknet_leaf_2_clk _0065_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5561__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3572__B2 cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3572__A1 cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3464__A cu.reg_file.reg_a\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6197__D net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4994__S _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4521__B1 _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5077__A1 _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output111_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3639__A _0587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3590_ cu.reg_file.reg_d\[4\] _0415_ _0432_ cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1
+ vccd1 _0666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3563__A1 cu.reg_file.reg_c\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5260_ _1144_ _1209_ _1666_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3315__A1 _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4211_ _2912_ _0583_ _1277_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__a31o_2
X_5191_ _2113_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4917__B cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5068__A1 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4142_ _0956_ _1205_ _1206_ _0957_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__o221a_1
XANTENNA__3079__B1 ih.t.timer_max\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4073_ _0811_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nand2_1
X_3024_ ih.t.timer_max\[24\] _2761_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__or2_2
XFILLER_0_78_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4975_ cu.pc.pc_o\[14\] cu.pc.pc_o\[13\] _1939_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__and3_1
XANTENNA__4579__B1 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _0981_ _0998_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__nand2_1
XANTENNA__6107__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3857_ _0865_ _0925_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__xnor2_1
X_3788_ cu.reg_file.reg_mem\[12\] _0640_ _0862_ _0863_ vssd1 vssd1 vccd1 vccd1 _0864_
+ sky130_fd_sc_hd__a211oi_2
X_5527_ net2 _2345_ _2346_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__a21o_1
XANTENNA__3554__A1 cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3284__A _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5458_ net60 _2085_ _2285_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__mux2_1
X_5389_ _2239_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
X_4409_ cu.reg_file.reg_sp\[7\] _0993_ _1344_ cu.id.cb_opcode_x\[1\] _1324_ vssd1
+ vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4806__A1 _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4843__A cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4034__A2 _0733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3793__A1 cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5534__A2 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3922__A _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3848__A2 _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output36_A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5470__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4430__C1 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4760_ net236 _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__or2_1
X_4691_ ih.t.count\[19\] _1711_ _1670_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__o21ai_1
X_3711_ _0759_ _0763_ _0783_ _0785_ _0786_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__a311o_2
XANTENNA__3784__A1 cu.reg_file.reg_a\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3784__B2 cu.reg_file.reg_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3642_ _0702_ _0716_ _0717_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__o21ai_2
X_5312_ _0619_ net92 _2195_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3573_ cu.reg_file.reg_c\[5\] _0427_ _0430_ cu.reg_file.reg_e\[5\] vssd1 vssd1 vccd1
+ vccd1 _0649_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6292_ clknet_leaf_42_clk _0274_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.alu_opcode\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_5243_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__buf_2
Xhold19 ih.t.next_count\[10\] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _1647_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__and2_1
X_4125_ _0942_ _0943_ _0944_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _0804_ _0811_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__and2_1
X_3007_ _2736_ _2737_ _2738_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__or4_4
XANTENNA__5759__A cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4958_ _1945_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__or2_1
X_4889_ cu.pc.pc_o\[7\] _1872_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__xor2_1
X_3909_ _0310_ _0328_ _0740_ _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__nor4_1
XFILLER_0_19_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3775__B2 cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3775__A1 cu.reg_file.reg_sp\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5494__A _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4724__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5452__A1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5452__B2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3636__B _0598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3518__A1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5343__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5930_ _2936_ _2448_ _2668_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__mux2_1
X_5861_ _2144_ ih.t.timer_max\[8\] _2636_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__mux2_1
X_4812_ _2948_ _1808_ _1813_ _1484_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__a22o_4
XANTENNA__5746__A2 _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5792_ cu.reg_file.reg_sp\[7\] _2535_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4743_ _2907_ _0311_ _0379_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4674_ net218 _1699_ _1701_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[13\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5708__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3625_ _0576_ _0695_ _0697_ _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3556_ _0623_ _0627_ _0630_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__o31a_4
X_6275_ clknet_leaf_15_clk _0257_ net175 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_5226_ _2135_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3487_ cu.pc.pc_o\[7\] _0501_ _0498_ cu.alu_f\[7\] _0504_ vssd1 vssd1 vccd1 vccd1
+ _0563_ sky130_fd_sc_hd__a221o_1
XANTENNA__4377__B _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5682__B2 ih.t.timer_max\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5157_ cu.reg_file.reg_l\[3\] _1187_ _2088_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__mux2_1
X_5088_ _2046_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
X_4108_ _0996_ _1003_ _1181_ _1010_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__or4b_2
X_4039_ _1060_ _0599_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nand2_1
XANTENNA__6193__RESET_B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4173__A1 _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5520__S1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4936__A0 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3647__A _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3410_ net148 _0460_ _0462_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ cu.reg_file.reg_sp\[6\] _0993_ _1344_ _0387_ _1324_ vssd1 vssd1 vccd1 vccd1
+ _1452_ sky130_fd_sc_hd__a221o_1
X_3341_ _0412_ _0405_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__or2_4
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A0 cu.reg_file.reg_e\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6060_ clknet_leaf_25_clk mc.rw.next_state\[0\] net194 vssd1 vssd1 vccd1 vccd1 mc.rw.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _2942_ _0345_ _0347_ _0336_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__o31a_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _1189_ _1213_ _0368_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3427__B1 _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5913_ _2947_ _1482_ _2664_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4941__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5844_ _1209_ _2622_ _2115_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5248__S _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2987_ _2721_ ih.ih.ih.prev_data\[9\] _2722_ ih.ih.ih.prev_data\[14\] _2725_ vssd1
+ vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5775_ cu.reg_file.reg_sp\[5\] _2535_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4726_ ih.t.count\[30\] _1732_ ih.t.count\[31\] vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__a21o_1
X_4657_ _1689_ _1690_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[7\] sky130_fd_sc_hd__nor2_1
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5352__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3608_ _0682_ _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4588_ mc.cl.cmp_o _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__or2b_2
X_3539_ _0572_ _0573_ _0608_ _0613_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__o2111a_1
XANTENNA__3902__B2 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6258_ clknet_leaf_4_clk _0240_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[14\]
+ sky130_fd_sc_hd__dfstp_2
X_6189_ clknet_leaf_22_clk _0222_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5209_ _1364_ _2125_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__or2_1
XANTENNA__5407__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4570__B _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4997__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5343__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5894__A1 _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5646__A1 _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4449__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4909__B1 _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3890_ _2917_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nand2_1
XANTENNA__5068__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5560_ net110 _2147_ _2225_ net118 _2377_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__a221o_1
X_4511_ _1566_ _1561_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__nand2_1
X_5491_ net100 _2205_ _2310_ _2257_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5592__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4442_ _1496_ _1500_ _1501_ _1371_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__a22o_1
X_4373_ _1396_ _1434_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6112_ clknet_leaf_13_clk _0146_ net173 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XANTENNA__4001__A _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _2950_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3255_ cu.id.opcode\[0\] cu.id.alu_opcode\[3\] cu.id.alu_opcode\[1\] _2892_ vssd1
+ vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__or4bb_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ clknet_leaf_4_clk _0081_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _2894_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout172_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4612__A2 _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5767__A cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5827_ _2606_ _2607_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5758_ _2547_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
X_4709_ ih.t.count\[25\] _1723_ _1670_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3584__C1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5689_ net3 _1650_ _2488_ _2498_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a31o_1
XANTENNA__4300__A1 cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4565__B _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4300__B2 cu.reg_file.reg_l\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5316__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5867__A1 ih.t.timer_max\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4119__B2 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5619__B2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5619__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output66_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ ih.t.count\[26\] _2763_ _2777_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4991_ cu.pc.pc_o\[15\] _1977_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__xor2_1
X_3942_ _1000_ _1008_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3873_ _0845_ _0910_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__xnor2_1
X_5612_ _1649_ _2427_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5543_ _1400_ _2361_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5474_ net64 _2085_ _2297_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__mux2_1
XANTENNA__3581__A2 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4425_ _1269_ _1484_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__or2_4
XFILLER_0_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4356_ _1332_ _1417_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nand2_1
X_3307_ _2905_ _0380_ _0381_ _0382_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__or4_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4287_ _1348_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__buf_4
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ clknet_leaf_9_clk _0064_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _2910_ _0313_ _0305_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__or3_1
X_3169_ _2887_ _2891_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4349__A1 cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4521__A1 cu.reg_file.reg_sp\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3911__C _0379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3639__B _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4042__A2_N _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3655__A _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ _2877_ _0336_ _0436_ _0293_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5190_ _2111_ _2112_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__and2_1
XANTENNA__5081__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4141_ _0817_ _0942_ _1210_ _0933_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__a22oi_1
XANTENNA__3079__A1 ih.t.timer_max\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4072_ _0808_ _0810_ _0805_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3023_ ih.t.timer_max\[22\] ih.t.timer_max\[23\] _2760_ vssd1 vssd1 vccd1 vccd1 _2761_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4579__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4579__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4974_ _1962_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__clkbuf_1
X_3925_ _0998_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5528__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3856_ _0829_ _0919_ _0931_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3787_ cu.reg_file.reg_b\[4\] _0426_ _0429_ cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1
+ vccd1 _0863_ sky130_fd_sc_hd__a22o_1
X_5526_ net16 _2179_ _2279_ ih.input_handler_enable vssd1 vssd1 vccd1 vccd1 _2346_
+ sky130_fd_sc_hd__a22o_1
X_5457_ _1633_ _2284_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4408_ cu.reg_file.reg_l\[7\] _1317_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__and2_1
XANTENNA__4503__A1 cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5388_ _1052_ net125 _2237_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__mux2_1
XANTENNA__5700__B1 cu.reg_file.reg_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4503__B2 cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4339_ _1393_ _1401_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6009_ clknet_leaf_31_clk _0047_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4806__A2 _1256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4843__B cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4990__A1 _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3793__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3475__A _0399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3710_ _0701_ _0694_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__and2b_1
X_4690_ _1711_ _1712_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[18\] sky130_fd_sc_hd__nor2_1
XFILLER_0_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _0694_ _0701_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5930__A0 _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3572_ cu.reg_file.reg_sp\[5\] _0636_ _0419_ cu.reg_file.reg_h\[5\] _0647_ vssd1
+ vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__a221o_1
X_5311_ net141 _2194_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__nand2_8
XFILLER_0_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6291_ clknet_leaf_42_clk _0273_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.alu_opcode\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_5242_ _2145_ _2149_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__or2_2
XANTENNA__4497__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5173_ mc.cl.next_data\[10\] net20 mc.count vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__mux2_1
X_4124_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__buf_4
Xinput1 interrupt_gpio_in vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__dlymetal6s2s_1
X_4055_ _1127_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3006_ _2739_ net33 ih.gpio_interrupt_mask\[6\] _2742_ _2743_ vssd1 vssd1 vccd1 vccd1
+ _2744_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5749__A0 cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4957_ _1920_ _1922_ _1932_ _1946_ _1921_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5775__A cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4888_ _1883_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__clkbuf_1
X_3908_ _2918_ _0966_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3839_ _0777_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__nand2_1
XANTENNA__3295__A _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5509_ _2169_ _2312_ _2328_ _2136_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__o211a_1
XANTENNA__4854__A _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5912__B1 _1484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5860_ _1667_ _2194_ _2635_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__o21ai_4
X_4811_ _1301_ _1775_ _1811_ _1812_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5791_ cu.reg_file.reg_sp\[7\] _2535_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4742_ _0314_ _1741_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__nor2_1
X_4673_ ih.t.count\[13\] _1699_ _1670_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3827__B _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3624_ cu.reg_file.reg_l\[3\] _0422_ _0698_ _0699_ _0440_ vssd1 vssd1 vccd1 vccd1
+ _0700_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3555_ _0295_ _2921_ _0536_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__o21ai_1
X_6274_ clknet_leaf_15_clk _0256_ net177 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3486_ cu.reg_file.reg_h\[7\] _0495_ _0539_ cu.reg_file.reg_sp\[7\] _0561_ vssd1
+ vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__a221o_1
X_5225_ _1261_ ih.gpio_interrupt_mask\[7\] _2127_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__mux2_1
X_5156_ _2091_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__clkbuf_1
X_5087_ cu.reg_file.reg_d\[3\] _2045_ _2039_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__mux2_1
X_4107_ _1018_ _1019_ _0395_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__a21oi_1
X_4038_ _0588_ _0610_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ clknet_leaf_29_clk _0027_ net188 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4584__A _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5189__A1 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5354__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output96_A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3340_ cu.reg_file.reg_sp\[0\] _0413_ _0415_ cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1
+ vccd1 _0416_ sky130_fd_sc_hd__a22o_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3271_ _0301_ _0346_ _0316_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__o21ai_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _1992_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__clkbuf_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5912_ _2663_ _1644_ _1484_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4941__B cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5843_ _2620_ _2621_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__xnor2_1
X_2986_ _2723_ ih.ih.ih.prev_data\[5\] _2724_ ih.ih.ih.prev_data\[10\] vssd1 vssd1
+ vccd1 vccd1 _2725_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5774_ _2561_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4725_ net207 _1732_ _1735_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[30\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4656_ net227 _1686_ _1687_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__o21ai_1
X_4587_ _1374_ _1625_ _1630_ _1417_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__a211o_1
XANTENNA__5352__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3607_ _0681_ _0671_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ _0549_ _0555_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3469_ _0537_ _0538_ _0543_ _0544_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__o31a_4
X_6257_ clknet_leaf_3_clk _0239_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[13\]
+ sky130_fd_sc_hd__dfstp_2
X_6188_ clknet_leaf_22_clk _0221_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5208_ _1634_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3666__A1 cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5139_ _2079_ cu.reg_file.reg_h\[5\] _2069_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__mux2_1
XANTENNA__3666__B2 cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5040__A0 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5591__A1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5591__B2 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5343__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5894__A2 _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6084__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3658__A _0733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5031__A0 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4510_ _1517_ _1530_ _1545_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__and3_1
X_5490_ net108 _2146_ _2193_ net92 vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4441_ _1478_ _1496_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__nor2_1
XANTENNA__5084__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4372_ _1396_ _1434_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__or2_1
X_6111_ clknet_leaf_31_clk _0145_ net183 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A0 _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3323_ _2893_ _0386_ _0324_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__a31o_2
XFILLER_0_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A2 _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3254_ _2894_ _2884_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__or2b_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ clknet_leaf_40_clk _0080_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_l\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _2920_ _2921_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3568__A _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5826_ _2597_ _2600_ _2598_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__a21bo_1
X_2969_ _2708_ vssd1 vssd1 vccd1 vccd1 mc.cc.enable sky130_fd_sc_hd__inv_2
XFILLER_0_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5757_ cu.reg_file.reg_sp\[2\] _2546_ _2539_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4708_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[24\] sky130_fd_sc_hd__nor2_1
XANTENNA__5783__A cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3584__B1 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5688_ _2497_ _1643_ cu.reg_file.reg_mem\[10\] _1646_ vssd1 vssd1 vccd1 vccd1 _2498_
+ sky130_fd_sc_hd__a2bb2o_1
X_4639_ _1672_ _1676_ _1677_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__and3_1
XANTENNA__3336__B1 cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6309_ clknet_leaf_20_clk _0291_ net182 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5089__A0 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5261__A0 ih.t.timer_max\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4581__B _1372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3909__C _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5316__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4119__A2 _1186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3327__B1 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5619__A2 _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4827__B1 cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4990_ _1233_ _1969_ _1976_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3802__B2 cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3941_ _1013_ _1014_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3872_ _0833_ _0912_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5611_ net12 _2345_ _2369_ net5 vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__a22o_1
X_5542_ ih.t.timer_max\[9\] _2193_ _2314_ ih.t.timer_max\[1\] _2360_ vssd1 vssd1 vccd1
+ vccd1 _2361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5473_ _2296_ _2284_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4424_ _1482_ _1483_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4355_ _1396_ _1415_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__nand2_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _2903_ _0313_ _0329_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o21bai_4
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ mc.rw.state\[1\] mc.rw.state\[0\] _2698_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__o21a_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ clknet_leaf_31_clk _0063_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _2892_ cu.id.opcode\[0\] vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__or2_2
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3168_ _2893_ _2896_ _2904_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3099_ ih.t.count\[0\] _2836_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5988__RESET_B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5809_ _2590_ _2591_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4285__A1 _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5482__A0 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4592__A _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5644__A_N _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5234__A0 ih.t.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3001__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3796__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5537__B2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5537__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3936__A _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5362__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4140_ _0817_ _0941_ _0776_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__a21o_1
X_4071_ _0765_ _0766_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3022_ ih.t.timer_max\[21\] _2759_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__or2_2
XANTENNA__5598__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5225__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4579__A2 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4973_ cu.pc.pc_o\[13\] _1961_ _1814_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3924_ _0976_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__nor2_1
XANTENNA__3787__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3855_ _0829_ _0919_ _0930_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3786_ cu.reg_file.reg_sp\[12\] _0636_ _0748_ cu.reg_file.reg_h\[4\] vssd1 vssd1
+ vccd1 vccd1 _0862_ sky130_fd_sc_hd__a22o_1
X_5525_ _1625_ _2344_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__nand2_2
XANTENNA__4751__A2 _1739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5456_ _2283_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4407_ cu.id.cb_opcode_x\[1\] _1295_ _1298_ cu.pc.pc_o\[7\] _1306_ vssd1 vssd1 vccd1
+ vccd1 _1468_ sky130_fd_sc_hd__a221o_1
XANTENNA__4503__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5387_ _2238_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5700__B2 _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4338_ _1356_ _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__o21ai_1
X_4269_ _1330_ _1334_ _1336_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6008_ clknet_leaf_5_clk _0046_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5519__A1 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5519__B2 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3491__A _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4258__A1 cu.reg_file.reg_sp\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4258__B2 _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4430__A1 cu.id.imm_i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4430__B2 cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _0711_ _0714_ _0715_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__a21oi_2
XANTENNA__5930__A1 _2448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3571_ cu.reg_file.reg_d\[5\] _0415_ _0432_ cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1
+ vccd1 _0647_ sky130_fd_sc_hd__a22o_1
X_5310_ _2193_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6290_ clknet_leaf_42_clk _0272_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.alu_opcode\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5241_ _1374_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__nor2_1
XANTENNA__5092__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4497__A1 cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4497__B2 cu.reg_file.reg_sp\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5172_ _2100_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
X_4123_ _1126_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__clkbuf_4
Xinput2 keypad_input[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
X_4054_ _1110_ _1126_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__and2_1
X_3005_ net75 net34 ih.gpio_interrupt_mask\[7\] vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__and3b_1
XANTENNA__3457__C1 cu.reg_file.reg_l\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ cu.pc.pc_o\[11\] _1521_ _1233_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4887_ cu.pc.pc_o\[6\] _1882_ _1815_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3907_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3838_ _0833_ _0912_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__o21a_1
XANTENNA__4171__S _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5508_ _2125_ _2325_ _2326_ ih.gpio_interrupt_mask\[0\] _2327_ vssd1 vssd1 vccd1
+ vccd1 _2328_ sky130_fd_sc_hd__a221o_1
XANTENNA__5791__A cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3769_ _0844_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__inv_2
X_5439_ _2269_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4854__B cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3448__C1 _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4176__A0 _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6038__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _1300_ _1768_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__xor2_1
XANTENNA__5600__B1 _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5790_ _2575_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4403__B2 cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4403__A1 cu.reg_file.reg_a\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5087__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4741_ _2922_ _0303_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4672_ _1699_ _1700_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[12\] sky130_fd_sc_hd__nor2_1
XFILLER_0_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5903__A1 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3623_ cu.reg_file.reg_mem\[3\] _0418_ _0433_ cu.reg_file.reg_a\[3\] vssd1 vssd1
+ vccd1 vccd1 _0699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ cu.reg_file.reg_b\[6\] _0502_ _0499_ cu.reg_file.reg_a\[6\] _0629_ vssd1 vssd1
+ vccd1 vccd1 _0630_ sky130_fd_sc_hd__a221o_1
X_6273_ clknet_leaf_15_clk _0255_ net175 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3485_ cu.reg_file.reg_b\[7\] _0502_ _0492_ cu.reg_file.reg_d\[7\] vssd1 vssd1 vccd1
+ vccd1 _0561_ sky130_fd_sc_hd__a22o_1
X_5224_ _2134_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout195_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5419__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5155_ cu.reg_file.reg_l\[2\] _1074_ _2088_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__mux2_1
X_5086_ _1187_ _1222_ _2035_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__mux2_1
X_4106_ cu.alu_f\[2\] _1013_ _1012_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__o21a_1
X_4037_ _0611_ _0643_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ clknet_leaf_29_clk _0026_ net188 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_4939_ _1521_ _1907_ cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4584__B _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output89_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3270_ _2874_ _2927_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__or2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4494__B _1545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5911_ cu.ir.idx\[0\] vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__inv_2
XANTENNA__5821__A0 cu.reg_file.reg_sp\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5842_ _2611_ _2614_ _2612_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5585__C1 _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5773_ cu.reg_file.reg_sp\[4\] _2560_ _2539_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__mux2_1
X_4724_ net207 _1732_ _1670_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2985_ net3 vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4655_ ih.t.count\[6\] ih.t.count\[7\] _1683_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__and3_1
XANTENNA__5888__A0 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4586_ _1434_ _1462_ _1473_ _1629_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__or4_2
XANTENNA__3899__C1 _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3606_ _0671_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3537_ _0610_ _0612_ net143 _0601_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a211o_1
X_3468_ _0294_ _0360_ _0536_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o21ai_1
X_6256_ clknet_leaf_2_clk _0238_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[12\]
+ sky130_fd_sc_hd__dfstp_2
X_5207_ _2124_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
X_6187_ clknet_leaf_22_clk _0220_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3666__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3399_ cu.id.cb_opcode_z\[1\] _2918_ _0364_ _0470_ _0474_ vssd1 vssd1 vccd1 vccd1
+ _0475_ sky130_fd_sc_hd__o221a_1
X_5138_ _1209_ _1144_ _2066_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5069_ _2032_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5812__A0 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5040__A1 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6312__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output127_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5031__A1 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3593__A1 cu.reg_file.reg_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3593__B2 cu.reg_file.reg_a\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4440_ _2701_ _1478_ _1353_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4489__B _1545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6110_ clknet_leaf_11_clk _0144_ net167 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XANTENNA__6200__D net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4371_ _1428_ _1429_ _1433_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__o21a_2
XANTENNA__5098__A1 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3322_ _0361_ _0388_ _0397_ _2891_ _2887_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__a311o_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _2925_ _2932_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__nor2_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ clknet_leaf_34_clk _0079_ net164 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_3184_ cu.id.cb_opcode_x\[0\] vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__inv_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout158_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5825_ _2604_ _2605_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__nand2_1
X_2968_ _2705_ _2707_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__and2_2
XFILLER_0_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5756_ _1073_ _2544_ _2545_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__mux2_1
X_4707_ net232 _1720_ _1687_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5275__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5687_ mc.cl.next_data\[10\] _2359_ _2490_ _2496_ vssd1 vssd1 vccd1 vccd1 _2497_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3584__A1 cu.reg_file.reg_e\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3584__B2 cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4638_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] vssd1 vssd1 vccd1 vccd1 _1677_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4569_ _1382_ _1616_ _1617_ _1621_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__a31o_1
XFILLER_0_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6308_ clknet_leaf_31_clk _0290_ net183 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5089__A1 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6239_ clknet_leaf_25_clk ih.t.next_count\[27\] net193 vssd1 vssd1 vccd1 vccd1 ih.t.count\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4619__S _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A1 _2163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3575__A1 cu.reg_file.reg_l\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5721__C1 _2870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4827__A1 _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5252__A1 _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3940_ _0976_ _0981_ _1008_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3802__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3871_ _0817_ _0945_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__and3_1
X_5610_ net72 _1648_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5541_ ih.t.timer_max\[25\] _2146_ _2204_ ih.t.timer_max\[17\] vssd1 vssd1 vccd1
+ vccd1 _2360_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5095__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5472_ _2147_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4423_ _1268_ _2947_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__or2_2
XFILLER_0_1_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4354_ _2701_ _1404_ _1417_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__and3_1
X_3305_ _0361_ _0376_ _2926_ _2928_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__a211o_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _1335_ _1349_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__o21a_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ clknet_leaf_5_clk _0062_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5491__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _2894_ _2916_ _2939_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_55_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167_ _2898_ _2903_ vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__or2_2
X_3098_ ih.t.timer_max\[1\] ih.t.count\[1\] vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4174__S _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_18_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5808_ cu.reg_file.reg_sp\[9\] _2536_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__nand2_1
XANTENNA__4754__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5739_ cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4203__A _1270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5482__A1 _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5234__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3796__A1 cu.reg_file.reg_sp\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__B2 cu.reg_file.reg_h\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5537__A2 _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3936__B _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5209__A _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output71_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _1143_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3021_ ih.t.timer_max\[19\] ih.t.timer_max\[20\] _2758_ vssd1 vssd1 vccd1 vccd1 _2759_
+ sky130_fd_sc_hd__or3_1
XANTENNA__4783__A _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5598__B _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4433__C1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4972_ _1953_ _1960_ _1808_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _0980_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__inv_2
XANTENNA__3787__B2 cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3787__A1 cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3854_ _0842_ _0929_ _0843_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3785_ cu.id.imm_i\[12\] _0739_ _0860_ _0653_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__a22oi_4
X_5524_ _1666_ _2191_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__nand2_1
X_5455_ _1364_ _2274_ _2275_ _2282_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4406_ _1271_ _1466_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__nor2_1
XANTENNA__5161__A0 cu.reg_file.reg_l\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5386_ _0619_ net124 _2237_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4337_ mc.rw.state\[1\] mc.rw.state\[0\] _2698_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__o21ai_4
XANTENNA__5692__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4268_ mc.rw.state\[2\] _2705_ _2707_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__o211a_1
X_6007_ clknet_2_3__leaf_clk _0045_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3219_ _0294_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6156__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4199_ _0323_ _1266_ _2912_ _2937_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4258__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3466__B1 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4718__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ _0295_ _0634_ _0373_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__or3b_1
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _1329_ _1372_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__or2_2
XANTENNA__5373__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4497__A2 _1282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5694__B2 ih.t.timer_max\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5171_ _1647_ _2099_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__and2_1
X_4122_ net208 _1186_ _0370_ _1192_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a22o_1
X_4053_ _1110_ _1126_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nor2_1
X_3004_ _2740_ net32 ih.gpio_interrupt_mask\[5\] _2741_ vssd1 vssd1 vccd1 vccd1 _2742_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__5402__A _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 keypad_input[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_4
XFILLER_0_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4955_ _1943_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3906_ _0976_ _0981_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__nand2_1
X_4886_ _1874_ _1881_ _1809_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__mux2_1
XANTENNA__4709__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3837_ _0829_ _0832_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3768_ _0842_ _0843_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__and2b_1
X_5507_ _1415_ _1629_ _1637_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__nor3_4
XFILLER_0_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5283__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3699_ _0620_ _0547_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5438_ _2022_ net73 _2268_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__mux2_1
XANTENNA__5685__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5369_ _1052_ net117 _2226_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3448__B1 _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5972__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5373__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4176__A1 _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5912__A2 _1644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4598__A _1415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6007__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4939__B1 cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__B2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4740_ _2908_ _0361_ _0968_ _0313_ _0326_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__o32a_1
X_4671_ ih.t.count\[12\] _1696_ _1687_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6203__D net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3622_ cu.reg_file.reg_c\[3\] _0427_ _0430_ cu.reg_file.reg_e\[3\] vssd1 vssd1 vccd1
+ vccd1 _0698_ sky130_fd_sc_hd__a22o_1
XANTENNA__3914__A1 _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3553_ cu.pc.pc_o\[6\] _0501_ _0628_ cu.reg_file.reg_mem\[6\] _0536_ vssd1 vssd1
+ vccd1 vccd1 _0629_ sky130_fd_sc_hd__a221o_1
X_6272_ clknet_leaf_15_clk _0254_ net175 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3484_ cu.reg_file.reg_c\[7\] _0485_ _0489_ cu.reg_file.reg_e\[7\] _0559_ vssd1 vssd1
+ vccd1 vccd1 _0560_ sky130_fd_sc_hd__a221o_1
X_5223_ _1194_ ih.gpio_interrupt_mask\[6\] _2127_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ _2090_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5419__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4105_ _0395_ _1169_ _1170_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout188_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5085_ _2044_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4036_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ clknet_leaf_28_clk _0025_ net186 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[9\] sky130_fd_sc_hd__dfrtp_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4938_ cu.pc.pc_o\[11\] _1521_ _1907_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__and3_1
XANTENNA_30 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4869_ _1851_ _1854_ _1852_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4158__B2 _0916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5107__A0 cu.reg_file.reg_e\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6171__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4584__C _1545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5594__A0 cu.reg_file.reg_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5897__A1 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4121__A _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4321__A1 cu.reg_file.reg_c\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ _2662_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4791__A _1186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5098__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5841_ _2618_ _2619_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2984_ net13 vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__inv_2
XANTENNA__4388__B2 cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4388__A1 _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5772_ _1160_ _2559_ _2545_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4723_ _1734_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[29\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__3200__A _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5337__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ _1686_ _1688_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4585_ _1393_ _1627_ _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__or3_4
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3605_ _0653_ _0673_ _0675_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__o22a_2
XFILLER_0_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4560__A1 cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3536_ _0447_ _0611_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6255_ clknet_leaf_2_clk _0237_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[11\]
+ sky130_fd_sc_hd__dfstp_2
X_5206_ _2122_ mc.cc.count\[3\] _2120_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__and3b_1
X_3467_ cu.reg_file.reg_sp\[1\] _0539_ _0540_ _0541_ _0542_ vssd1 vssd1 vccd1 vccd1
+ _0543_ sky130_fd_sc_hd__a2111o_1
XANTENNA__4966__A _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6186_ clknet_leaf_22_clk _0219_ net190 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3398_ _2900_ _2878_ _0301_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__a21o_1
X_5137_ _2078_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__clkbuf_1
X_5068_ cu.reg_file.reg_c\[6\] _1193_ _2025_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__mux2_1
X_4019_ _0801_ _0812_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5576__B1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4876__A cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4595__B _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3290__A1 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4370_ cu.reg_file.reg_c\[5\] _1313_ _1430_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__4542__B2 cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4542__A1 cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3321_ _0375_ _0396_ cu.id.cb_opcode_x\[1\] _0387_ vssd1 vssd1 vccd1 vccd1 _0397_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__5381__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4786__A _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _2887_ _2891_ _0323_ _0327_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__or4b_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6040_ clknet_leaf_33_clk _0078_ net164 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5824_ cu.reg_file.reg_sp\[11\] _2536_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2967_ _2701_ _2706_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__nor2_1
X_5755_ _2115_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__clkbuf_4
X_4706_ ih.t.count\[24\] _1720_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__and2_1
X_5686_ ih.t.timer_max\[26\] _2151_ _2320_ ih.t.timer_max\[10\] vssd1 vssd1 vccd1
+ vccd1 _2496_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4637_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] vssd1 vssd1 vccd1 vccd1 _1676_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4568_ _1618_ _1619_ _1620_ _1614_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5291__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6307_ clknet_leaf_7_clk _0289_ net165 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_4499_ cu.id.imm_i\[12\] _1294_ _1297_ cu.pc.pc_o\[12\] _1488_ vssd1 vssd1 vccd1
+ vccd1 _1555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3519_ cu.id.cb_opcode_y\[1\] _0361_ _0437_ _0340_ _0583_ vssd1 vssd1 vccd1 vccd1
+ _0595_ sky130_fd_sc_hd__a221o_1
X_6238_ clknet_leaf_24_clk ih.t.next_count\[26\] net193 vssd1 vssd1 vccd1 vccd1 ih.t.count\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ clknet_leaf_3_clk _0203_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5797__A0 cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4524__A1 _1304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4827__A2 cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3015__A ih.t.timer_max\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5788__A0 _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3870_ _0833_ _0930_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5540_ _2313_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5960__A0 cu.id.imm_i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5471_ _2295_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
X_4422_ _1301_ _1300_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__or2_1
X_4353_ _1306_ _1410_ _1414_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4284_ _2696_ _1333_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__or2_2
X_3304_ _0296_ _2891_ _0318_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__or3_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ clknet_leaf_31_clk _0061_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3235_ _2885_ _2927_ _0309_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__and3_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5491__A2 _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _2901_ _2902_ _2884_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__or3b_2
X_3097_ ih.t.timer_max\[4\] _2747_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3999_ _1063_ _1070_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5807_ cu.reg_file.reg_sp\[9\] _2535_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__or2_1
X_5738_ net25 _2519_ _2529_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5669_ _2169_ _2474_ _2481_ _2136_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5942__A0 cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5924__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5170__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output64_A net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3020_ ih.t.timer_max\[18\] _2757_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3484__A1 cu.reg_file.reg_c\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6206__D net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4433__B1 _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4971_ _1958_ _1959_ _1798_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3922_ _0986_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__nor2_1
XANTENNA__3787__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3853_ _0854_ _0927_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3784_ cu.reg_file.reg_a\[4\] _0625_ _0628_ cu.reg_file.reg_mem\[12\] _0859_ vssd1
+ vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__a221o_1
X_5523_ _2275_ _2342_ _1648_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__and3b_1
X_5454_ _1369_ _2276_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__o21ai_1
X_5385_ net141 _2236_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__nand2_8
X_4405_ cu.reg_file.reg_c\[7\] _1281_ _1465_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5161__A1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4677__C _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4336_ _1348_ _1373_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__nor2_8
XFILLER_0_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4267_ _1329_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__inv_2
X_6006_ clknet_leaf_31_clk _0044_ net183 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_3218_ _0293_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__clkbuf_4
X_4198_ _2877_ _0436_ _0469_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__and3_1
X_3149_ cu.id.opcode\[6\] cu.id.opcode\[7\] cu.id.opcode\[2\] cu.id.opcode\[1\] vssd1
+ vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3702__A2 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3466__B2 cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4124__A _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5654__S _1739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5170_ mc.cl.next_data\[9\] net19 mc.count vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__mux2_1
X_4121_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__clkbuf_8
X_4052_ _1115_ _1116_ _1119_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__or4b_4
X_3003_ net72 net31 ih.gpio_interrupt_mask\[4\] vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__and3b_1
Xinput4 keypad_input[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_4954_ _1233_ cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3905_ _0350_ _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4885_ _1879_ _1880_ _1799_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3836_ _0845_ _0910_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3767_ _0841_ _0838_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__or2b_1
X_5506_ _1489_ _2125_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3698_ _0514_ _0605_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__or2_2
X_5437_ _2139_ _2225_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__nand2_1
X_5368_ _2227_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5685__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5299_ _1190_ net88 _2182_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4319_ cu.reg_file.reg_a\[3\] _1276_ _1287_ cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1
+ vccd1 _1384_ sky130_fd_sc_hd__a22o_1
XANTENNA__4645__B1 _1670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__A0 cu.reg_file.reg_c\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3620__A1 cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3620__B2 cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5373__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4879__A _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4884__A0 _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4939__A1 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3958__A _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__A2 _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3611__A1 cu.reg_file.reg_c\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3611__B2 cu.reg_file.reg_e\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4670_ ih.t.count\[12\] _1696_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4789__A _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3621_ cu.reg_file.reg_sp\[3\] _0413_ _0419_ cu.reg_file.reg_h\[3\] _0696_ vssd1
+ vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3552_ _0494_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6271_ clknet_leaf_15_clk _0253_ net175 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_3483_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[7\] vssd1 vssd1 vccd1 vccd1 _0559_
+ sky130_fd_sc_hd__o211a_1
X_5222_ _2133_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
X_5153_ cu.reg_file.reg_l\[1\] _1051_ _2088_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4104_ _0547_ _0833_ _1176_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a211o_1
X_5084_ cu.reg_file.reg_d\[2\] _2043_ _2039_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__mux2_1
X_4035_ _1099_ _1105_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5986_ clknet_leaf_28_clk _0024_ net186 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[8\] sky130_fd_sc_hd__dfrtp_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4937_ _1928_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3602__B2 cu.reg_file.reg_a\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3602__A1 cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_31 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _1863_ _1864_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3819_ cu.reg_file.reg_mem\[9\] _0640_ _0893_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_
+ sky130_fd_sc_hd__a211oi_4
X_4799_ _0310_ _0311_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5307__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5107__A1 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3669__A1 cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5291__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5043__A0 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5594__A1 _2410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5932__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3018__A ih.t.timer_max\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5379__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5624__A_N _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5034__A0 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5840_ cu.reg_file.reg_sp\[13\] _2536_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__nand2_1
X_2983_ net7 vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__inv_2
X_5771_ _2557_ _2558_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__xor2_1
X_4722_ _1732_ _1733_ _1669_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5337__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4653_ net229 _1683_ _1687_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3348__B1 _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4584_ _1511_ _1530_ _1545_ _1496_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__or4b_1
XANTENNA__3899__A1 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3604_ _0677_ _0679_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__or2_1
X_3535_ _0377_ _0602_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nor2_4
XFILLER_0_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3466_ cu.reg_file.reg_mem\[1\] _0482_ _0493_ _0495_ cu.reg_file.reg_h\[1\] vssd1
+ vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__a32o_1
X_6254_ clknet_leaf_2_clk _0236_ net155 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[10\]
+ sky130_fd_sc_hd__dfstp_2
X_5205_ net223 mc.cc.enable_edge_detector.prev_data _2122_ _2123_ vssd1 vssd1 vccd1
+ vccd1 _0099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4966__B cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6185_ clknet_leaf_35_clk _0218_ net162 vssd1 vssd1 vccd1 vccd1 ih.interrupt_source\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3397_ net149 _0469_ _0453_ _0472_ _0293_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__a41o_4
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5136_ _2077_ cu.reg_file.reg_h\[4\] _2069_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__mux2_1
X_5067_ _2031_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_1
X_4018_ _0776_ _0801_ _1091_ _0768_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5025__A0 _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__A2 _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5576__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5576__B2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5969_ _2694_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4921__S _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5053__A _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3275__C1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3814__A1 cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5228__A _1415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _0373_ _0374_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3251_ _0324_ _0325_ _2897_ _2909_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__a2111o_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ cu.id.cb_opcode_z\[0\] cu.id.cb_opcode_z\[1\] cu.id.cb_opcode_z\[2\] vssd1
+ vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__and3b_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6209__D net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3805__A1 cu.reg_file.reg_a\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5823_ cu.reg_file.reg_sp\[11\] _2536_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2966_ _2698_ mc.rw.state\[1\] mc.rw.state\[0\] vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__and3_1
X_5754_ _2530_ _2543_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__xnor2_1
X_4705_ _1722_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[23\] sky130_fd_sc_hd__clkbuf_1
X_5685_ net17 _1650_ _2488_ _2495_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__a31o_1
X_4636_ _1675_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5730__A1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4533__A2 _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4567_ _2701_ _1618_ _1353_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__a21o_1
X_6306_ clknet_leaf_9_clk _0288_ net165 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4498_ cu.reg_file.reg_b\[4\] net144 _1284_ cu.reg_file.reg_h\[4\] _1553_ vssd1 vssd1
+ vccd1 vccd1 _1554_ sky130_fd_sc_hd__a221o_1
X_3518_ _0340_ _0443_ _0336_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__a21o_1
X_6237_ clknet_leaf_24_clk ih.t.next_count\[25\] net193 vssd1 vssd1 vccd1 vccd1 ih.t.count\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_3449_ _0359_ _0386_ _2887_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ clknet_leaf_3_clk _0202_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _2034_ _2023_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__or2_1
X_6099_ clknet_leaf_9_clk _0133_ net165 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_2
XANTENNA__4049__B2 _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4217__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5549__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4221__A1 cu.reg_file.reg_e\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4221__B2 cu.reg_file.reg_l\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3015__B ih.t.timer_max\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output132_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4460__B2 _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3966__A _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5960__A1 _2410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5470_ net63 _2085_ _2294_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4421_ _1423_ _1437_ _1456_ _1474_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__or4_1
XANTENNA__4797__A _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5392__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6243__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4352_ _1356_ _1404_ _1402_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4283_ _1335_ _1349_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nand2_1
X_3303_ _0378_ _0309_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__and2_2
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4279__A1 cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6022_ clknet_leaf_31_clk _0060_ net183 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _2923_ _2874_ _0309_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__and3_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4279__B2 cu.reg_file.reg_e\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ cu.id.alu_opcode\[1\] vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__buf_4
X_3096_ ih.t.count\[5\] _2833_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout163_A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4451__A1 cu.reg_file.reg_b\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3006__A2 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5400__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3998_ _0531_ _1071_ _1040_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__mux2_1
X_5806_ _2589_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_5737_ _2518_ mc.cl.next_data\[7\] _2111_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ ih.gpio_interrupt_mask\[7\] _2326_ _2480_ _2125_ _2327_ vssd1 vssd1 vccd1
+ vccd1 _2481_ sky130_fd_sc_hd__a221o_1
X_4619_ _1650_ _1657_ _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__mux2_1
X_5599_ net104 _2205_ _2414_ _1401_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5219__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4442__A1 _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3402__C1 _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5942__A1 _2410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5506__A _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5458__A0 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5940__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output57_A net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5241__A _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4433__A1 cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4970_ _1209_ _1953_ _1794_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__mux2_1
XANTENNA__4433__B2 cu.id.imm_i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3921_ _0989_ _0994_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3852_ _0853_ _0850_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5522_ _2336_ _2341_ _2282_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3783_ cu.pc.pc_o\[12\] _0740_ _0857_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5453_ _1374_ _2278_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__or3_1
X_5384_ _2235_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4404_ cu.reg_file.reg_e\[7\] _1283_ _1285_ cu.reg_file.reg_l\[7\] _1464_ vssd1 vssd1
+ vccd1 vccd1 _1465_ sky130_fd_sc_hd__a221o_1
X_4335_ _1393_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__clkbuf_4
X_4266_ _2697_ _1333_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6005_ clknet_leaf_31_clk _0043_ net183 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3217_ cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__clkbuf_4
X_4197_ _0370_ _1261_ _1262_ _1264_ _1265_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a221o_1
X_3148_ cu.id.alu_opcode\[0\] cu.id.opcode\[0\] vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__and2_2
XANTENNA__3337__A_N _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3079_ ih.t.timer_max\[10\] _2752_ ih.t.timer_max\[11\] vssd1 vssd1 vccd1 vccd1 _2817_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5297__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5924__A1 _2391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4188__A0 cu.alu_f\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4514__A2_N _1561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5000__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3280__A1_N _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4120_ _1144_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__buf_4
X_4051_ _0570_ _0644_ _1124_ _1069_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o22a_1
XANTENNA__4103__B1 _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 keypad_input[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_4
X_3002_ net73 vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__inv_2
XANTENNA__5851__A0 cu.reg_file.reg_sp\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _2920_ cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__and2_1
XANTENNA__3614__C1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3904_ _0449_ _0971_ _0979_ _2935_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__and4b_2
XFILLER_0_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4884_ _1126_ _1874_ _1795_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3835_ _0838_ _0841_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nor2_1
X_3766_ _0838_ _0841_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__and2b_1
X_5505_ mc.cl.next_data\[0\] _2313_ _2323_ net237 vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__a22o_1
X_5436_ _2267_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3697_ _0772_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__clkbuf_4
X_5367_ _0619_ net116 _2226_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _1377_ _1379_ _1378_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__a21bo_1
X_5298_ _2186_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
X_4249_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__A1 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__A _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4879__B cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3136__A1 _2745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3304__A _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3620_ cu.reg_file.reg_d\[3\] _0415_ _0432_ cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1
+ vccd1 _0696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3551_ cu.reg_file.reg_h\[6\] _0495_ _0624_ cu.reg_file.reg_sp\[6\] _0626_ vssd1
+ vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__a221o_1
X_6270_ clknet_leaf_13_clk _0252_ net174 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3482_ _0547_ _0549_ _0552_ _0554_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__a2111o_4
X_5221_ _1192_ ih.gpio_interrupt_mask\[5\] _2127_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__mux2_1
X_5152_ _2089_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__clkbuf_1
X_4103_ _0547_ _0833_ _0824_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4627__B2 _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5083_ _1074_ _1226_ _2035_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__mux2_1
X_4034_ _0570_ _0733_ _1106_ _1107_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5985_ clknet_leaf_28_clk _0023_ net186 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _1521_ _1927_ _1814_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3602__A2 _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 programmable_gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _0373_ cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4158__A3 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ cu.reg_file.reg_b\[1\] _0426_ _0429_ cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1
+ vccd1 _0894_ sky130_fd_sc_hd__a22o_1
X_4798_ _1789_ _1796_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__mux2_1
X_3749_ cu.reg_file.reg_d\[7\] _0488_ _0741_ cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1
+ vccd1 _0825_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5419_ _1261_ net139 _2248_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3669__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5291__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5043__A1 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6180__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4554__B1 _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5704__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5034__A1 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2982_ net17 vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__inv_2
X_5770_ _2550_ _2551_ _2549_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__a21o_1
X_4721_ ih.t.count\[27\] ih.t.count\[28\] _1726_ ih.t.count\[29\] vssd1 vssd1 vccd1
+ vccd1 _1733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4652_ _1669_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput30 programmable_gpio_in[3] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3603_ cu.reg_file.reg_sp\[4\] _0539_ _0492_ cu.reg_file.reg_d\[4\] _0678_ vssd1
+ vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4312__B _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4583_ _1561_ _1626_ _1598_ _1614_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3534_ _0609_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3465_ cu.reg_file.reg_e\[1\] _0480_ _0487_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__and3_1
X_6253_ clknet_leaf_2_clk _0235_ net155 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[9\]
+ sky130_fd_sc_hd__dfstp_2
X_5204_ mc.cc.count\[1\] _2118_ _2120_ mc.cc.count\[2\] vssd1 vssd1 vccd1 vccd1 _2123_
+ sky130_fd_sc_hd__o211a_1
X_6184_ clknet_leaf_35_clk net199 net162 vssd1 vssd1 vccd1 vccd1 ih.interrupt_source\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3396_ _2918_ _0355_ _0470_ _2902_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout193_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5135_ _1213_ _1160_ _2066_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ cu.reg_file.reg_c\[5\] _1191_ _2025_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__mux2_1
XANTENNA__5273__A1 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4017_ _0770_ _0773_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5025__A1 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5968_ cu.id.imm_i\[15\] _2486_ _2686_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__mux2_1
XANTENNA__5576__A2 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4919_ _1910_ _1911_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__xor2_1
X_5899_ ih.t.timer_max\[18\] _1074_ _2654_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3511__A1 _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4067__A2 _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3814__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3750__B2 cu.reg_file.reg_sp\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3250_ _2899_ _2900_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__nand2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _2916_ _2917_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__nand2b_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3502__B2 cu.reg_file.reg_a\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5822_ _2603_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
X_5753_ _2541_ _2542_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__and2_1
X_4704_ _1720_ _1721_ _1672_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__and3b_1
XFILLER_0_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2965_ _2704_ _2699_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5684_ _2494_ _1643_ cu.reg_file.reg_mem\[9\] _1646_ vssd1 vssd1 vccd1 vccd1 _2495_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4635_ _1672_ _1673_ _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__and3_1
X_4566_ _1356_ _1614_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6305_ clknet_leaf_9_clk _0287_ net165 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3517_ cu.reg_file.reg_l\[1\] _0422_ _0592_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__a21o_1
X_4497_ cu.reg_file.reg_d\[4\] _1282_ _1286_ cu.reg_file.reg_sp\[12\] vssd1 vssd1
+ vccd1 vccd1 _1553_ sky130_fd_sc_hd__a22o_1
X_6236_ clknet_leaf_24_clk ih.t.next_count\[24\] net192 vssd1 vssd1 vccd1 vccd1 ih.t.count\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_3448_ _0372_ _0522_ _0523_ _0387_ _2918_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__a311o_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _0298_ _2923_ _2901_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or3_1
X_6167_ clknet_leaf_3_clk _0201_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _2064_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__clkbuf_1
X_6098_ clknet_leaf_9_clk _0132_ net165 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_4
X_5049_ _1260_ _1263_ _2002_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5549__A2 _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output125_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4408__A cu.reg_file.reg_l\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3312__A cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5003__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5938__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3420__B1 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4143__A _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3971__A1 _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4420_ _1440_ _1462_ _1473_ _1332_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4920__A0 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4250__D_N _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ _1306_ _1410_ _1414_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__o21a_4
X_4282_ _1332_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__xnor2_1
X_3302_ _2892_ _2894_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__and2b_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ clknet_leaf_31_clk _0059_ net183 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3233_ cu.id.opcode\[1\] cu.id.opcode\[6\] cu.id.opcode\[7\] cu.id.opcode\[2\] vssd1
+ vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__and4b_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5421__B _1372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3164_ _2899_ _2875_ _2876_ _2900_ vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__or4b_4
X_3095_ ih.t.timer_max\[5\] _2749_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout156_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5400__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3997_ _0588_ _1044_ _1061_ _0610_ _1045_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__o221a_1
XANTENNA__5149__A _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5805_ cu.reg_file.reg_sp\[8\] _2588_ _2539_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__mux2_1
X_5736_ net24 _2519_ _2528_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4053__A _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5667_ mc.cl.next_data\[7\] _2313_ net142 _2479_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__a22o_1
XANTENNA__4988__A cu.pc.pc_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4618_ _1660_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3892__A _0379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5598_ net88 _1330_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__or2_1
X_4549_ _1581_ _1601_ _1588_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__nand3_1
X_6219_ clknet_leaf_14_clk ih.t.next_count\[7\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5612__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2971__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3134__B_N _2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5155__A0 cu.reg_file.reg_l\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5458__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5630__A1 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3977__A _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _0995_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3696__B _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3851_ _0866_ _0925_ _0926_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__o21a_1
XANTENNA__5394__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3782_ cu.reg_file.reg_b\[4\] _0743_ _0624_ cu.reg_file.reg_sp\[12\] vssd1 vssd1
+ vccd1 vccd1 _0858_ sky130_fd_sc_hd__a22o_1
X_5521_ _2337_ _2338_ _2339_ _2340_ _1369_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5697__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5452_ net71 _1638_ _2279_ net70 vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__a22o_1
X_5383_ _1369_ _2191_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__nor2_1
X_4403_ cu.reg_file.reg_a\[7\] _1276_ _1287_ cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1
+ vccd1 _1464_ sky130_fd_sc_hd__a22o_1
X_4334_ _1397_ _1394_ _1383_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__a21o_1
XANTENNA__3217__A cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4265_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__clkbuf_4
X_6004_ clknet_leaf_20_clk _0042_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3216_ _2896_ _2952_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__nand2_2
X_4196_ cu.alu_f\[7\] _1027_ _1184_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__and3_1
X_3147_ cu.id.alu_opcode\[3\] vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ _2754_ _2814_ ih.t.count\[12\] vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5621__B2 _2435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5621__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3887__A _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3632__B1 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4188__A1 _1256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3935__A1 _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5719_ _2514_ _2519_ _2520_ _2518_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5688__B2 _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4112__A1 _1027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__A1 _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4179__A1 _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4050_ _1120_ _1096_ _1097_ _0754_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__o221a_1
X_3001_ net74 vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__inv_2
Xinput6 keypad_input[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5603__A1 ih.t.timer_max\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5398__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _1213_ _1941_ _1795_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__mux2_1
X_4883_ _1877_ _1878_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__xor2_1
X_3903_ _0308_ _0525_ _0977_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__and4b_1
XANTENNA__5367__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3834_ _0856_ _0908_ _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3765_ cu.reg_file.reg_mem\[14\] _0640_ _0839_ _0840_ vssd1 vssd1 vccd1 vccd1 _0841_
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5504_ _1374_ _1625_ _1630_ _1489_ _1417_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__a2111oi_1
X_3696_ _0512_ _0528_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5435_ _2022_ net72 _2266_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__mux2_1
XANTENNA__4342__A1 cu.reg_file.reg_a\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5366_ net141 _2225_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__nand2_8
XANTENNA__4342__B2 cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4317_ _1370_ _1375_ _1381_ _1382_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__a22o_1
X_5297_ _1188_ net87 _2182_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__mux2_1
X_4248_ _1309_ _1311_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nor2b_2
X_4179_ _0574_ _0545_ _0447_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3605__B1 _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5358__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6315__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3136__A2 _2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5800__A cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5011__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3320__A _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5946__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4135__B _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3550_ cu.reg_file.reg_d\[6\] _0492_ _0625_ cu.alu_f\[6\] vssd1 vssd1 vccd1 vccd1
+ _0626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5220_ _2132_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3481_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5151_ cu.reg_file.reg_l\[0\] _2085_ _2088_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__mux2_1
X_5082_ _2042_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
X_4102_ _0829_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__xnor2_1
X_4033_ _0822_ _0632_ _0566_ _0531_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ clknet_leaf_29_clk _0022_ net188 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[6\] sky130_fd_sc_hd__dfrtp_4
X_4935_ _1917_ _1926_ _1808_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_22 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _0373_ cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_11 programmable_gpio_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4797_ _1798_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3817_ cu.reg_file.reg_sp\[9\] _0636_ _0748_ cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1
+ vccd1 _0893_ sky130_fd_sc_hd__a22o_1
X_3748_ _0384_ _0392_ _0400_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__and3_2
XFILLER_0_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3679_ _0684_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__inv_2
X_5418_ _2255_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
X_5349_ _2216_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4935__S _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3287__D1 _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4554__B2 cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5006__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3817__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2981_ _2715_ ih.ih.ih.prev_data\[6\] _2716_ ih.ih.ih.prev_data\[12\] _2719_ vssd1
+ vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4720_ ih.t.count\[28\] ih.t.count\[29\] _1729_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_41_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4651_ ih.t.count\[6\] _1683_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 memory_data_in[2] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
X_3602_ cu.pc.pc_o\[4\] _0501_ _0499_ cu.reg_file.reg_a\[4\] _0504_ vssd1 vssd1 vccd1
+ vccd1 _0678_ sky130_fd_sc_hd__a221o_1
Xinput31 programmable_gpio_in[4] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_2
X_4582_ _1579_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__inv_2
X_3533_ _0548_ _0393_ _0529_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3464_ cu.reg_file.reg_a\[1\] _0499_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__and2_1
X_6252_ clknet_leaf_1_clk _0234_ net155 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[8\]
+ sky130_fd_sc_hd__dfstp_2
X_5203_ mc.cc.count\[2\] mc.cc.count\[1\] _2118_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__nor3_1
X_6183_ clknet_leaf_22_clk _0216_ net190 vssd1 vssd1 vccd1 vccd1 mc.count sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3395_ _2878_ _0402_ _0301_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__a21o_1
X_5134_ _2076_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5440__A _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5065_ _2030_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3808__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4016_ _1073_ _1089_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4481__B1 _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5967_ _2693_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4918_ _1899_ _1902_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _2656_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4849_ _1840_ _1847_ _1809_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__mux2_1
XANTENNA__4536__A1 cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5543__A_N _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3983__C1 _1027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4413__B _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3750__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _2899_ _2900_ _2875_ _2876_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__and4b_2
XFILLER_0_28_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5821_ cu.reg_file.reg_sp\[10\] _2602_ _2539_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__mux2_1
X_2964_ _2695_ mc.rw.state\[0\] vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__and2_1
XANTENNA__4604__A _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5752_ cu.reg_file.reg_sp\[2\] _2534_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ ih.t.count\[21\] ih.t.count\[22\] _1714_ ih.t.count\[23\] vssd1 vssd1 vccd1
+ vccd1 _1721_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_14_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5683_ mc.cl.next_data\[9\] _2359_ _2490_ _2493_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__o2bb2a_1
X_4634_ ih.t.count\[0\] ih.t.count\[1\] vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__or2_1
XANTENNA__4518__B2 cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4565_ _1567_ _1579_ _1598_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__or3b_1
X_6304_ clknet_leaf_9_clk _0286_ net165 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[9\] sky130_fd_sc_hd__dfrtp_4
X_3516_ cu.reg_file.reg_b\[1\] _0432_ _0433_ cu.reg_file.reg_a\[1\] vssd1 vssd1 vccd1
+ vccd1 _0592_ sky130_fd_sc_hd__a22o_1
X_4496_ _1351_ _1550_ _1551_ _1371_ _1552_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__a221o_1
XFILLER_0_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6235_ clknet_leaf_23_clk ih.t.next_count\[23\] net179 vssd1 vssd1 vccd1 vccd1 ih.t.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3447_ _0373_ cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _0379_ _0450_ _0451_ _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__or4b_2
X_6166_ clknet_leaf_3_clk _0200_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ clknet_leaf_27_clk _0131_ net195 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ cu.reg_file.reg_e\[7\] _1260_ _2056_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__mux2_1
X_5048_ _2019_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4206__B1 _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5954__A0 cu.id.imm_i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3312__B _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output118_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5954__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3420__B2 cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3420__A1 cu.reg_file.reg_sp\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5173__A1 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ cu.reg_file.reg_c\[4\] _1313_ _1411_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3301_ _0371_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__nor2_1
X_4281_ _1340_ _1341_ _1347_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__o21a_4
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ clknet_leaf_20_clk _0058_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _2902_ _0304_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__o21ai_2
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__A1 cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3163_ cu.id.opcode\[1\] vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__buf_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3094_ _2750_ _2830_ ih.t.count\[6\] vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5421__C _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5936__A0 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5804_ _1622_ _2587_ _2545_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3996_ _0570_ _0759_ _1068_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__o22a_1
X_5735_ _2518_ mc.cl.next_data\[6\] _2111_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4053__B _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5666_ _1665_ _2477_ _2478_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__o21a_1
X_4617_ _0315_ _1658_ _1659_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5597_ net96 _2194_ _2412_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4548_ _1581_ _1588_ _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__a21o_1
X_4479_ _1382_ _1532_ _1533_ _1536_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__a31o_1
XFILLER_0_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6218_ clknet_leaf_14_clk ih.t.next_count\[6\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6149_ clknet_leaf_8_clk _0183_ net172 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4427__B1 _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3650__A1 cu.reg_file.reg_c\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5975__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3953__A2 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5155__A1 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5014__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5630__A2 _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _0861_ _0864_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__or2b_1
XANTENNA__5394__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3781_ cu.reg_file.reg_d\[4\] _0488_ _0741_ cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1
+ vccd1 _0857_ sky130_fd_sc_hd__a22o_1
XANTENNA__4197__A2 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5520_ net28 net30 net27 net29 _1354_ _1330_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5451_ _1335_ _1372_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5382_ _2234_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5697__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4402_ _1333_ _1462_ _1457_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__o21a_1
X_4333_ _1395_ _1397_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4264_ _1331_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__clkbuf_4
X_3215_ _2938_ _2932_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6003_ clknet_leaf_5_clk _0041_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4195_ _0516_ _1260_ _1263_ _1027_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__a22o_1
X_3146_ cu.id.alu_opcode\[1\] vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__inv_2
X_3077_ ih.t.count\[12\] _2754_ _2814_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5621__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3632__A1 cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5604__A_N _1400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5718_ _2351_ _2514_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__nor2_1
X_3979_ _0372_ _0371_ _0774_ _1019_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o2111a_1
XANTENNA__5594__S _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4511__B _1561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5649_ _2169_ _2455_ _2462_ _2136_ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__o211a_1
XANTENNA__4112__A2 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__A2 _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2982__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3623__B2 cu.reg_file.reg_a\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3623__A1 cu.reg_file.reg_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5517__B _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5009__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4887__A0 cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output62_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3000_ net71 net30 ih.gpio_interrupt_mask\[3\] vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__and3b_1
Xinput7 keypad_input[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_4
X_4951_ _1939_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__nor2_1
XANTENNA__3614__A1 cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3614__B2 cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4882_ _1863_ _1866_ _1864_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3902_ _2886_ _0965_ _0521_ _0359_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5367__A1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3833_ _0850_ _0853_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3764_ cu.reg_file.reg_b\[6\] _0426_ _0429_ cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1
+ vccd1 _0840_ sky130_fd_sc_hd__a22o_1
X_5503_ _1661_ _2318_ _2322_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3695_ _0768_ _0770_ _0753_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__or3b_1
X_5434_ _2139_ _2147_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__nand2_1
XANTENNA__3228__A _2936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5443__A _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5365_ _2224_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4316_ _1351_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__clkbuf_4
X_5296_ _2185_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__clkbuf_1
X_4247_ _1314_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__buf_2
X_4178_ _1246_ _1247_ _0600_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__mux2_1
X_3129_ ih.t.count\[30\] _2866_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__nor2_1
XANTENNA__5055__B1 _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4506__B _1561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5358__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__C _1269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5618__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2977__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5046__A0 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5597__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output100_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3320__B _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5962__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3480_ _0550_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__nand2_1
XANTENNA__5521__B2 _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6025__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5150_ _2087_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__clkbuf_4
X_5081_ cu.reg_file.reg_d\[1\] _2041_ _2039_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4101_ _0918_ _0948_ _1172_ _1174_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5285__A0 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4032_ alu.Cin _0554_ _0556_ _0509_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5037__A0 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ clknet_leaf_28_clk _0021_ net186 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[5\] sky130_fd_sc_hd__dfrtp_4
X_4934_ _1924_ _1925_ _1798_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4260__A1 cu.reg_file.reg_c\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _1860_ _1861_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_34 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4796_ _2948_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__nand2_8
XFILLER_0_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3816_ cu.id.imm_i\[9\] _0739_ _0891_ _0653_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__a22oi_4
X_3747_ _0574_ _0558_ _0822_ _0566_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3678_ _0645_ _0722_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5417_ _1194_ net138 _2248_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__mux2_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ss6[6] sky130_fd_sc_hd__buf_2
XANTENNA__5512__B2 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5512__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5348_ _0619_ net108 _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__mux2_1
X_5279_ net80 _1189_ _2170_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__mux2_1
XANTENNA__5028__B1 _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5579__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5579__B2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5503__A1 _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3817__A1 cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3817__B2 cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2980_ _2717_ ih.ih.ih.prev_data\[4\] _2718_ ih.ih.ih.prev_data\[13\] vssd1 vssd1
+ vccd1 vccd1 _2719_ sky130_fd_sc_hd__o22a_1
XANTENNA__3450__C1 _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4650_ _1685_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4162__A _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput21 memory_data_in[3] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
Xinput10 keypad_input[2] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_2
X_3601_ cu.reg_file.reg_b\[4\] _0502_ _0494_ cu.reg_file.reg_mem\[4\] _0676_ vssd1
+ vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__a221o_1
Xinput32 programmable_gpio_in[5] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
X_4581_ _1329_ _1372_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3532_ _0574_ _0604_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__o21ai_1
X_3463_ _0480_ _0493_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__and2_2
X_6251_ clknet_leaf_1_clk _0233_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_5202_ net228 _2118_ _2121_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a21o_1
X_6182_ clknet_leaf_7_clk _0215_ net172 vssd1 vssd1 vccd1 vccd1 ih.input_handler_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3394_ _0378_ _0309_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__nand2_1
X_5133_ _2075_ cu.reg_file.reg_h\[3\] _2069_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5064_ cu.reg_file.reg_c\[4\] _1189_ _2025_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__mux2_1
XANTENNA__5440__B _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4015_ _1081_ _1082_ _1085_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout179_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4481__A1 cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4481__B2 cu.reg_file.reg_h\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5966_ cu.id.imm_i\[14\] _2467_ _2686_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__mux2_1
X_5897_ ih.t.timer_max\[17\] _1051_ _2654_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__mux2_1
X_4917_ _2920_ cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__xor2_1
XANTENNA__5168__A _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4848_ _1845_ _1846_ _1799_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3992__B1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _1775_ _1779_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4946__S _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2990__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5724__A1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4527__A2 _1561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5017__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5660__B1 _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5820_ _1226_ _2601_ _2545_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2963_ _2703_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_5751_ cu.reg_file.reg_sp\[2\] _2534_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__nand2_1
X_4702_ ih.t.count\[22\] ih.t.count\[23\] _1717_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5682_ ih.t.timer_max\[25\] _2151_ _2320_ ih.t.timer_max\[9\] vssd1 vssd1 vccd1 vccd1
+ _2493_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ ih.t.count\[0\] ih.t.count\[1\] vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4564_ _1599_ _1602_ _1615_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__nand3_1
XANTENNA__6040__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6303_ clknet_leaf_7_clk _0285_ net170 vssd1 vssd1 vccd1 vccd1 cu.id.imm_i\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3515_ cu.reg_file.reg_sp\[1\] _0413_ _0419_ cu.reg_file.reg_h\[1\] _0590_ vssd1
+ vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__a221o_1
X_6234_ clknet_leaf_17_clk ih.t.next_count\[22\] net179 vssd1 vssd1 vccd1 vccd1 ih.t.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_4495_ _1402_ _1545_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3446_ _0373_ cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nand2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3377_ _0452_ _0303_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__nor2_1
X_6165_ clknet_leaf_0_clk _0199_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ clknet_leaf_10_clk _0130_ net166 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_4
X_5116_ _2063_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__clkbuf_1
X_5047_ cu.reg_file.reg_b\[6\] _2018_ _2006_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5954__A1 _2350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5949_ _2683_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3414__C1 cu.reg_file.reg_l\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5706__B2 ih.t.timer_max\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3193__A1 _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5890__A0 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2985__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__A1 cu.reg_file.reg_b\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__B2 cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3956__B1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output92_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _0372_ _2921_ _0375_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4280_ cu.reg_file.reg_c\[1\] _1313_ _1342_ _1346_ vssd1 vssd1 vccd1 vccd1 _1347_
+ sky130_fd_sc_hd__a211o_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _2897_ _2917_ _0305_ _0306_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o2bb2a_2
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4133__B1 _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3162_ cu.id.opcode\[2\] vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__buf_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__A2 _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3093_ ih.t.count\[6\] _2750_ _2830_ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4615__A _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5803_ _2585_ _2586_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3995_ _0620_ _0824_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3947__B1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5936__A1 _2350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5734_ net23 _2519_ _2527_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a21o_1
X_5665_ ih.t.timer_max\[23\] _2150_ _2319_ ih.t.timer_max\[7\] _1660_ vssd1 vssd1
+ vccd1 vccd1 _2478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4616_ _2923_ _2903_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__or2_1
X_5596_ net128 _2236_ _2247_ net136 vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5880__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4547_ _1599_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__nand2_1
Xmax_cap151 net243 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xmax_cap140 _2873_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_1
X_4478_ _1530_ _1534_ _1535_ _1356_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6217_ clknet_leaf_14_clk ih.t.next_count\[5\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3429_ cu.pc.pc_o\[0\] _0501_ _0502_ cu.reg_file.reg_b\[0\] _0504_ vssd1 vssd1 vccd1
+ vccd1 _0505_ sky130_fd_sc_hd__a221o_1
X_6148_ clknet_leaf_20_clk _0182_ net182 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ clknet_leaf_23_clk _0113_ net192 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4427__B2 cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4427__A1 cu.reg_file.reg_b\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4244__B _1309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5863__A0 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4418__A1 _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output130_A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ _0854_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5450_ net68 _2277_ _2179_ net69 vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4401_ _1455_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__inv_2
X_5381_ _1261_ net123 _2226_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4332_ _1396_ _1393_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ mc.rw.state\[2\] _2699_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__and2_1
XANTENNA__5713__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6002_ clknet_leaf_20_clk _0040_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_b\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3214_ _2882_ _2906_ _2945_ _2948_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__o311a_4
XANTENNA__4329__B _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4194_ _0516_ _1175_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__nor2_4
X_3145_ _2874_ _2881_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__nor2_1
XANTENNA__4409__A1 cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4409__B2 cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3076_ ih.t.timer_max\[12\] _2753_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5909__A1 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3978_ _1021_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__inv_2
X_5717_ _2518_ _2351_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__nor2_4
XANTENNA__3396__A1 _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5648_ ih.gpio_interrupt_mask\[6\] _2326_ _2461_ _2125_ _2327_ vssd1 vssd1 vccd1
+ vccd1 _2462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5579_ net103 _2205_ _2395_ _1401_ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3424__A cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5845__A0 cu.reg_file.reg_sp\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5517__C _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5025__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5836__A0 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output55_A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 keypad_input[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_2
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5064__A1 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4950_ cu.pc.pc_o\[12\] _1929_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__nor2_1
XANTENNA__3614__A2 _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4881_ _1875_ _1876_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__or2b_1
X_3901_ _0361_ _0332_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3832_ _0866_ _0906_ _0907_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4575__B1 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5502_ ih.t.timer_max\[0\] _2320_ _2321_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3763_ cu.reg_file.reg_sp\[14\] _0636_ _0748_ cu.reg_file.reg_h\[6\] vssd1 vssd1
+ vccd1 vccd1 _0839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _0769_ _0734_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__xnor2_2
X_5433_ _2265_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5364_ _1374_ _2179_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__and2_1
XANTENNA__5443__B _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4315_ _1377_ _1380_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3550__A1 cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5295_ _1075_ net86 _2182_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__mux2_1
XANTENNA__3550__B2 cu.alu_f\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4246_ _1309_ _1311_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__nor2_2
X_4177_ _0663_ _0681_ _1060_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__mux2_1
X_3128_ _2766_ _2865_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__nor2_1
XANTENNA__5055__A1 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3059_ ih.t.count\[19\] _2796_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__xnor2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5618__B _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3369__A1 cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3369__B2 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5046__A1 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5597__A2 _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4309__B1 _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4100_ _0960_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__nand2_1
X_5080_ _1051_ _1623_ _2035_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__mux2_1
XANTENNA__5285__A1 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _1102_ _1103_ _1104_ _0566_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5037__A1 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5982_ clknet_leaf_28_clk _0020_ net186 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4933_ _1226_ _1917_ _1794_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4864_ cu.pc.pc_o\[4\] _1838_ cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_35 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _0986_ _1005_ _1786_ _0983_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_24 _0651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3815_ cu.reg_file.reg_a\[1\] _0625_ _0628_ cu.reg_file.reg_mem\[9\] _0890_ vssd1
+ vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__a221o_1
X_3746_ _0550_ _0820_ _0821_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__a21o_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3771__B2 cu.reg_file.reg_sp\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3771__A1 cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5416_ _2254_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3677_ _0737_ _0752_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__xor2_1
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ss5[4] sky130_fd_sc_hd__clkbuf_4
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ss6[7] sky130_fd_sc_hd__clkbuf_4
X_5347_ _2147_ net141 vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__nand2_8
X_5278_ _2174_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4229_ _1296_ _1294_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__nor2_2
XANTENNA__5028__A1 _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5579__A2 _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3762__A1 cu.id.imm_i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5364__A _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2988__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3514__B2 cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5303__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4162__B _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput11 keypad_input[3] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 memory_data_in[4] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_2
X_4580_ _2702_ _1261_ _1263_ _2697_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__a22o_1
X_3600_ cu.reg_file.reg_h\[4\] _0495_ _0498_ cu.alu_f\[4\] vssd1 vssd1 vccd1 vccd1
+ _0676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3531_ _0603_ _0606_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__or2_2
Xinput33 programmable_gpio_in[6] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3753__A1 cu.id.imm_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3462_ cu.reg_file.reg_d\[1\] _0492_ _0498_ cu.alu_f\[1\] vssd1 vssd1 vccd1 vccd1
+ _0538_ sky130_fd_sc_hd__a22o_1
X_6250_ clknet_leaf_1_clk _0232_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_5201_ mc.cc.count\[1\] _2118_ _2120_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__o21ai_1
X_6181_ clknet_leaf_25_clk _0214_ vssd1 vssd1 vccd1 vccd1 mc.cl.cmp_o sky130_fd_sc_hd__dfxtp_1
X_3393_ _0312_ _0449_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__nor2_4
XANTENNA__3505__A1 cu.reg_file.reg_l\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5132_ _1222_ _1089_ _2066_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__mux2_1
XANTENNA__4618__A _1660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5063_ _2029_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4466__C1 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3808__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4014_ _0558_ _0681_ _0822_ _1040_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5449__A _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5965_ _2692_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5896_ _2655_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
X_4916_ _1907_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__nor2_1
X_4847_ _1089_ _1840_ _1795_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__mux2_1
X_4778_ net140 _1783_ net203 vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3729_ _0755_ _0787_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3135__C _2870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5249__A1 _2155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4962__S _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5488__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5488__B2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4160__A1 _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5660__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5660__B2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5968__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2962_ _2697_ _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__or2_1
X_5750_ _2540_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
X_4701_ net219 _1717_ _1719_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[22\] sky130_fd_sc_hd__a21oi_1
X_5681_ net16 _1650_ _2488_ _2492_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a31o_1
X_4632_ _1669_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4923__A0 cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4563_ _1599_ _1602_ _1615_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4494_ _1535_ _1545_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6302_ clknet_leaf_36_clk _0284_ net161 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_x\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3514_ cu.reg_file.reg_mem\[1\] _0418_ _0415_ cu.reg_file.reg_d\[1\] vssd1 vssd1
+ vccd1 vccd1 _0590_ sky130_fd_sc_hd__a22o_1
X_6233_ clknet_leaf_17_clk ih.t.next_count\[21\] net179 vssd1 vssd1 vccd1 vccd1 ih.t.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3445_ _2936_ _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__nor2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _2884_ _2885_ _2941_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__and3_1
X_6164_ clknet_leaf_41_clk _0198_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__B _1372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6095_ clknet_leaf_10_clk _0129_ net166 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
X_5115_ cu.reg_file.reg_e\[6\] _1193_ _2056_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5046_ _1193_ _1624_ _2002_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__mux2_1
XANTENNA__5878__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5651__B2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5651__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5948_ _0387_ _2467_ _2666_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5879_ _2646_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4530__B _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4390__A1 cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4390__B2 _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5536__B _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5552__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _2892_ _2899_ _2900_ _2923_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__or4bb_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _2893_ _2897_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__nand2_1
XANTENNA__4168__A _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3092_ ih.t.timer_max\[5\] _2749_ ih.t.timer_max\[6\] vssd1 vssd1 vccd1 vccd1 _2830_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5802_ _2576_ _2579_ _2577_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3994_ _0918_ _0760_ _1065_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__a2bb2o_1
X_5733_ _2518_ mc.cl.next_data\[5\] _2111_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5664_ _1400_ _2476_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__and2b_1
X_4615_ _0350_ _2940_ _0379_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__or3_2
X_5595_ _2411_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4546_ _1333_ _1598_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap141 _2181_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4477_ _1517_ _1530_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__nand2_1
X_6216_ clknet_leaf_14_clk ih.t.next_count\[4\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_3428_ _2948_ _0501_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__a21bo_2
X_6147_ clknet_leaf_31_clk _0181_ net183 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_4
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _2940_ _2942_ _0379_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__nor3_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ clknet_leaf_23_clk _0112_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[26\]
+ sky130_fd_sc_hd__dfrtp_2
X_5029_ cu.reg_file.reg_b\[0\] _2003_ _2006_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__mux2_1
XANTENNA__4525__B _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5388__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4244__C _1311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3938__A1 alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4363__A1 cu.reg_file.reg_e\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5560__B1 _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4363__B2 cu.reg_file.reg_l\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2996__A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5312__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5984__RESET_B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5863__A1 ih.t.timer_max\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output123_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5379__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ _1382_ _1457_ _1458_ _1461_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__a31o_2
XFILLER_0_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5380_ _2233_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3343__C_N _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4331_ _1376_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4262_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__buf_4
XANTENNA__5303__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3213_ _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__buf_4
X_6001_ clknet_leaf_3_clk _0039_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4193_ _1184_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__inv_2
XANTENNA__5606__A1 _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3144_ _2877_ _2880_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__and2_1
XANTENNA__4409__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3075_ ih.t.count\[13\] _2812_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3617__B1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3977_ _1051_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4042__B1 _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5716_ mc.count vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__buf_2
XANTENNA__5457__A _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5647_ mc.cl.next_data\[6\] _2313_ net142 _2460_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__a22o_1
X_5578_ net87 _1330_ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__or2_1
X_4529_ _1580_ _1581_ _1582_ _1334_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__a31oi_1
XANTENNA__3553__C1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3705__A _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2997__A_N net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4033__B1 _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5781__A0 cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 keypad_input[1] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
XANTENNA_output48_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5041__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4880_ _0387_ cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__nand2_1
X_3900_ _0321_ _0970_ _0972_ _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__or4_4
XFILLER_0_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3831_ _0861_ _0864_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nor2_1
XANTENNA__5772__A0 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4575__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3762_ cu.id.imm_i\[14\] _0739_ _0837_ _0653_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__a22oi_4
X_5501_ ih.t.enable _2257_ _2150_ ih.t.timer_max\[16\] _1660_ vssd1 vssd1 vccd1 vccd1
+ _2321_ sky130_fd_sc_hd__a221o_1
XANTENNA__4575__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3693_ _0645_ _0722_ _0735_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5432_ _2022_ net71 _2264_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__mux2_1
XANTENNA__4327__A1 cu.reg_file.reg_c\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5363_ _2223_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__clkbuf_1
X_4314_ _1378_ _1379_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__nand2_1
XANTENNA__3550__A2 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5294_ _2184_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4245_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__clkbuf_4
X_4176_ _0566_ _0632_ _1060_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__mux2_1
X_3127_ ih.t.timer_max\[30\] _2765_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__and2_1
X_3058_ ih.t.timer_max\[19\] _2758_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__xor2_1
XANTENNA__5886__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3435__A alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5126__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4266__A _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4557__A1 cu.pc.pc_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _0599_ _0603_ _1101_ _0729_ _0606_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__a32o_1
X_5981_ clknet_leaf_28_clk _0019_ net187 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4904__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4932_ _1920_ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6034__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4863_ cu.pc.pc_o\[5\] cu.pc.pc_o\[4\] _1838_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__and3_1
XANTENNA_14 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4794_ _0617_ _1788_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3814_ cu.pc.pc_o\[9\] _0740_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__a21o_1
X_3745_ _0614_ _0573_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3771__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5415_ _1192_ net137 _2248_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__mux2_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ss4[2] sky130_fd_sc_hd__clkbuf_4
X_3676_ _0747_ _0751_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__xor2_4
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ss7[0] sky130_fd_sc_hd__clkbuf_4
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ss5[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5346_ _2214_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5277_ net79 _1187_ _2170_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__mux2_1
X_4228_ _1271_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__inv_2
X_4159_ _0954_ _0778_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4539__A1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4162__C _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 keypad_input[4] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_2
Xinput23 memory_data_in[5] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
X_3530_ _0519_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__nor2_2
Xinput34 programmable_gpio_in[7] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
X_3461_ cu.reg_file.reg_c\[1\] _0485_ _0533_ _0535_ _0536_ vssd1 vssd1 vccd1 vccd1
+ _0537_ sky130_fd_sc_hd__a2111o_1
X_5200_ mc.cc.enable_edge_detector.prev_data _2708_ vssd1 vssd1 vccd1 vccd1 _2120_
+ sky130_fd_sc_hd__or2_1
X_6180_ clknet_leaf_36_clk _0000_ net161 vssd1 vssd1 vccd1 vccd1 ih.interrupt_source\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3392_ _0465_ net149 _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__nor3_2
X_5131_ _2074_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__clkbuf_1
X_5062_ cu.reg_file.reg_c\[3\] _1187_ _2025_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__mux2_1
XANTENNA__6286__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4013_ _0607_ _1086_ _0694_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__o21a_1
XANTENNA__3269__A1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5966__A0 cu.id.imm_i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5449__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5964_ cu.id.imm_i\[13\] _2448_ _2686_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5895_ ih.t.timer_max\[16\] _0618_ _2654_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__mux2_1
X_4915_ cu.pc.pc_o\[9\] _1894_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4846_ _1843_ _1844_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4777_ net200 _1782_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3728_ _0664_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__xnor2_1
X_3659_ _0632_ _0643_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5329_ _2204_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4202__C_N _1269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4339__A_N _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3432__A1 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5314__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5645__C1 _1660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5948__A0 _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3671__A1 cu.id.imm_i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2961_ _2698_ _2699_ _2701_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__a21o_4
XFILLER_0_60_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ ih.t.count\[22\] _1717_ _1670_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__o21ai_1
X_5680_ _2491_ _1643_ cu.reg_file.reg_mem\[8\] _2111_ vssd1 vssd1 vccd1 vccd1 _2492_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4631_ _1671_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[0\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__5176__A1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4562_ _1396_ _1614_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4493_ _1548_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6301_ clknet_leaf_38_clk _0283_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3513_ cu.reg_file.reg_c\[1\] _0427_ _0430_ cu.reg_file.reg_e\[1\] vssd1 vssd1 vccd1
+ vccd1 _0589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6232_ clknet_leaf_17_clk ih.t.next_count\[20\] net179 vssd1 vssd1 vccd1 vccd1 ih.t.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_6_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3444_ _2886_ _0378_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nand2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ clknet_leaf_10_clk _0197_ net166 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_2
X_3375_ _2878_ _0301_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nor2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ clknet_leaf_28_clk _0128_ net186 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_4
X_5114_ _2062_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__clkbuf_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _2017_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout184_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5947_ _2682_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
X_5878_ _2022_ ih.t.timer_max\[0\] _2645_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__mux2_1
XANTENNA__5167__A1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4829_ _0341_ cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4390__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4973__S _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4850__A0 cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4381__A2 _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5044__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _2894_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__inv_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4168__B _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3091_ ih.t.count\[7\] _2828_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__xnor2_1
Xhold1 ih.ip_ed.prev_data vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4615__C _0379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5801_ _2583_ _2584_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__nand2_1
X_5732_ net22 _2519_ _2526_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__a21o_1
X_3993_ _1033_ _1066_ _0806_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5663_ ih.t.timer_max\[23\] _2204_ _2314_ ih.t.timer_max\[7\] _2475_ vssd1 vssd1
+ vccd1 vccd1 _2476_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4614_ _1656_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5594_ cu.reg_file.reg_mem\[3\] _2410_ _2351_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4545_ _1333_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__or2_1
Xmax_cap142 net237 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4476_ _1356_ _1517_ _1402_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6215_ clknet_leaf_14_clk ih.t.next_count\[3\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3427_ _2913_ _2952_ _0307_ _0293_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__a31o_1
XANTENNA__3263__A _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6146_ clknet_leaf_11_clk _0180_ net167 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ cu.reg_file.reg_b\[0\] _0432_ _0433_ cu.reg_file.reg_a\[0\] vssd1 vssd1 vccd1
+ vccd1 _0434_ sky130_fd_sc_hd__a22o_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6077_ clknet_leaf_23_clk _0111_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_3289_ _2940_ _2953_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__o21bai_1
X_5028_ _2002_ _2005_ _2951_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__o21a_4
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5388__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5129__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4348__C1 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5560__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5560__B2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5312__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output116_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5379__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4587__C1 _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5000__A0 cu.reg_file.reg_a\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5551__A1 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5551__B2 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4330_ _1383_ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4261_ _1291_ _1307_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__o21bai_4
XANTENNA__5303__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3314__B1 _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3212_ cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__inv_2
X_6000_ clknet_leaf_4_clk _0038_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_4192_ _1260_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__buf_4
X_3143_ _2878_ _2879_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__or2_2
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3074_ ih.t.timer_max\[13\] _2754_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__xor2_1
XANTENNA__4814__A0 _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3976_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5457__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5715_ _2517_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5646_ _1665_ _2458_ _2459_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5542__A1 ih.t.timer_max\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5542__B2 ih.t.timer_max\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5577_ net95 _2194_ _2393_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4528_ _1580_ _1581_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__a21o_1
X_4459_ _1356_ _1501_ _1402_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__o21a_1
XANTENNA__4502__C1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6129_ clknet_leaf_21_clk _0163_ net182 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XANTENNA__4817__A _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5058__A0 cu.reg_file.reg_c\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5383__A _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5297__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5322__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__A0 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4272__A1 cu.reg_file.reg_c\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5558__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5221__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4024__A1 _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _0877_ _0904_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__a21o_1
XANTENNA__4575__A2 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3761_ cu.reg_file.reg_a\[6\] _0625_ _0628_ cu.reg_file.reg_mem\[14\] _0836_ vssd1
+ vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__a221o_1
X_5500_ _2319_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3692_ _0754_ _0757_ _0767_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5431_ _2139_ _2205_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5362_ _1261_ net115 _2215_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4313_ _1332_ _1368_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5293_ _1052_ net85 _2182_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__mux2_1
X_4244_ _0992_ _1309_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__and3b_2
X_4175_ _1241_ _1244_ _0588_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__mux2_1
X_3126_ _2770_ _2771_ _2863_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__or3_1
XANTENNA__4356__B _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3057_ ih.t.count\[20\] _2759_ _2793_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5468__A _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _0758_ _1031_ _1033_ _0918_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5629_ _2169_ _2436_ _2443_ _2136_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5407__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5279__A0 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5142__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4557__A2 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3214__C1 _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4309__A2 _1372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output60_A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5980_ clknet_leaf_30_clk _0018_ net187 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4904__B cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4931_ _1921_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__nand2_1
XANTENNA__4192__A _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5288__A _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4862_ _1859_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3813_ cu.reg_file.reg_d\[1\] _0488_ _0741_ cu.reg_file.reg_h\[1\] _0888_ vssd1 vssd1
+ vccd1 vccd1 _0889_ sky130_fd_sc_hd__a221o_1
XANTENNA__6074__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3744_ _0605_ _0553_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3675_ cu.reg_file.reg_mem\[8\] _0640_ _0749_ _0750_ vssd1 vssd1 vccd1 vccd1 _0751_
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5414_ _2253_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 ss3[0] sky130_fd_sc_hd__clkbuf_4
XANTENNA__3536__A _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 ss7[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ss5[6] sky130_fd_sc_hd__clkbuf_4
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ss4[3] sky130_fd_sc_hd__clkbuf_4
X_5345_ _1261_ net107 _2206_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5751__A cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5276_ _2173_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
X_4227_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__buf_2
XANTENNA__4367__A cu.reg_file.reg_l\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4484__A1 cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4158_ _0771_ _0954_ _0779_ _0935_ _0916_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__o32a_1
X_3109_ ih.t.count\[3\] _2846_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__xor2_1
X_4089_ _1161_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4830__A _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3446__A _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4277__A _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 keypad_input[5] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_2
Xinput24 memory_data_in[6] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
XANTENNA__5047__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3460_ _0504_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__clkbuf_4
X_3391_ _2923_ _0354_ net151 _0382_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__a311o_1
X_5130_ _2073_ cu.reg_file.reg_h\[2\] _2069_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__mux2_1
X_5061_ _2028_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4466__B2 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4466__A1 cu.id.imm_i\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4012_ _0610_ _1083_ _0701_ _0611_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3269__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4915__A cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5415__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5966__A1 _2467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5963_ _2691_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4769__A2 _1644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4914_ cu.pc.pc_o\[9\] _1894_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5894_ _1667_ _2205_ _2152_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__o21a_2
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4845_ _1829_ _1832_ _1830_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4776_ _0980_ _1781_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5465__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3727_ _0684_ _0787_ _0682_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3658_ _0733_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__inv_2
X_3589_ _0294_ _0634_ _0374_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__or3b_1
XANTENNA_clkbuf_leaf_27_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5328_ _2149_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5700__A2_N _1643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5259_ _2162_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5709__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5978__RESET_B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2999__B net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout190 net196 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4454__B _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5948__A1 _2467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ _2700_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__clkbuf_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4630_ ih.t.count\[0\] _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4561_ _1305_ _1610_ _1613_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6300_ clknet_leaf_38_clk _0282_ net162 vssd1 vssd1 vccd1 vccd1 cu.id.cb_opcode_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4492_ _1332_ _1530_ _1532_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3512_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__buf_2
X_6231_ clknet_leaf_17_clk net214 net179 vssd1 vssd1 vccd1 vccd1 ih.t.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_3443_ _0384_ _0392_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__or2_1
XANTENNA__5884__A0 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ clknet_leaf_10_clk _0196_ net166 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _0312_ net242 _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__or3_1
XANTENNA__4151__A3 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5113_ cu.reg_file.reg_e\[5\] _1191_ _2056_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__mux2_1
X_6093_ clknet_leaf_13_clk _0127_ net173 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__B1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ cu.reg_file.reg_b\[5\] _2016_ _2006_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout177_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__A1 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5946_ _0373_ _2448_ _2666_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__mux2_1
X_5877_ _1667_ _2180_ _2635_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5476__A _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4828_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3708__B _0587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6007__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4759_ _1760_ _1766_ _1767_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5415__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3090_ ih.t.timer_max\[7\] _2750_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__xor2_1
Xhold2 _0217_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5060__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3992_ _0816_ _0807_ _0776_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5800_ cu.reg_file.reg_sp\[8\] _2535_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__nand2_1
X_5731_ _2518_ mc.cl.next_data\[4\] _2111_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5662_ ih.t.timer_max\[31\] _2145_ _2192_ ih.t.timer_max\[15\] vssd1 vssd1 vccd1
+ vccd1 _2475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4613_ mc.cl.cmp_o _1364_ _1613_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__or3b_1
X_5593_ _2406_ _2407_ _2409_ _1641_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__o22a_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4544_ _1305_ _1594_ _1597_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap143 _0509_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
XFILLER_0_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6214_ clknet_leaf_13_clk ih.t.next_count\[2\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_4475_ _1512_ _1531_ _1520_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__nand3_1
XANTENNA__5857__A0 cu.reg_file.reg_sp\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3426_ net147 _0473_ _0479_ _0486_ _0458_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__o2111a_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ clknet_leaf_10_clk _0179_ net166 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_2
XANTENNA__3332__A1 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3357_ _0412_ _0405_ _0424_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__and3_2
X_6076_ clknet_leaf_23_clk _0110_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _2902_ _2884_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__xnor2_4
X_5027_ _1792_ _2004_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__nor2_1
XANTENNA__4832__A1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5929_ _2673_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4060__A2 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5560__A2 _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3571__A1 cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3571__B2 cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5145__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3323__A1 _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3087__B1 ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5993__RESET_B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output90_A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3562__A1 cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3364__A _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3562__B2 cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4260_ cu.reg_file.reg_c\[0\] _1313_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4191_ _1110_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__buf_4
X_3211_ _2946_ _2947_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__nor2_8
XFILLER_0_5_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3142_ _2875_ _2876_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3073_ _2755_ _2809_ ih.t.count\[14\] vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3975_ _0517_ _1038_ _1039_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__a211o_4
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5714_ ih.input_handler_enable _0618_ _2516_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__mux2_1
X_5645_ ih.t.timer_max\[22\] _2150_ _2319_ ih.t.timer_max\[6\] _1660_ vssd1 vssd1
+ vccd1 vccd1 _2459_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5576_ net127 _2236_ _2247_ net135 vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__a22o_1
XANTENNA__5473__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3553__A1 cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4527_ _1333_ _1561_ _1565_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3274__A _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4458_ _1501_ _1511_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__and2_1
XANTENNA__4502__B1 _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3409_ _0464_ _0480_ _0482_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__a22o_2
X_6128_ clknet_leaf_22_clk _0162_ net190 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_4
X_4389_ cu.reg_file.reg_l\[6\] _1317_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__and2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__B cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5058__A1 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4805__A1 _0359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6059_ clknet_leaf_4_clk _0096_ net157 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3792__B2 cu.reg_file.reg_h\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3792__A1 cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5049__A1 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5839__A cu.reg_file.reg_sp\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5558__B _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ cu.pc.pc_o\[14\] _0740_ _0834_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3783__A1 cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5430_ _2263_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3691_ _0765_ _0766_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5361_ _2222_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4732__A0 cu.alu_f\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5292_ _2183_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4312_ _1376_ _1374_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__nand2_1
XANTENNA__3525__C _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4243_ _2883_ _0320_ _1310_ _0295_ _2914_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__a2111o_2
X_4174_ _1242_ _1243_ _0600_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3125_ _2773_ _2775_ _2776_ _2862_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__or4_1
X_3056_ _2759_ _2793_ ih.t.count\[20\] vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4372__B _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3958_ _1032_ _0807_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5484__A _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3889_ _2897_ _0324_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__nor2_1
X_5628_ ih.gpio_interrupt_mask\[5\] _2326_ _2442_ _2125_ _2327_ vssd1 vssd1 vccd1
+ vccd1 _2443_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5559_ net102 _2205_ _2376_ _1401_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5279__A1 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4282__B _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3214__B1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4962__A0 cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3517__A1 cu.reg_file.reg_l\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6302__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5333__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5690__B2 ih.t.timer_max\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4930_ _1902_ _1910_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__or2b_1
X_4861_ cu.pc.pc_o\[4\] _1858_ _1815_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3812_ cu.reg_file.reg_b\[1\] _0743_ _0624_ cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1
+ vccd1 _0888_ sky130_fd_sc_hd__a22o_1
XANTENNA_27 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3756__A1 cu.reg_file.reg_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4792_ _1793_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3743_ _0753_ _0778_ _0780_ _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3674_ cu.reg_file.reg_b\[0\] _0426_ _0429_ cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1
+ vccd1 _0750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5413_ _1190_ net136 _2248_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__mux2_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 ss3[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__3508__B2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ss5[7] sky130_fd_sc_hd__buf_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 ss7[2] sky130_fd_sc_hd__clkbuf_4
X_5344_ _2213_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__clkbuf_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ss4[4] sky130_fd_sc_hd__clkbuf_4
X_5275_ net78 _1074_ _2170_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4226_ _1293_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__buf_2
XANTENNA__5681__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4484__A2 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4157_ _0935_ _0813_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__xnor2_1
X_3108_ _2747_ _2845_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__nand2_1
X_4088_ _0617_ _1050_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__xor2_1
X_3039_ ih.t.timer_max\[25\] _2762_ ih.t.timer_max\[26\] vssd1 vssd1 vccd1 vccd1 _2777_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__4944__A0 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4830__B cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3747__B2 _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3446__B cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5121__A0 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6195__D net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 keypad_input[6] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 memory_data_in[7] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_1
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3356__B _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5360__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3390_ _0300_ _0353_ _2912_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5060_ cu.reg_file.reg_c\[2\] _1074_ _2025_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__mux2_1
X_4011_ _0606_ _0701_ _1083_ _0603_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__a221o_1
XANTENNA__3674__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5415__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5962_ cu.id.imm_i\[12\] _2429_ _2686_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__mux2_1
X_4913_ _1906_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__clkbuf_1
X_5893_ _2653_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4844_ _1841_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__and2b_1
X_4775_ _0976_ _0989_ _1780_ _0994_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3726_ _0645_ _0799_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4982__B1_N _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3657_ _0732_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__buf_2
X_3588_ _0652_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__xnor2_4
X_5327_ _2203_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5481__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5103__A0 cu.reg_file.reg_e\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ ih.t.timer_max\[28\] _2161_ _2153_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__mux2_1
XANTENNA__5654__A1 _2467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5189_ mc.cl.next_data\[15\] net25 mc.count vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__mux2_1
X_4209_ _2883_ _2937_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5709__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5672__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout191 net193 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_4
XANTENNA_output139_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5847__A cu.reg_file.reg_sp\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ cu.reg_file.reg_h\[7\] _1316_ _1312_ cu.reg_file.reg_b\[7\] _1612_ vssd1 vssd1
+ vccd1 vccd1 _1613_ sky130_fd_sc_hd__a221o_1
XANTENNA__5058__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4384__B2 cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4491_ _1546_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3511_ _0576_ _0581_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__o21ai_2
X_6230_ clknet_leaf_17_clk ih.t.next_count\[18\] net178 vssd1 vssd1 vccd1 vccd1 ih.t.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5333__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3442_ _0401_ _0511_ _0513_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__o211a_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ clknet_leaf_10_clk _0195_ net167 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
X_3373_ _2894_ _2874_ _0309_ _2941_ _0378_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__a32o_2
XANTENNA__4198__A _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5112_ _2061_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
X_6092_ clknet_leaf_24_clk _0126_ net192 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__B2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5043_ _1191_ _1209_ _2002_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__mux2_1
XANTENNA__4926__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4611__A2 _1644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5945_ _2681_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
X_5876_ _2644_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4827_ _1299_ cu.pc.pc_o\[1\] cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758_ _1268_ _1300_ _1756_ _1301_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__and4bb_1
X_4689_ ih.t.count\[18\] _1708_ _1687_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__o21ai_1
X_3709_ _0762_ _0784_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5324__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4127__A1 _0916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4127__B2 _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5875__A1 ih.t.timer_max\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3638__B1 _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4290__B _1354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4366__A1 _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4366__B2 cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3337__D _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5341__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 cu.id.interrupt_requested vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ _0758_ _0760_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__o21bai_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5730_ net21 _2519_ _2525_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5661_ net83 _1633_ _2470_ _2473_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4612_ _2704_ _1647_ _1655_ vssd1 vssd1 vccd1 vccd1 mc.rw.next_state\[0\] sky130_fd_sc_hd__a21o_1
X_5592_ _1649_ _2408_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4543_ cu.reg_file.reg_h\[6\] _1317_ _1313_ cu.reg_file.reg_b\[6\] _1596_ vssd1 vssd1
+ vccd1 vccd1 _1597_ sky130_fd_sc_hd__a221o_1
Xmax_cap144 net238 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6213_ clknet_leaf_14_clk ih.t.next_count\[1\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_4474_ _1512_ _1520_ _1531_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3425_ _0500_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ clknet_leaf_9_clk _0178_ net165 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_4
X_3356_ _0412_ _0405_ _0424_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__and3b_4
X_6075_ clknet_leaf_18_clk _0109_ net180 vssd1 vssd1 vccd1 vccd1 ih.t.enable sky130_fd_sc_hd__dfrtp_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _0360_ _0361_ _0362_ _0297_ _0296_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__5251__S _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5026_ _1790_ _0352_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__nand2_1
XANTENNA__4832__A2 cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5928_ _0359_ _2429_ _2668_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__mux2_1
XANTENNA__3399__A2 _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5859_ _2141_ _2320_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__and2b_2
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4348__A1 cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4348__B2 _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4520__A1 cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__A _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4587__A1 _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output83_A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3210_ cu.id.state\[1\] cu.id.state\[0\] vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4190_ _1259_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__clkbuf_1
X_3141_ cu.id.opcode\[0\] cu.id.opcode\[2\] cu.id.opcode\[1\] vssd1 vssd1 vccd1 vccd1
+ _2878_ sky130_fd_sc_hd__nand3b_4
X_3072_ ih.t.count\[14\] _2755_ _2809_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3974_ _0558_ _1040_ _1043_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5713_ _1328_ _1354_ _2274_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__and3_1
X_5644_ _1400_ _2457_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5575_ _2392_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_4526_ _1396_ _1579_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__nand2_1
XANTENNA__4750__B2 _1269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3553__A2 _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4457_ _1512_ _1513_ _1514_ _1334_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__a31o_1
XANTENNA__4502__B2 cu.id.imm_i\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4502__A1 cu.reg_file.reg_sp\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3408_ _0483_ _0463_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__nor2_1
X_6127_ clknet_leaf_10_clk _0161_ net167 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_4
X_4388_ _0387_ _1295_ _1298_ cu.pc.pc_o\[6\] _1306_ vssd1 vssd1 vccd1 vccd1 _1450_
+ sky130_fd_sc_hd__a221o_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _0414_ _0405_ _0412_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__and3b_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ clknet_leaf_25_clk mc.cc.enable net194 vssd1 vssd1 vccd1 vccd1 mc.cc.enable_edge_detector.prev_data
+ sky130_fd_sc_hd__dfrtp_1
X_5009_ cu.reg_file.reg_a\[3\] _1991_ _1985_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5518__B1 _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3792__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3465__A cu.reg_file.reg_e\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6198__D net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__S _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output121_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5839__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5757__A0 cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5855__A cu.reg_file.reg_sp\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3783__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3690_ _0718_ _0684_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5066__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5360_ _1194_ net114 _2215_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__mux2_1
XANTENNA__4732__A1 alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5291_ _0619_ net84 _2182_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__mux2_1
X_4311_ _1376_ _1348_ _1349_ _1335_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4242_ _2908_ _0361_ _0968_ _0336_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__o31a_1
XFILLER_0_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _0747_ _0892_ _0447_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__mux2_1
X_3124_ _2778_ _2779_ _2861_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__or3_1
X_3055_ ih.t.timer_max\[19\] _2758_ ih.t.timer_max\[20\] vssd1 vssd1 vccd1 vccd1 _2793_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ _0401_ _0528_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__or2_4
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3888_ _0620_ _0819_ _0823_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5627_ mc.cl.next_data\[5\] _2313_ net142 _2441_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__a22o_1
X_5558_ net86 _1330_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__or2_1
XANTENNA__5920__A0 _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4509_ _1546_ _1563_ _1562_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5489_ net124 _2236_ _2247_ net132 _2308_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__a221o_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3462__A1 cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5614__S _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output46_A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4473__B _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4860_ _1850_ _1857_ _1809_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3811_ _0886_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__inv_2
XANTENNA_28 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4791_ _1186_ _1790_ _0352_ _1792_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__or4_2
XFILLER_0_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3742_ _0776_ _0798_ _0815_ _0817_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ cu.reg_file.reg_sp\[8\] _0636_ _0748_ cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1
+ vccd1 _0749_ sky130_fd_sc_hd__a22o_1
X_5412_ _2252_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5343_ _1194_ net106 _2206_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__mux2_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 ss3[2] sky130_fd_sc_hd__clkbuf_4
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ss4[5] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ss6[0] sky130_fd_sc_hd__buf_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 ss7[3] sky130_fd_sc_hd__clkbuf_4
X_5274_ _2172_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5130__A1 cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4225_ _2950_ _1292_ _1269_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__and3_2
XANTENNA__5681__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4156_ _0516_ _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__nor2_4
X_3107_ ih.t.timer_max\[3\] _2746_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__nand2_1
X_4087_ _1144_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__xor2_1
X_3038_ ih.t.count\[27\] _2764_ _2774_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4989_ cu.pc.pc_o\[14\] _1968_ _1233_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4839__A cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5121__A1 _0617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput26 nrst vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput15 keypad_input[7] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5360__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4010_ _0531_ _0694_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4871__A0 _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3674__A1 cu.reg_file.reg_b\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3674__B2 cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _2690_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__clkbuf_1
X_4912_ cu.pc.pc_o\[8\] _1905_ _1815_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__mux2_1
X_5892_ _1260_ ih.t.timer_max\[7\] _2645_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__mux2_1
XANTENNA__5179__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4843_ cu.id.cb_opcode_y\[0\] cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__nand2_1
X_4774_ _2948_ _0986_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3725_ _0733_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3656_ _0730_ _0731_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__or2_1
XANTENNA__5254__S _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3587_ _0653_ _0655_ _0657_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__o22a_4
X_5326_ _1261_ net99 _2195_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__mux2_1
X_5257_ _1160_ _1213_ _1667_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__mux2_1
XANTENNA__5103__A1 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4208_ _2912_ _2937_ _0583_ _1274_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__a31o_2
X_5188_ _1646_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__clkbuf_2
X_4139_ _1203_ _1208_ _0516_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5590__A1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5953__A _2685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout181 net197 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5339__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5581__A1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3510_ _0294_ _0585_ _0576_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__o21ai_1
X_4490_ _1333_ _1545_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5333__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5074__S _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3441_ _0395_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ clknet_leaf_20_clk _0194_ net172 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_4
X_3372_ _2925_ _0313_ _0325_ _2910_ _2879_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__a2111oi_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ cu.reg_file.reg_e\[4\] _1189_ _2056_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__mux2_1
XANTENNA__3895__A1 _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3895__B2 _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ clknet_leaf_21_clk _0125_ net183 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_4
XANTENNA__5636__A2 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _2015_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4926__B _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _0374_ _2429_ _2666_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5875_ _2167_ ih.t.timer_max\[15\] _2636_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4826_ _1299_ cu.pc.pc_o\[1\] cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5021__A0 cu.reg_file.reg_a\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4757_ _1761_ _1764_ _1765_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__a21oi_1
X_4688_ ih.t.count\[18\] _1708_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__and2_1
X_3708_ _0710_ _0587_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5324__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3639_ _0587_ _0710_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3335__B1 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3293__A _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5309_ _2192_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__clkbuf_4
X_6289_ clknet_leaf_42_clk _0271_ net153 vssd1 vssd1 vccd1 vccd1 cu.id.opcode\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__3740__B _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4852__A cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5260__A0 _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5012__A0 cu.reg_file.reg_a\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3187__B _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5563__A1 ih.t.timer_max\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5563__B2 ih.t.timer_max\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4584__D_N _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 _0001_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3629__A1 cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3629__B2 cu.reg_file.reg_a\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5251__A0 _1073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3990_ _0761_ _0772_ _0777_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5660_ net115 _2146_ _2225_ net123 _2472_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__a221o_1
XANTENNA__3378__A _0379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5003__A0 cu.reg_file.reg_a\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4611_ _1650_ _1644_ _1651_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__a31o_1
X_5591_ net11 _2345_ _2369_ net4 vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__a22o_1
XANTENNA__5554__A1 _2372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4542_ cu.pc.pc_o\[14\] _1322_ _1315_ cu.reg_file.reg_d\[6\] _1595_ vssd1 vssd1 vccd1
+ vccd1 _1596_ sky130_fd_sc_hd__a221o_1
X_4473_ _1332_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6212_ clknet_leaf_14_clk ih.t.next_count\[0\] net176 vssd1 vssd1 vccd1 vccd1 ih.t.count\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3424_ cu.id.starting_int_service net150 vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__or2_1
X_6143_ clknet_leaf_12_clk _0177_ net168 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5532__S _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3355_ cu.reg_file.reg_c\[0\] _0427_ _0430_ cu.reg_file.reg_e\[0\] vssd1 vssd1 vccd1
+ vccd1 _0431_ sky130_fd_sc_hd__a22o_1
X_6074_ clknet_leaf_16_clk _0108_ net180 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _2888_ _2890_ _2933_ _2934_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__and4_1
X_5025_ _0618_ _1622_ _2002_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__mux2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4293__A1 cu.reg_file.reg_e\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4293__B2 cu.reg_file.reg_l\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5768__A cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5927_ _2672_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ _2634_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5545__A1 _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4809_ _1301_ _1775_ _1779_ _1268_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__o22ai_1
X_5789_ cu.reg_file.reg_sp\[6\] _2574_ _2539_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__mux2_1
XANTENNA__4348__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4520__A2 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__B _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5678__A _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4582__A _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5352__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3140_ _2875_ _2876_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__nand2b_4
X_3071_ ih.t.timer_max\[13\] _2754_ ih.t.timer_max\[14\] vssd1 vssd1 vccd1 vccd1 _2809_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3483__C1 cu.reg_file.reg_l\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5712_ net190 _2707_ _2514_ _2515_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__a31o_1
X_3973_ _0574_ _0822_ _1046_ _0545_ _1047_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__a221o_1
XANTENNA__3786__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6037__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5643_ ih.t.timer_max\[14\] _2193_ _2314_ ih.t.timer_max\[6\] _2456_ vssd1 vssd1
+ vccd1 vccd1 _2457_ sky130_fd_sc_hd__a221o_1
XANTENNA__5527__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5574_ cu.reg_file.reg_mem\[2\] _2391_ _2351_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__mux2_1
X_4525_ _1396_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4456_ _1512_ _1513_ _1514_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4387_ _1271_ _1448_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3407_ net149 _0454_ _0457_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__a21o_1
X_6126_ clknet_leaf_11_clk _0160_ net167 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_4
X_3338_ _0293_ _0407_ _0408_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__or3b_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ clknet_leaf_22_clk _0095_ net190 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3269_ _0340_ _0341_ _0342_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5008_ _1187_ _1222_ _0368_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5215__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5518__A1 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_25_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4257__A1 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output114_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4743__C _0379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3359__C _0379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4310_ mc.rw.state\[2\] _2699_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__nand2_1
X_5290_ _2180_ _2181_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__nand2_8
XFILLER_0_77_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4241_ _0336_ _0436_ _1308_ _0295_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__a211o_2
X_4172_ _0871_ _0902_ _1060_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__mux2_1
X_3123_ _2781_ _2783_ _2784_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__or4_1
X_3054_ _2760_ _2790_ ih.t.count\[21\] vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4950__A cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3956_ _1030_ _1029_ _0773_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5626_ _1666_ _2439_ _2440_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__o21a_1
XANTENNA__5257__S _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3887_ _0824_ _0915_ _0962_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__and3_1
X_5557_ net94 _2194_ _2374_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__a21o_1
XANTENNA__5920__A1 _2350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4508_ _1546_ _1562_ _1563_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__nand3_1
X_5488_ net84 _2180_ _2224_ net116 vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__a22o_1
X_4439_ _1497_ _1480_ _1481_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__nand3_1
Xwire2 _1280_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4487__A1 cu.reg_file.reg_h\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4487__B2 cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6109_ clknet_leaf_28_clk _0143_ net186 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4239__A1 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4239__B2 _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3462__A2 _0492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__A1 cu.reg_file.reg_c\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3476__A _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4478__A1 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6311__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4790_ _1791_ _0366_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__or2_2
X_3810_ _0882_ _0885_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__xor2_1
XANTENNA_29 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3741_ _0816_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3610__C1 cu.reg_file.reg_l\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3672_ _0417_ _0421_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__nor2_4
XFILLER_0_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5411_ _1188_ net135 _2248_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ss4[6] sky130_fd_sc_hd__clkbuf_4
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ss6[1] sky130_fd_sc_hd__clkbuf_4
X_5342_ _2212_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3913__B1 _0296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ss3[3] sky130_fd_sc_hd__clkbuf_4
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 ss7[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5273_ net77 _1051_ _2170_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__mux2_1
XANTENNA__4469__B2 cu.id.imm_i\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4469__A1 cu.reg_file.reg_sp\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4224_ _2904_ _2924_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__nand2_1
X_4155_ _0955_ _1215_ _1216_ _0952_ _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__o221a_1
X_3106_ _2749_ _2835_ ih.t.count\[4\] vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4086_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__buf_4
X_3037_ _2764_ _2774_ ih.t.count\[27\] vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5776__A cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4988_ cu.pc.pc_o\[15\] _1963_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3296__A cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3939_ _0983_ _0996_ _1003_ _1011_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5609_ _2169_ _2417_ _2424_ _2136_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__o211a_1
XANTENNA__5409__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4590__A _1415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3821__B_N _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput27 programmable_gpio_in[0] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput16 keypad_input[8] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_2
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5360__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3674__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5960_ cu.id.imm_i\[11\] _2410_ _2686_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__mux2_1
XANTENNA__3595__A1_N _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5820__A0 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5891_ _2652_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
X_4911_ _1896_ _1904_ _1809_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4842_ cu.id.cb_opcode_y\[0\] cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4773_ net206 _1779_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _0644_ _0799_ _0790_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3655_ _0566_ _0729_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__nor2_1
XANTENNA__4139__B1 _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3844__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3586_ _0659_ _0660_ _0661_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__or3_2
X_5325_ _2202_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
X_5256_ _2160_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_1
X_4207_ _2912_ _0583_ _1273_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__a31o_1
X_5187_ _2110_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3356__A_N _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4394__B _1455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4138_ _0916_ _0943_ _1206_ _0950_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4069_ _1135_ _1138_ _1141_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5590__A2 _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5878__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3904__D _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout182 net184 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4585__A _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout171 net172 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout193 net196 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5581__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3664__A _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3440_ _0515_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__buf_8
X_3371_ _0416_ _0420_ _0441_ _0446_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__o31a_4
XANTENNA__3344__B2 cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ clknet_leaf_7_clk _0124_ net171 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_4
X_5110_ _2060_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ cu.reg_file.reg_b\[4\] _2014_ _2006_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__mux2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5090__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5943_ _2680_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
X_5874_ _2643_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
X_4825_ _1825_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4756_ _1268_ _1301_ _1300_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3583__A1 cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4687_ _1710_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__4780__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3707_ _0781_ _0712_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3638_ _0712_ _0713_ _0545_ _0599_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3293__B _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3569_ _0644_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__inv_2
X_5308_ _1374_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3886__A2 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6288_ clknet_leaf_42_clk _0270_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.opcode\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_5239_ _2146_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5260__A1 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3574__B2 cu.reg_file.reg_a\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3629__A2 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5 ih.interrupt_source\[1\] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5251__A1 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3659__A _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4610_ _2701_ _2706_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5590_ net71 _1648_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4541_ cu.reg_file.reg_sp\[14\] _0992_ _1344_ cu.id.imm_i\[14\] _1324_ vssd1 vssd1
+ vccd1 vccd1 _1595_ sky130_fd_sc_hd__a221o_1
X_4472_ _1305_ _1526_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6211_ clknet_leaf_7_clk ih.ih.int_f.data_in net181 vssd1 vssd1 vccd1 vccd1 ih.ih.int_f.prev_data
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap146 net240 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
X_3423_ net147 _0473_ net146 _0486_ _0458_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__o2111a_4
X_6142_ clknet_leaf_13_clk _0176_ net173 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3354_ _0425_ _0414_ _0429_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6073_ clknet_leaf_19_clk _0107_ net180 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3841__B _0916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3285_ _0342_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__clkbuf_4
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _2001_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__buf_4
XANTENNA__5490__B2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5490__A1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4953__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5926_ _2893_ _2410_ _2668_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5784__A cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5857_ cu.reg_file.reg_sp\[15\] _2633_ _2538_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__mux2_1
X_4808_ _1788_ _1800_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__mux2_1
X_5788_ _1126_ _2573_ _2545_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__mux2_1
X_4739_ _1012_ _1747_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4863__A cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3492__B1 _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4992__A0 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3795__A1 cu.id.imm_i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3547__A1 cu.reg_file.reg_c\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output69_A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3070_ ih.t.count\[15\] _2756_ _2806_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__and3_1
XANTENNA__5971__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5711_ net190 mc.cl.cmp_o vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__and2b_1
XANTENNA__4983__A0 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3972_ _0531_ _0545_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__nor2_1
XANTENNA__3786__A1 cu.reg_file.reg_sp\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3786__B2 cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5642_ ih.t.timer_max\[30\] _2146_ _2149_ ih.t.timer_max\[22\] vssd1 vssd1 vccd1
+ vccd1 _2456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5573_ _2387_ _2388_ _2390_ _1641_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__o22a_2
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4524_ _1304_ _1575_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__o21a_2
X_4455_ _1396_ _1496_ _1498_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__a21bo_1
X_4386_ cu.reg_file.reg_c\[6\] _1281_ _1447_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__a21oi_1
X_3406_ _0468_ _0473_ net146 vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__nor3_4
X_6125_ clknet_leaf_13_clk _0159_ net173 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_3337_ _0405_ _0407_ _0409_ _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__and4bb_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ clknet_leaf_22_clk _0094_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3268_ _0343_ cu.id.cb_opcode_z\[1\] cu.id.cb_opcode_z\[2\] vssd1 vssd1 vccd1 vccd1
+ _0344_ sky130_fd_sc_hd__nand3_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3199_ _2884_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__clkbuf_4
X_5007_ _1990_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3299__A _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3777__A1 cu.reg_file.reg_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5909_ ih.t.timer_max\[23\] _1260_ _2654_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4032__A1_N alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5151__A0 cu.reg_file.reg_l\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5454__A1 _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4257__A2 _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4593__A _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3002__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output107_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6170__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5390__A0 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4240_ _0359_ _0320_ _0336_ _2914_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__a211oi_1
XANTENNA__5693__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4171_ _1239_ _1240_ _0600_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__mux2_1
X_3122_ _2786_ _2787_ _2859_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3053_ ih.t.count\[21\] _2760_ _2790_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__and3_1
XANTENNA__3824__A1_N _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4956__B1 _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3955_ _0511_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__inv_2
XANTENNA__3759__B2 cu.reg_file.reg_sp\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3759__A1 cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5625_ ih.t.timer_max\[21\] _2150_ _2319_ ih.t.timer_max\[5\] _1661_ vssd1 vssd1
+ vccd1 vccd1 _2440_ sky130_fd_sc_hd__a221o_1
X_3886_ _0918_ _0779_ _0932_ _0947_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__a311o_1
XFILLER_0_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5381__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5556_ net126 _2236_ _2247_ net134 vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5273__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4507_ _1333_ _1545_ _1549_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__a21o_1
X_5487_ _2307_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4438_ _1480_ _1481_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__a21o_1
XANTENNA__5684__B2 _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ cu.pc.pc_o\[5\] _1322_ _1315_ cu.reg_file.reg_e\[5\] _1431_ vssd1 vssd1 vccd1
+ vccd1 _1432_ sky130_fd_sc_hd__a221o_1
X_6108_ clknet_leaf_28_clk _0142_ net195 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ clknet_leaf_33_clk _0077_ net163 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4947__A0 cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3989__B2 _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5358__S _2215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_19 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _0401_ _0528_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3671_ cu.id.imm_i\[8\] _0739_ _0746_ _0653_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__a22oi_4
X_5410_ _2251_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ss4[7] sky130_fd_sc_hd__buf_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ss3[4] sky130_fd_sc_hd__clkbuf_4
X_5341_ _1192_ net105 _2206_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__mux2_1
XANTENNA__5093__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 ss7[5] sky130_fd_sc_hd__clkbuf_4
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ss6[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5666__A1 _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5272_ _2171_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4223_ _1271_ _1290_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__nor2_1
X_4154_ _0817_ _0939_ _1223_ _0938_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__o2bb2a_1
X_3105_ ih.t.count\[4\] _2749_ _2835_ _2842_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__a31o_1
X_4085_ _1150_ _1151_ _1152_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__or4b_1
X_3036_ ih.t.timer_max\[27\] _2763_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4929__B1 _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4987_ _1974_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__clkbuf_1
X_3938_ alu.Cin _1013_ _1012_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5792__A cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3869_ _0942_ _0943_ _0944_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__and3_1
XANTENNA__5354__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5608_ ih.gpio_interrupt_mask\[4\] _2326_ _2423_ _2125_ _2327_ vssd1 vssd1 vccd1
+ vccd1 _2424_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5539_ net77 _1633_ _2354_ _2357_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5657__A1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3716__A1_N _0733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 keypad_input[9] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_4
Xinput28 programmable_gpio_in[1] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
XANTENNA__5345__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4320__A1 cu.reg_file.reg_e\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4320__B2 cu.reg_file.reg_l\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5890_ _1193_ ih.t.timer_max\[6\] _2645_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__mux2_1
X_4910_ _1799_ _1897_ _1902_ _1903_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__a22o_1
X_4841_ _1838_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4772_ _1301_ _1777_ _1778_ _1303_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3723_ _0664_ _0684_ _0787_ _0794_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3654_ _0566_ _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3585_ cu.reg_file.reg_c\[5\] _0485_ _0621_ cu.reg_file.reg_l\[5\] vssd1 vssd1 vccd1
+ vccd1 _0661_ sky130_fd_sc_hd__a22o_1
XANTENNA__5639__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5324_ _1194_ net98 _2195_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5255_ ih.t.timer_max\[27\] _2159_ _2153_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__mux2_1
XANTENNA__5639__B2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4311__B2 _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4206_ _0336_ _1266_ _0293_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__a21o_1
X_5186_ _1647_ _2109_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _0950_ _1204_ _0773_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4068_ _0570_ _0664_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__nor2_1
X_3019_ ih.t.timer_max\[16\] ih.t.timer_max\[17\] _2756_ vssd1 vssd1 vccd1 vccd1 _2757_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5878__A1 ih.t.timer_max\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4866__A _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout172 net181 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_4
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4369__A1 cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4369__B2 cu.reg_file.reg_e\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5318__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5869__A1 ih.t.timer_max\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output99_A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ _2949_ _0445_ _0440_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4541__A1 cu.reg_file.reg_sp\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4541__B2 cu.id.imm_i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5371__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5040_ _1189_ _1213_ _2002_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__mux2_1
XANTENNA__4495__B _1545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5942_ cu.id.cb_opcode_y\[0\] _2410_ _2666_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5873_ _2165_ ih.t.timer_max\[14\] _2636_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4824_ cu.pc.pc_o\[1\] _1824_ _1815_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4016__A _1073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4755_ _1756_ _1763_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _0545_ _0600_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4686_ _1708_ _1709_ _1672_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3637_ _0575_ net143 vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3568_ _0632_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__xnor2_2
X_5307_ _1329_ _1354_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5281__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ clknet_leaf_42_clk _0269_ net152 vssd1 vssd1 vccd1 vccd1 cu.id.opcode\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3499_ _0416_ _0420_ _0441_ _0446_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__o31ai_2
X_5238_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__clkbuf_4
X_5169_ _2098_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4048__B1 _0916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5796__A0 _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4523__A1 cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4523__B2 cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 cu.id.can_be_interrupted vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output137_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4540_ cu.pc.pc_o\[14\] _1485_ _1593_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4471_ cu.reg_file.reg_h\[2\] _1317_ _1312_ cu.reg_file.reg_b\[2\] _1528_ vssd1 vssd1
+ vccd1 vccd1 _1529_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6201__D net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6210_ clknet_leaf_9_clk net8 net166 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap147 _0468_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_4
X_3422_ net147 _0473_ net239 _0486_ _0483_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6141_ clknet_leaf_24_clk _0175_ net192 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _0428_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__clkbuf_4
X_6072_ clknet_leaf_16_clk _0106_ net174 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _0340_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__inv_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _1790_ _0352_ _1791_ _0366_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__and4b_1
XANTENNA__4953__B cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5925_ _2671_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5856_ _1263_ _2632_ _2115_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__mux2_1
X_4807_ _1808_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__buf_4
X_2999_ net70 net29 ih.gpio_interrupt_mask\[2\] vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__and3b_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5787_ _2571_ _2572_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5950__A0 _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4738_ _0456_ _1746_ _2950_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__o21ai_2
X_4669_ _1698_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4863__B cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5678__C _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4680__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3971_ _0600_ _1044_ _1042_ _0610_ _1045_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_85_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5710_ _2708_ _1653_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ net82 _1633_ _2451_ _2454_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__o22a_1
XANTENNA__5096__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5572_ _1649_ _2389_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__and2_1
X_4523_ cu.reg_file.reg_h\[5\] _1316_ _1312_ cu.reg_file.reg_b\[5\] _1577_ vssd1 vssd1
+ vccd1 vccd1 _1578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4454_ _1332_ _1511_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3405_ net149 _0476_ _0478_ _0382_ _0465_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__a2111oi_1
X_4385_ cu.reg_file.reg_e\[6\] _1283_ _1285_ cu.reg_file.reg_l\[6\] _1446_ vssd1 vssd1
+ vccd1 vccd1 _1447_ sky130_fd_sc_hd__a221o_1
X_6124_ clknet_leaf_23_clk _0158_ net192 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
X_3336_ _0410_ _0411_ cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__a21o_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ clknet_leaf_24_clk _0093_ net191 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4964__A cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3267_ cu.id.cb_opcode_z\[0\] vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__buf_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ cu.reg_file.reg_a\[2\] _1989_ _1985_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__mux2_1
XANTENNA__4671__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3198_ _2888_ _2890_ _2933_ _2934_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__nand4_4
XANTENNA__3299__B _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5908_ _2661_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5839_ cu.reg_file.reg_sp\[13\] _2536_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5151__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4662__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4114__A _1089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5390__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output81_A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5142__A1 cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5693__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4170_ _0850_ _0861_ _1060_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__mux2_1
X_3121_ _2789_ _2791_ _2792_ _2858_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__or4_1
XANTENNA__4653__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3052_ ih.t.timer_max\[21\] _2759_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4956__A1 cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3954_ _0712_ _0713_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__xor2_1
XANTENNA__3759__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4420__A3 _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3885_ _0914_ _0960_ _0773_ _0777_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5624_ _1400_ _2438_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5381__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5554__S _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5555_ _2373_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4506_ _1333_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__xnor2_1
X_5486_ net67 _0618_ _2306_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__mux2_1
X_4437_ _1396_ _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5133__A1 cu.reg_file.reg_h\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire4 _0481_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_1
X_6107_ clknet_leaf_27_clk _0141_ net195 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ cu.reg_file.reg_sp\[5\] _0993_ _1344_ _0373_ _1364_ vssd1 vssd1 vccd1 vccd1
+ _1431_ sky130_fd_sc_hd__a221o_1
X_3319_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__buf_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ cu.reg_file.reg_sp\[2\] _0993_ _1344_ _0341_ _1364_ vssd1 vssd1 vccd1 vccd1
+ _1365_ sky130_fd_sc_hd__a221o_1
X_6038_ clknet_leaf_33_clk _0076_ net164 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5124__A1 cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3570__C_N _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3670_ cu.reg_file.reg_a\[0\] _0625_ _0628_ cu.reg_file.reg_mem\[8\] _0745_ vssd1
+ vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ss5[0] sky130_fd_sc_hd__buf_2
X_5340_ _2211_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__clkbuf_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ss3[5] sky130_fd_sc_hd__buf_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 ss7[6] sky130_fd_sc_hd__clkbuf_4
X_5271_ net76 _2085_ _2170_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ss6[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5115__A1 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4222_ cu.reg_file.reg_c\[0\] _1281_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4874__A0 cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4153_ _0816_ _0936_ _0776_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__a21oi_1
X_3104_ _2837_ _2838_ _2840_ _2841_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__or4_1
X_4084_ _1045_ _0681_ _1155_ _1157_ _0531_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__a32o_1
XANTENNA__3429__A1 cu.pc.pc_o\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3035_ ih.t.count\[28\] _2772_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3429__B2 cu.reg_file.reg_b\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4986_ cu.pc.pc_o\[14\] _1973_ _1814_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__mux2_1
XANTENNA__4929__A1 cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3937_ _0372_ _2921_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3601__A1 cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3601__B2 cu.reg_file.reg_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3868_ _0844_ _0929_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__xnor2_1
X_5607_ mc.cl.next_data\[4\] _2313_ net142 _2422_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__a22o_1
XANTENNA__5354__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3799_ _0871_ _0874_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__and2b_1
X_5538_ net109 _2147_ _2225_ net117 _2356_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__a221o_1
XANTENNA__4379__B1_N _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5469_ _2293_ _2284_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__nor2_1
XANTENNA__3668__A1 cu.reg_file.reg_b\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3668__B2 cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4590__C _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3918__D _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 memory_data_in[0] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5345__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 programmable_gpio_in[2] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3008__A ih.t.timer_max\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5922__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output44_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5281__A0 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5369__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4840_ cu.pc.pc_o\[3\] _1826_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__nor2_1
XANTENNA__6204__D net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _1268_ _1012_ _1646_ _1301_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3722_ _0796_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3653_ _0576_ _0723_ _0725_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5323_ _2201_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3584_ cu.reg_file.reg_e\[5\] _0489_ _0495_ cu.reg_file.reg_h\[5\] _0536_ vssd1 vssd1
+ vccd1 vccd1 _0660_ sky130_fd_sc_hd__a221o_1
X_5254_ _1089_ _1222_ _1667_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__mux2_1
XANTENNA__4847__A0 _1089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5185_ mc.cl.next_data\[14\] net24 mc.count vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__mux2_1
XANTENNA__4311__A2 _1348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4205_ _0359_ _2937_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__or2_1
X_4136_ _0918_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__and2_1
X_4067_ _0558_ _0632_ _0663_ _1139_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__a221o_1
X_3018_ ih.t.timer_max\[15\] _2755_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__or2_2
XANTENNA__5279__S _2170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4969_ _1956_ _1957_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5308__A _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4866__B cu.pc.pc_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3510__B1 _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout162 net197 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5263__A0 _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3813__A1 cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__B2 cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5015__A0 cu.reg_file.reg_a\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5566__A1 _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5318__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3329__B1 cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5254__A0 _1089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4792__A _1793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _2679_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5099__S _2039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3804__A1 cu.pc.pc_o\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5872_ _2642_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5006__A0 cu.reg_file.reg_a\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5557__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4823_ _1817_ _1823_ _1809_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__mux2_1
XANTENNA__4016__B _1089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4754_ _2904_ _2924_ _1318_ _1762_ _0350_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__a41o_1
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3705_ _0447_ net143 vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4685_ ih.t.count\[15\] ih.t.count\[16\] _1702_ ih.t.count\[17\] vssd1 vssd1 vccd1
+ vccd1 _1709_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3636_ _0545_ _0598_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3567_ _0576_ _0635_ _0638_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__o2bb2a_2
X_5306_ _2190_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__clkbuf_1
X_6286_ clknet_leaf_37_clk _0268_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.can_be_interrupted
+ sky130_fd_sc_hd__dfrtp_1
X_5237_ _1369_ _1625_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__nor2_1
X_3498_ net143 vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__inv_2
XANTENNA__4178__S _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4296__A1 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4296__B2 cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5168_ _1647_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__and2_1
X_5099_ cu.reg_file.reg_d\[7\] _2053_ _2039_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__mux2_1
X_4119_ net212 _1186_ _0370_ _1190_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a22o_1
XANTENNA__4048__A1 _1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4220__A1 cu.reg_file.reg_a\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4220__B2 cu.reg_file.reg_sp\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4877__A cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 cu.id.is_interrupted vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3005__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5236__A0 _0617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4117__A _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4470_ _1521_ _1321_ _1314_ cu.reg_file.reg_d\[2\] _1527_ vssd1 vssd1 vccd1 vccd1
+ _1528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4787__A _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3421_ cu.reg_file.reg_d\[0\] _0492_ _0494_ cu.reg_file.reg_mem\[0\] _0496_ vssd1
+ vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__a221o_1
X_6140_ clknet_leaf_24_clk _0174_ net192 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3352_ _0412_ _0405_ _0409_ _0407_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__and4b_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6071_ clknet_leaf_12_clk _0105_ net174 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3283_ _2902_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4278__B2 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4278__A1 cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _2000_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4450__A1 cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5924_ _2899_ _2391_ _2668_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__mux2_1
XANTENNA__4450__B2 cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5855_ cu.reg_file.reg_sp\[15\] _2631_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4806_ _2935_ _1256_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__o21ai_4
X_2998_ _2734_ net28 ih.gpio_interrupt_mask\[1\] _2735_ vssd1 vssd1 vccd1 vccd1 _2736_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5786_ _2562_ _2565_ _2563_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5950__A1 _2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4737_ _0302_ _1266_ _1745_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4668_ _1696_ _1697_ _1672_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__and3b_1
XANTENNA__3961__B1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3619_ _0294_ _0692_ _0634_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__or3_1
X_4599_ _1634_ _1636_ _1641_ _1642_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__nand4_4
XFILLER_0_86_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6269_ clknet_leaf_15_clk _0251_ net175 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4269__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5466__A0 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3952__B1 _1027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5930__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3016__A ih.t.timer_max\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4432__A1 cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3970_ _0603_ _0606_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5377__S _2226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5640_ net114 _2147_ _2225_ net122 _2453_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5571_ net10 _2345_ _2369_ net3 vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5932__A1 _2467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4522_ cu.pc.pc_o\[13\] _1321_ _1314_ cu.reg_file.reg_d\[5\] _1576_ vssd1 vssd1 vccd1
+ vccd1 _1577_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4453_ _1332_ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__or2_1
XANTENNA__5696__B1 cu.reg_file.reg_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4499__A1 cu.id.imm_i\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4499__B2 cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3404_ net147 _0473_ _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor3_2
XFILLER_0_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4384_ cu.reg_file.reg_a\[6\] _1276_ _1287_ cu.reg_file.reg_sp\[6\] vssd1 vssd1 vccd1
+ vccd1 _1446_ sky130_fd_sc_hd__a22o_1
X_6123_ clknet_leaf_16_clk _0157_ net174 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XANTENNA__5448__A0 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3335_ _2900_ _2878_ _2877_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a21o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ clknet_leaf_22_clk _0092_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3266_ _2885_ _2927_ _2917_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__and3_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _1074_ _1226_ _0368_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__mux2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3197_ cu.id.alu_opcode\[0\] cu.id.opcode\[0\] vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5907_ ih.t.timer_max\[22\] _1193_ _2654_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5620__B1 _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3631__C1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5838_ _2617_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
X_5769_ _2555_ _2556_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4890__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5914__A1 _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output74_A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3120_ _2794_ _2795_ _2857_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3051_ ih.t.count\[22\] _2788_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5850__A0 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6207__D net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4405__A1 cu.reg_file.reg_c\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4956__A2 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3953_ _0370_ _0619_ _1026_ _1028_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3884_ _0948_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5623_ ih.t.timer_max\[13\] _2193_ _2314_ ih.t.timer_max\[5\] _2437_ vssd1 vssd1
+ vccd1 vccd1 _2438_ sky130_fd_sc_hd__a221o_1
XANTENNA__5905__A1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5554_ cu.reg_file.reg_mem\[1\] _2372_ _2351_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__mux2_1
X_5485_ _2305_ _2284_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__nor2_1
X_4505_ _1305_ _1557_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4436_ _1305_ _1492_ _1495_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__o21a_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4367_ cu.reg_file.reg_l\[5\] _1317_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__and2_1
XANTENNA__4975__A cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6106_ clknet_leaf_28_clk _0140_ net186 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3318_ _0377_ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _1324_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__buf_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[3\] vssd1 vssd1 vccd1 vccd1 _0325_
+ sky130_fd_sc_hd__or2_1
X_6037_ clknet_leaf_33_clk _0075_ net163 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4215__A _1282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4580__B1 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3013__B ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output112_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5060__A1 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ss3[6] sky130_fd_sc_hd__buf_2
XANTENNA__4571__B1 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _2169_ _2140_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__nor2_4
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ss5[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 ss7[7] sky130_fd_sc_hd__buf_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ss6[4] sky130_fd_sc_hd__clkbuf_4
X_4221_ cu.reg_file.reg_e\[0\] _1283_ _1285_ cu.reg_file.reg_l\[0\] _1288_ vssd1 vssd1
+ vccd1 vccd1 _1289_ sky130_fd_sc_hd__a221o_1
XANTENNA__5390__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ _1217_ _1221_ _0824_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__o21a_4
X_3103_ _2746_ _2839_ ih.t.count\[2\] vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__a21oi_1
X_4083_ _0606_ _0671_ _0681_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__a211oi_1
XANTENNA__3429__A2 _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3034_ ih.t.timer_max\[28\] _2764_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4985_ _1965_ _1972_ _1808_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__mux2_1
XANTENNA__4929__A2 cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3936_ _0296_ _2918_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3867_ _0856_ _0927_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__xnor2_2
X_5606_ _1666_ _2420_ _2421_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__o21a_1
X_3798_ cu.reg_file.reg_mem\[11\] _0640_ _0872_ _0873_ vssd1 vssd1 vccd1 vccd1 _0874_
+ sky130_fd_sc_hd__a211oi_2
X_5537_ net101 _2205_ _2355_ _1401_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3365__A1 cu.reg_file.reg_l\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5468_ _2205_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__inv_2
X_5399_ _2244_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
X_4419_ _1382_ _1475_ _1476_ _1479_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__a31o_1
XANTENNA__3668__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput19 memory_data_in[1] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4553__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3008__B ih.t.timer_max\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5805__A0 cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output37_A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5281__A1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4770_ _1300_ _1761_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3721_ _0752_ _0789_ _0792_ _0795_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nand4_1
XFILLER_0_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3652_ cu.reg_file.reg_l\[7\] _0422_ _0726_ _0727_ _0440_ vssd1 vssd1 vccd1 vccd1
+ _0728_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_2_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3583_ cu.reg_file.reg_sp\[5\] _0539_ _0494_ cu.reg_file.reg_mem\[5\] _0658_ vssd1
+ vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__a221o_1
X_5322_ _1192_ net97 _2195_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5253_ _2158_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__clkbuf_1
X_5184_ _2108_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
X_4204_ _0469_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__inv_2
X_4135_ _1204_ _0779_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__or2_1
XANTENNA__4075__A2 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4066_ _0531_ _0663_ _0681_ _0822_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__a2bb2o_1
X_3017_ ih.t.timer_max\[13\] ih.t.timer_max\[14\] _2754_ vssd1 vssd1 vccd1 vccd1 _2755_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4968_ _1943_ _1948_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__and2b_1
XANTENNA__5295__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4899_ _1893_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3919_ _0986_ _0989_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nand3b_1
XANTENNA__6282__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6211__RESET_B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4299__C1 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout174 net177 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_4
Xfanout163 net164 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_4
Xfanout196 net197 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
Xfanout185 net196 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5263__A1 _1624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3501__B2 cu.reg_file.reg_e\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5254__A1 _1222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5940_ _0341_ _2391_ _2666_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__mux2_1
XANTENNA__3804__A2 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5871_ _2163_ ih.t.timer_max\[13\] _2636_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5557__A2 _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4822_ _1821_ _1822_ _1799_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__mux2_1
X_4753_ net150 _2952_ _0307_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3704_ _0768_ _0770_ _0753_ _0779_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__nor4_1
X_4684_ ih.t.count\[16\] ih.t.count\[17\] _1705_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4517__B1 _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3635_ _0587_ _0710_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3566_ cu.reg_file.reg_l\[6\] _0422_ _0639_ _0641_ _0576_ vssd1 vssd1 vccd1 vccd1
+ _0642_ sky130_fd_sc_hd__a2111o_1
X_5305_ _1261_ net91 _2182_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__mux2_1
X_3497_ _0514_ _0529_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__or2_1
X_6285_ clknet_leaf_38_clk _0267_ net161 vssd1 vssd1 vccd1 vccd1 cu.ir.idx\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__4686__C _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5236_ _0617_ _1622_ _1667_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5167_ mc.cl.next_data\[8\] net18 mc.count vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__mux2_1
XANTENNA__5245__A1 _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4118_ _1189_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__buf_4
X_5098_ _1110_ _1263_ _2035_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__mux2_1
X_4049_ _0802_ _1122_ _0812_ _1032_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold8 ih.interrupt_source\[2\] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5236__A1 _1622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__A0 cu.pc.pc_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3798__A1 cu.reg_file.reg_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5928__S _2668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5539__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4787__B _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap149 net241 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3420_ cu.reg_file.reg_sp\[0\] _0480_ _0493_ _0495_ cu.reg_file.reg_h\[0\] vssd1
+ vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3351_ _0423_ _0424_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a21o_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6070_ clknet_leaf_12_clk _0104_ net168 vssd1 vssd1 vccd1 vccd1 ih.gpio_interrupt_mask\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _2915_ _0353_ _0357_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__o21ba_1
XANTENNA__4278__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ cu.reg_file.reg_a\[7\] _1999_ _1985_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__mux2_1
XANTENNA__4986__A0 cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3212__A cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5923_ _2670_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5854_ _1589_ _2630_ _2626_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4805_ _0359_ _0304_ _1801_ _1804_ _1806_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__o2111a_2
XANTENNA__4738__B1 _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2997_ net68 net27 ih.gpio_interrupt_mask\[0\] vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5785_ _2569_ _2570_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__nand2_1
X_4736_ _2897_ _2941_ _1742_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4667_ ih.t.count\[10\] _1693_ ih.t.count\[11\] vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__a21o_1
XANTENNA__4978__A _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3618_ _0687_ _0689_ _0691_ _0693_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__o31a_4
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4598_ _1415_ _1629_ _1637_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__or3_2
XANTENNA__4189__S _1027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3549_ _0498_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__clkbuf_4
X_6268_ clknet_leaf_13_clk _0250_ net174 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5466__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5219_ _1190_ ih.gpio_interrupt_mask\[4\] _2127_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__mux2_1
X_6199_ clknet_leaf_11_clk net12 net168 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3952__A1 alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4901__B1 cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3468__B1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__6314__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4432__A2 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ net70 _1648_ _2137_ _2274_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4521_ cu.reg_file.reg_sp\[13\] _0992_ _1343_ cu.id.imm_i\[13\] _1323_ vssd1 vssd1
+ vccd1 vccd1 _1576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4452_ _1505_ _1506_ _1510_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5696__B2 _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3403_ net241 _0476_ _0478_ _0382_ _0465_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__a2111o_2
X_4383_ _1423_ _1437_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6122_ clknet_leaf_11_clk _0156_ net167 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_4
X_3334_ _2925_ _2932_ _0364_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__or3_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ clknet_leaf_22_clk _0091_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3265_ cu.id.cb_opcode_z\[2\] vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__buf_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _1988_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__clkbuf_1
X_3196_ _2899_ _2900_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4959__B1 _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ _2660_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5620__B2 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5620__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5837_ cu.reg_file.reg_sp\[12\] _2616_ _2538_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5768_ cu.reg_file.reg_sp\[4\] _2534_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__and2_1
X_4719_ net221 _1729_ _1731_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[28\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5699_ mc.cl.next_data\[13\] _2359_ _2490_ _2505_ vssd1 vssd1 vccd1 vccd1 _2506_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4890__B cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5611__B2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5611__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5375__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5507__A _1415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3653__A1_N _0576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output67_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3050_ ih.t.timer_max\[22\] _2760_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5388__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3952_ alu.Cin _1023_ _1027_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3883_ _0949_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5622_ ih.t.timer_max\[29\] _2146_ _2204_ ih.t.timer_max\[21\] vssd1 vssd1 vccd1
+ vccd1 _2437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5553_ _2367_ _2368_ _2371_ _1641_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__o22a_2
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4504_ cu.reg_file.reg_h\[4\] _1316_ _1312_ cu.reg_file.reg_b\[4\] _1559_ vssd1 vssd1
+ vccd1 vccd1 _1560_ sky130_fd_sc_hd__a221o_1
X_5484_ _2247_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__inv_2
X_4435_ cu.reg_file.reg_h\[0\] _1316_ _1312_ cu.reg_file.reg_b\[0\] _1494_ vssd1 vssd1
+ vccd1 vccd1 _1495_ sky130_fd_sc_hd__a221o_1
X_4366_ _0373_ _1295_ _1298_ cu.pc.pc_o\[5\] _1306_ vssd1 vssd1 vccd1 vccd1 _1429_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire6 _0448_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_1
X_6105_ clknet_leaf_9_clk _0139_ net165 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4975__B cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3317_ _0384_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__or2b_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ cu.reg_file.reg_e\[2\] _1315_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__and2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[3\] vssd1 vssd1 vccd1 vccd1 _0324_
+ sky130_fd_sc_hd__nand2_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ clknet_leaf_33_clk _0074_ net163 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4991__A cu.pc.pc_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3179_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[3\] cu.id.opcode\[0\] cu.id.alu_opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__or4bb_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5109__A0 cu.reg_file.reg_e\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4580__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4580__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4231__A cu.pc.pc_o\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4399__A1 _1455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output105_A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5596__B1 _2247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3310__A _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3071__A1 ih.t.timer_max\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5348__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5936__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5899__A1 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5237__A _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4571__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4571__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ss3[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ss6[5] sky130_fd_sc_hd__clkbuf_4
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ss5[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__4323__A1 cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4323__B2 cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4220_ cu.reg_file.reg_a\[0\] _1276_ _1287_ cu.reg_file.reg_sp\[0\] vssd1 vssd1 vccd1
+ vccd1 _1288_ sky130_fd_sc_hd__a22o_1
X_4151_ _0951_ _1214_ _0773_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__a31o_1
X_3102_ ih.t.count\[2\] _2746_ _2839_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__and3_1
X_4082_ _1153_ _1117_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__nor2_1
X_3033_ _2765_ _2769_ ih.t.count\[29\] vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4626__A2 _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4984_ _1969_ _1970_ _1971_ _1799_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__a2bb2o_1
X_3935_ _0986_ _1006_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5339__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5605_ ih.t.timer_max\[20\] _2150_ _2319_ ih.t.timer_max\[4\] _1661_ vssd1 vssd1
+ vccd1 vccd1 _2421_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3866_ _0933_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5147__A _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3797_ cu.reg_file.reg_b\[3\] _0426_ _0429_ cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1
+ vccd1 _0873_ sky130_fd_sc_hd__a22o_1
X_5536_ net85 _1330_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__or2_1
X_5467_ _2292_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
X_4418_ _1473_ _1477_ _1478_ _1356_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__o22ai_1
X_5398_ _1194_ net130 _2237_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__mux2_1
X_4349_ cu.pc.pc_o\[4\] _1322_ _1315_ cu.reg_file.reg_e\[4\] _1412_ vssd1 vssd1 vccd1
+ vccd1 _1413_ sky130_fd_sc_hd__a221o_1
X_6019_ clknet_leaf_6_clk _0057_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4226__A _1293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4553__B2 cu.reg_file.reg_sp\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3008__C ih.t.timer_max\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3720_ _0789_ _0792_ _0795_ _0752_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ cu.reg_file.reg_mem\[7\] _0418_ _0433_ cu.reg_file.reg_a\[7\] vssd1 vssd1
+ vccd1 vccd1 _0727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3582_ cu.reg_file.reg_b\[5\] _0502_ _0499_ cu.reg_file.reg_a\[5\] vssd1 vssd1 vccd1
+ vccd1 _0658_ sky130_fd_sc_hd__a22o_1
X_5321_ _2200_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_1
X_5252_ ih.t.timer_max\[26\] _2157_ _2153_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5183_ _1647_ _2107_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__and2_1
X_4203_ _1270_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4134_ _0956_ _0957_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__nor2_1
X_4065_ _0610_ _1136_ _0652_ _0611_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3807__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3016_ ih.t.timer_max\[12\] _2753_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__or2_2
XFILLER_0_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4480__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4967_ _1954_ _1955_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__nor2_1
XANTENNA__3230__D_N _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4898_ cu.pc.pc_o\[7\] _1892_ _1815_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3918_ _0449_ _0972_ _0990_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__or4_2
XFILLER_0_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3849_ _0876_ _0924_ _0875_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5519_ net31 _1625_ _2148_ net34 vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout153 net159 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
Xfanout164 net197 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_2
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
Xfanout197 net26 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_4
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5515__A _1374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5974__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5870_ _2641_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4821_ _1050_ _1817_ _1795_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5396__S _2237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5962__A0 cu.id.imm_i\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4752_ _2880_ _2913_ _2935_ _0977_ _0350_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4683_ net217 _1705_ _1707_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[16\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3703_ _0512_ _0528_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4517__A1 cu.reg_file.reg_b\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4517__B2 cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3634_ _0704_ _0706_ _0708_ _0709_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5425__A _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6009__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3565_ cu.reg_file.reg_mem\[6\] _0640_ _0433_ cu.reg_file.reg_a\[6\] vssd1 vssd1
+ vccd1 vccd1 _0641_ sky130_fd_sc_hd__a22o_1
X_5304_ _2189_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__clkbuf_1
X_3496_ alu.Cin vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__inv_2
X_6284_ clknet_leaf_36_clk _0266_ net161 vssd1 vssd1 vccd1 vccd1 cu.ir.idx\[0\] sky130_fd_sc_hd__dfrtp_2
X_5235_ _2143_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _2096_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__clkbuf_1
X_4117_ _1160_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__buf_4
X_5097_ _2052_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5245__A2 _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4048_ _1032_ _1121_ _0916_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5999_ clknet_leaf_2_clk _0037_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold9 cu.id.is_halted vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5944__A0 _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5944__S _2666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output97_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3972__B _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3350_ _0425_ _0421_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__nor2_4
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _0354_ _2953_ _0297_ _0356_ _2942_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a2111o_1
X_5020_ _1260_ _1263_ _0368_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__mux2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__A1 cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3486__B2 cu.reg_file.reg_sp\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5922_ _2900_ _2372_ _2668_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5853_ cu.reg_file.reg_sp\[14\] _1287_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4324__A cu.reg_file.reg_l\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4804_ _0306_ _0305_ _1805_ _2950_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o211a_1
X_5784_ cu.reg_file.reg_sp\[6\] _2535_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__nand2_1
X_2996_ net69 vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4735_ _0303_ _0449_ _1743_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4666_ ih.t.count\[10\] ih.t.count\[11\] _1693_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4978__B cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4597_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__clkinv_4
XANTENNA__5163__A1 _1193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3617_ _0294_ _0692_ _0536_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3548_ _0539_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__clkbuf_4
X_6267_ clknet_leaf_23_clk _0249_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_3479_ _0400_ _0546_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__and2_1
X_5218_ _2131_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
X_6198_ clknet_leaf_11_clk net11 net168 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5149_ _2951_ _2004_ _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__and3_1
XANTENNA__4426__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5926__A0 _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4901__A1 cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output135_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5231__C _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3313__A _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5090__A0 cu.reg_file.reg_d\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5674__S _1739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4520_ cu.pc.pc_o\[13\] _1485_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4451_ cu.reg_file.reg_b\[1\] _1313_ _1507_ _1509_ vssd1 vssd1 vccd1 vccd1 _1510_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__5145__A1 cu.reg_file.reg_h\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3402_ _2896_ _0364_ _0477_ _2935_ _2949_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__o2111ai_2
X_4382_ _1382_ _1438_ _1439_ _1444_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__a31o_2
X_6121_ clknet_leaf_21_clk _0155_ net184 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3333_ cu.id.starting_int_service _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ clknet_leaf_22_clk _0090_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5448__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3264_ cu.id.cb_opcode_z\[1\] vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__buf_4
XANTENNA__3459__A1 cu.reg_file.reg_e\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3459__B2 cu.reg_file.reg_b\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ cu.reg_file.reg_a\[1\] _1987_ _1985_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__mux2_1
X_3195_ _2931_ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__buf_2
XANTENNA__5605__C1 _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5081__A0 cu.reg_file.reg_d\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5905_ ih.t.timer_max\[21\] _1191_ _2654_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5620__A2 _2147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3631__A1 cu.pc.pc_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4054__A _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5836_ _1213_ _2615_ _2115_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__mux2_1
X_2979_ net6 vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5767_ cu.reg_file.reg_sp\[4\] _2534_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__nor2_1
X_4718_ ih.t.count\[28\] _1729_ _1670_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__o21ai_1
X_5698_ ih.t.timer_max\[29\] _2151_ _2320_ ih.t.timer_max\[13\] vssd1 vssd1 vccd1
+ vccd1 _2505_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4649_ _1683_ _1684_ _1672_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5136__A1 cu.reg_file.reg_h\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4895__A0 _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4229__A _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3133__A _2870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2972__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3622__A1 cu.reg_file.reg_c\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3622__B2 cu.reg_file.reg_e\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5375__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5127__A1 cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3027__B ih.t.timer_max\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _2951_ _0368_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nand2_4
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3613__B2 cu.reg_file.reg_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3882_ _0950_ _0956_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5621_ net81 _1633_ _2432_ _2435_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5552_ _1649_ _2370_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4503_ cu.pc.pc_o\[12\] _1321_ _1314_ cu.reg_file.reg_d\[4\] _1558_ vssd1 vssd1 vccd1
+ vccd1 _1559_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483_ _2304_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3218__A _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4434_ cu.pc.pc_o\[8\] _1321_ _1314_ cu.reg_file.reg_d\[0\] _1493_ vssd1 vssd1 vccd1
+ vccd1 _1494_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4365_ _1271_ _1427_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__nor2_1
Xwire7 _2895_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6104_ clknet_leaf_9_clk _0138_ net166 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _2887_ _0391_ _2950_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__o21ai_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4296_ _0341_ _1295_ _1298_ cu.pc.pc_o\[2\] _1361_ vssd1 vssd1 vccd1 vccd1 _1362_
+ sky130_fd_sc_hd__a221o_1
X_6035_ clknet_leaf_34_clk _0073_ net163 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3247_ _2878_ _2907_ _2908_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__and3b_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3178_ _2908_ _2914_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__nor2_1
XANTENNA__6276__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5819_ _2599_ _2600_ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5109__A1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4580__A2 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5293__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5596__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5596__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5348__A1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4571__A2 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ss4[0] sky130_fd_sc_hd__buf_2
XFILLER_0_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ss5[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5520__A1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4150_ _0916_ _0940_ _1219_ _0817_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__a2bb2o_1
X_3101_ ih.t.timer_max\[0\] ih.t.timer_max\[1\] ih.t.timer_max\[2\] vssd1 vssd1 vccd1
+ vccd1 _2839_ sky130_fd_sc_hd__o21ai_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 ss1[6] sky130_fd_sc_hd__clkbuf_4
X_4081_ _1153_ _1112_ _1154_ _0610_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__a2bb2o_1
X_3032_ ih.t.count\[29\] _2765_ _2769_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__and3_1
X_4983_ _1624_ _1965_ _1795_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3934_ _1007_ _0981_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3865_ _0939_ _0940_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__nand2_1
X_5604_ _1400_ _2419_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__and2b_1
XANTENNA__5428__A _2139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3796_ cu.reg_file.reg_sp\[11\] _0636_ _0748_ cu.reg_file.reg_h\[3\] vssd1 vssd1
+ vccd1 vccd1 _0872_ sky130_fd_sc_hd__a22o_1
X_5535_ net93 _2194_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5466_ net62 _2085_ _2291_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4417_ _1460_ _1473_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__nand2_1
XANTENNA__5511__A1 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5511__B2 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5397_ _2243_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5192__C_N _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4348_ cu.reg_file.reg_sp\[4\] _0993_ _1344_ _0374_ _1364_ vssd1 vssd1 vccd1 vccd1
+ _1412_ sky130_fd_sc_hd__a221o_1
X_4279_ cu.pc.pc_o\[1\] _1322_ _1315_ cu.reg_file.reg_e\[1\] _1345_ vssd1 vssd1 vccd1
+ vccd1 _1346_ sky130_fd_sc_hd__a221o_1
X_6018_ clknet_leaf_31_clk _0056_ net185 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_d\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4538__C1 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4553__A2 _1282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5502__A1 ih.t.timer_max\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5266__A0 _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3816__A1 cu.id.imm_i\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5012__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ cu.reg_file.reg_c\[7\] _0427_ _0430_ cu.reg_file.reg_e\[7\] vssd1 vssd1 vccd1
+ vccd1 _0726_ sky130_fd_sc_hd__a22o_1
X_3581_ cu.reg_file.reg_d\[5\] _0492_ _0625_ cu.alu_f\[5\] _0656_ vssd1 vssd1 vccd1
+ vccd1 _0657_ sky130_fd_sc_hd__a221o_1
X_5320_ _1190_ net96 _2195_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__mux2_1
X_5251_ _1073_ _1226_ _1667_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4202_ _0294_ _1267_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__or3b_2
X_5182_ mc.cl.next_data\[13\] net23 mc.count vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5257__A0 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4133_ _1201_ _1202_ _1032_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _0719_ _1137_ _1045_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__a21oi_1
X_3015_ ih.t.timer_max\[10\] ih.t.timer_max\[11\] _2752_ vssd1 vssd1 vccd1 vccd1 _2753_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3807__B2 cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3807__A1 cu.reg_file.reg_sp\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4480__B2 cu.reg_file.reg_sp\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4480__A1 cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5009__A0 cu.reg_file.reg_a\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4966_ _1233_ cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__and2_1
X_4897_ _1884_ _1891_ _1809_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__mux2_1
X_3917_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3848_ _0882_ _0885_ _0923_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__a21boi_1
XANTENNA__5732__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3779_ _0853_ _0850_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__or2b_1
X_5518_ net33 _2191_ _1374_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5449_ _1335_ _1354_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__nor2_1
XANTENNA__4299__A1 cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4299__B2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5248__A0 _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4936__S _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_4
Xfanout176 net177 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_4
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
XANTENNA__4471__A1 cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4237__A _1304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5531__A _1739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output42_A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820_ _1819_ _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5411__A0 _1188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5962__A1 _2429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4751_ _1300_ _1739_ _1740_ _1759_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4682_ ih.t.count\[16\] _1705_ _1670_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3702_ _0771_ _0773_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__a21o_1
XANTENNA__5714__A1 _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3633_ _2950_ _0341_ _0507_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3564_ _0418_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__clkbuf_8
X_6283_ clknet_leaf_16_clk _0265_ net178 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5478__A0 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5303_ _1194_ net90 _2182_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3495_ _0570_ _0510_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__and2b_1
X_5234_ ih.t.enable _2085_ _2142_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__mux2_1
X_5165_ cu.reg_file.reg_l\[7\] _1260_ _2088_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout196_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4116_ net209 _1186_ _0370_ _1188_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5096_ cu.reg_file.reg_d\[6\] _2051_ _2039_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4047_ _0804_ _0811_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3896__A _2935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5998_ clknet_leaf_2_clk _0036_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4949_ cu.pc.pc_o\[12\] _1929_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5705__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4444__A1 cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4444__B2 cu.reg_file.reg_h\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5944__A1 _2429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5960__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _2918_ _0355_ _2883_ _2940_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__a2bb2o_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5880__A0 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3486__A2 _0495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4435__A1 cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4435__B2 cu.reg_file.reg_b\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5921_ _2669_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4605__A _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5852_ _2629_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
X_4803_ _2939_ _2916_ _2932_ _0331_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5783_ cu.reg_file.reg_sp\[6\] _2535_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2995_ _2714_ _2733_ vssd1 vssd1 vccd1 vccd1 ih.ih.int_f.data_in sky130_fd_sc_hd__nand2_1
XFILLER_0_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4734_ _2939_ _2916_ _2878_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ net215 _1693_ _1695_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[10\] sky130_fd_sc_hd__a21oi_1
X_4596_ _1629_ _1639_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3616_ cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3547_ cu.reg_file.reg_c\[6\] _0485_ _0622_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__a21o_1
X_6266_ clknet_leaf_23_clk _0248_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3478_ _0514_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__nor2_1
XANTENNA__5871__A0 _2163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5171__A _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5217_ _1188_ ih.gpio_interrupt_mask\[3\] _2127_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__mux2_1
X_6197_ clknet_leaf_11_clk net10 net168 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5148_ _2023_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__inv_2
X_5079_ _2040_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4426__B2 cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4426__A1 cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5926__A1 _2410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4250__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3313__B cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output128_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__A0 cu.reg_file.reg_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4425__A _1269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5020__S _0368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4450_ cu.pc.pc_o\[9\] _1322_ _1315_ cu.reg_file.reg_d\[1\] _1508_ vssd1 vssd1 vccd1
+ vccd1 _1509_ sky130_fd_sc_hd__a221o_1
X_4381_ _1353_ _1434_ _1443_ _1371_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__a22o_1
X_3401_ _2902_ _0300_ _2912_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6120_ clknet_leaf_13_clk _0154_ net173 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3332_ _2877_ _2878_ _2932_ _2925_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ clknet_leaf_22_clk _0089_ net189 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5448__A3 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3263_ _0296_ _0297_ _0337_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__or4_2
XANTENNA__3459__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ cu.id.opcode\[2\] cu.id.opcode\[1\] cu.id.opcode\[6\] cu.id.opcode\[7\] vssd1
+ vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__or4_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _1051_ _1623_ _0368_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5904_ _2659_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4335__A _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3631__A2 _0501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5835_ _2613_ _2614_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4054__B _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2978_ net12 vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5766_ _2554_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
X_4717_ _1729_ _1730_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[27\] sky130_fd_sc_hd__nor2_1
X_5697_ net5 _1650_ _2488_ _2504_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4648_ ih.t.count\[4\] _1679_ ih.t.count\[5\] vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4579_ _2702_ _1194_ _1624_ _2697_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__a22o_1
X_6249_ clknet_leaf_1_clk _0231_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5844__A0 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3308__B _0379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3324__A _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5015__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3950_ _0964_ _1015_ _1016_ _1017_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3881_ _0866_ _0906_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5620_ net113 _2147_ _2225_ net121 _2434_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5551_ net9 _2345_ _2369_ net17 vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4574__B1 _1226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4502_ cu.reg_file.reg_sp\[12\] _0992_ _1343_ cu.id.imm_i\[12\] _1323_ vssd1 vssd1
+ vccd1 vccd1 _1558_ sky130_fd_sc_hd__a221o_1
X_5482_ net66 _0618_ _2303_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4433_ cu.reg_file.reg_sp\[8\] _0992_ _1343_ cu.id.imm_i\[8\] _1323_ vssd1 vssd1
+ vccd1 vccd1 _1493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4364_ cu.reg_file.reg_c\[5\] _1281_ _1426_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__a21oi_1
X_6103_ clknet_leaf_31_clk _0137_ net183 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_4
X_4295_ _1271_ _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__nor2_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _2936_ _0385_ _0386_ _2928_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__a311o_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3234__A _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _2896_ _2911_ _2935_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__nand3_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ clknet_leaf_33_clk _0072_ net163 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_h\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _2912_ _2913_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4801__A1 _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5818_ _2590_ _2593_ _2591_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4512__B _1561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5749_ cu.reg_file.reg_sp\[1\] _2531_ _2539_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3144__A _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2983__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5596__A2 _2236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ss4[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5520__A2 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output72_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 ss0[4] sky130_fd_sc_hd__clkbuf_4
X_3100_ _2836_ ih.t.count\[0\] ih.t.timer_max\[0\] vssd1 vssd1 vccd1 vccd1 _2838_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 ss1[7] sky130_fd_sc_hd__clkbuf_4
X_4080_ _0611_ _0671_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__nand2_1
X_3031_ ih.t.timer_max\[28\] _2764_ ih.t.timer_max\[29\] vssd1 vssd1 vccd1 vccd1 _2769_
+ sky130_fd_sc_hd__o21ai_1
X_4982_ _1966_ _1968_ _1798_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3933_ _0998_ _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3864_ _0877_ _0924_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__xnor2_1
X_5603_ ih.t.timer_max\[12\] _2193_ _2314_ ih.t.timer_max\[4\] _2418_ vssd1 vssd1
+ vccd1 vccd1 _2419_ sky130_fd_sc_hd__a221o_1
XANTENNA__5428__B _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4332__B _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3795_ cu.id.imm_i\[11\] _0739_ _0870_ _0653_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__a22oi_4
X_5534_ net125 _2236_ _2247_ net133 vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5465_ _2290_ _2284_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__nor2_1
XANTENNA__3770__A1 cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3770__B2 cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4416_ _1356_ _1460_ _1402_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__o21a_1
X_5396_ _1192_ net129 _2237_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4347_ cu.reg_file.reg_l\[4\] _1317_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__and2_1
XANTENNA__5275__A1 _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4278_ cu.reg_file.reg_sp\[1\] _0993_ _1344_ _0340_ _1324_ vssd1 vssd1 vccd1 vccd1
+ _1345_ sky130_fd_sc_hd__a221o_1
X_6017_ clknet_leaf_7_clk _0055_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_3229_ _2902_ _2884_ _2875_ _2876_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__or4bb_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2978__A net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3513__A1 cu.reg_file.reg_c\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3513__B2 cu.reg_file.reg_e\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5266__A1 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4417__B _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output110_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_20_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3580_ cu.pc.pc_o\[5\] _0501_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3752__A1 cu.reg_file.reg_a\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3752__B2 cu.reg_file.reg_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5250_ _2156_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4201_ cu.id.state\[1\] cu.id.state\[0\] _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__and3b_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5181_ _2106_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3504__B2 cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4132_ _0942_ _0943_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__or2_1
XANTENNA__5257__A1 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4063_ _0603_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__nand2_1
X_3014_ ih.t.timer_max\[9\] _2751_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__or2_2
XANTENNA__3512__A _0587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4480__A2 _1282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4965_ _1233_ cu.pc.pc_o\[13\] vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3916_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__buf_2
X_4896_ _1889_ _1890_ _1798_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3847_ _0887_ _0922_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__or2_1
X_3778_ _0850_ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__or2b_1
X_5517_ net32 _1330_ _1354_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5174__A _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5448_ net73 net75 net72 net74 _1354_ _1330_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__mux4_1
XANTENNA__4299__A2 _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5379_ _1194_ net122 _2226_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__mux2_1
Xfanout155 net159 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout177 net181 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net196 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout166 net169 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5248__A1 _1623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4428__A _1269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5958__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output35_A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5411__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4750_ _1645_ _1755_ _1758_ _1269_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__o22a_1
XANTENNA__4163__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4681_ _1705_ _1706_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[15\] sky130_fd_sc_hd__nor2_1
X_3701_ _0512_ _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__nor2_2
XANTENNA__3973__B2 _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3632_ cu.reg_file.reg_sp\[2\] _0624_ _0492_ cu.reg_file.reg_d\[2\] _0707_ vssd1
+ vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5302_ _2188_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__clkbuf_1
X_3563_ cu.reg_file.reg_c\[6\] _0427_ _0430_ cu.reg_file.reg_e\[6\] vssd1 vssd1 vccd1
+ vccd1 _0639_ sky130_fd_sc_hd__a22o_1
X_6282_ clknet_leaf_16_clk _0264_ net180 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5478__A1 _0618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3494_ _0569_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__buf_2
X_5233_ _2140_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__nor2_1
XANTENNA__3489__B1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5164_ _2095_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__clkbuf_1
X_4115_ _1187_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__buf_4
X_5095_ _1193_ _1624_ _2035_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4989__B1 _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3354__B1_N _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ _0757_ _0767_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5650__A1 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6018__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5997_ clknet_leaf_2_clk _0035_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4948_ _1938_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3413__B1 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4879_ _0387_ cu.pc.pc_o\[6\] vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5705__A2 _1650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4947__S _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5632__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4248__A _1309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5641__A1 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2991__A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5157__A0 cu.reg_file.reg_l\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5807__A cu.reg_file.reg_sp\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5018__S _1985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5880__A1 ih.t.timer_max\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _2923_ _2350_ _2668_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5851_ cu.reg_file.reg_sp\[14\] _2628_ _2538_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__mux2_1
X_2994_ _2720_ _2726_ _2732_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__and3_1
XANTENNA__5396__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4802_ _1803_ _1742_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5782_ _2568_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4733_ _2893_ _1741_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4664_ ih.t.count\[10\] _1693_ _1670_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4595_ _1373_ _1417_ _1637_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__or4_1
X_3615_ cu.reg_file.reg_sp\[3\] _0539_ _0492_ cu.reg_file.reg_d\[3\] _0690_ vssd1
+ vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__a221o_1
X_3546_ cu.reg_file.reg_e\[6\] _0489_ _0621_ cu.reg_file.reg_l\[6\] vssd1 vssd1 vccd1
+ vccd1 _0622_ sky130_fd_sc_hd__a22o_1
X_6265_ clknet_leaf_18_clk _0247_ net193 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_5216_ _2130_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5320__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3477_ _0400_ _0528_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__or2b_1
XANTENNA__5871__A1 ih.t.timer_max\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6196_ clknet_leaf_10_clk net9 net167 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5147_ _0618_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__clkbuf_4
X_5078_ cu.reg_file.reg_d\[0\] _2036_ _2039_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__mux2_1
XANTENNA__5623__A1 ih.t.timer_max\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4426__A2 _1282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4029_ _0611_ _0729_ _0607_ _0552_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4362__B2 cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4362__A1 cu.reg_file.reg_a\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__A1 _2429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5301__S _2182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4425__B _1484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5917__A2 _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire150 net242 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_1
XFILLER_0_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4380_ _1441_ _1442_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3400_ _0452_ _0303_ _0450_ _0475_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__or4b_1
X_3331_ _0299_ _0329_ _0406_ _2877_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ clknet_leaf_22_clk _0088_ net190 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3262_ _2907_ _2914_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__and2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _2918_ _2919_ _2922_ _2924_ _2929_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__o311a_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _1986_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4616__A _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5903_ ih.t.timer_max\[20\] _1189_ _2654_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5369__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5834_ _2604_ _2607_ _2605_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5447__A _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2977_ net5 vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__inv_2
XANTENNA__4041__B1 _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5765_ cu.reg_file.reg_sp\[3\] _2553_ _2539_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4716_ net231 _1726_ _1687_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__o21ai_1
X_5696_ _2503_ _1643_ cu.reg_file.reg_mem\[12\] _1646_ vssd1 vssd1 vccd1 vccd1 _2504_
+ sky130_fd_sc_hd__a2bb2o_1
X_4647_ ih.t.count\[4\] ih.t.count\[5\] _1679_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _0516_ _1200_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__nor2_4
X_3529_ _0399_ _0546_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__or2_1
X_6248_ clknet_leaf_42_clk _0230_ net152 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_6179_ clknet_leaf_21_clk _0213_ net182 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4804__C1 _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5121__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5780__A0 _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5523__C _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4099__B1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3324__B _0399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5031__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5966__S _2686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3880_ _0951_ _0952_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__or3_1
X_5550_ _1335_ _1372_ _1661_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__and3_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4574__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5481_ _2302_ _2284_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__nor2_1
X_4501_ cu.pc.pc_o\[12\] _1485_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4432_ cu.pc.pc_o\[8\] _1485_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4326__A1 cu.pc.pc_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4326__B2 cu.reg_file.reg_e\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ cu.reg_file.reg_e\[5\] _1283_ _1285_ cu.reg_file.reg_l\[5\] _1425_ vssd1 vssd1
+ vccd1 vccd1 _1426_ sky130_fd_sc_hd__a221o_1
X_6102_ clknet_leaf_13_clk _0136_ net173 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_2
X_4294_ cu.reg_file.reg_c\[2\] _1281_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__a21oi_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _0388_ _0389_ _2918_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__a21oi_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _0318_ _0319_ _0320_ _2913_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__or4b_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ clknet_leaf_4_clk _0071_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _2909_ _2878_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__or2_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5177__A _1647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5817_ _2597_ _2598_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__nand2_1
X_5748_ _2538_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ mc.cl.next_data\[8\] _2359_ _2489_ _2490_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__6285__RESET_B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4150__A1_N _0916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4256__A _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4795__A1_N _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3461__D1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4005__B1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4556__A1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5815__A cu.reg_file.reg_sp\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[2] sky130_fd_sc_hd__buf_2
XANTENNA__5520__A3 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output65_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 ss0[5] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 ss2[0] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5550__A _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3030_ ih.t.timer_max\[31\] _2767_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _1966_ _1968_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3932_ _1004_ _0986_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__and2b_1
XANTENNA__4613__B _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3863_ _0936_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__and2b_1
X_5602_ ih.t.timer_max\[28\] _2146_ _2204_ ih.t.timer_max\[20\] vssd1 vssd1 vccd1
+ vccd1 _2418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5533_ _2352_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
X_3794_ cu.reg_file.reg_a\[3\] _0625_ _0628_ cu.reg_file.reg_mem\[11\] _0869_ vssd1
+ vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5464_ _2194_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__inv_2
XANTENNA__3770__A2 _0488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4415_ _1463_ _1474_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__nand2_1
X_5395_ _2242_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
X_4346_ _0374_ _1295_ _1298_ cu.pc.pc_o\[4\] _1409_ vssd1 vssd1 vccd1 vccd1 _1410_
+ sky130_fd_sc_hd__a221o_2
XANTENNA__5460__A _1369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4277_ _1343_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__buf_2
X_6016_ clknet_leaf_7_clk _0054_ net171 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_3228_ _2936_ _2885_ _2941_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__nand3_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ _2894_ net243 vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__nand2_4
XFILLER_0_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4538__A1 cu.id.imm_i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4538__B2 cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output103_A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4200_ cu.id.state\[2\] vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__buf_2
X_5180_ _1647_ _2105_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__and2_1
X_4131_ _0942_ _0943_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__nand2_1
X_4062_ _0599_ _1100_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__nor2_1
X_3013_ ih.t.timer_max\[7\] ih.t.timer_max\[8\] _2750_ vssd1 vssd1 vccd1 vccd1 _2751_
+ sky130_fd_sc_hd__or3_1
XANTENNA__4465__B1 _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_16_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4624__A _1665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ cu.pc.pc_o\[13\] _1939_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3915_ _0295_ _0968_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__or2_1
X_4895_ _1110_ _1884_ _1794_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3846_ _0920_ _0896_ _0796_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3777_ cu.reg_file.reg_mem\[13\] _0640_ _0851_ _0852_ vssd1 vssd1 vccd1 vccd1 _0853_
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__5455__A _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5516_ _1369_ _2331_ _2332_ _2335_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__o31a_1
X_5447_ _1417_ _2136_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5378_ _2232_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4329_ _1376_ _1393_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__or2_1
Xfanout156 net159 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_4
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_4
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
Xfanout167 net168 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A0 cu.id.imm_i\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5708__B1 cu.reg_file.reg_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2989__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4428__B _1484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3670__A1 cu.reg_file.reg_a\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3700_ _0774_ _0775_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__nand2_4
X_4680_ net235 _1702_ _1687_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3631_ cu.pc.pc_o\[2\] _0501_ _0502_ cu.reg_file.reg_b\[2\] _0536_ vssd1 vssd1 vccd1
+ vccd1 _0707_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3562_ cu.reg_file.reg_sp\[6\] _0636_ _0419_ cu.reg_file.reg_h\[6\] _0637_ vssd1
+ vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__a221o_1
X_5301_ _1192_ net89 _2182_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__mux2_1
X_6281_ clknet_leaf_17_clk _0263_ net178 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3493_ _0519_ _0553_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__or2_1
X_5232_ _1364_ _1631_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_5_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5163_ cu.reg_file.reg_l\[6\] _1193_ _2088_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__mux2_1
X_4114_ _1089_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3523__A _0598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5094_ _2050_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4989__A1 cu.pc.pc_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4045_ _0606_ _0643_ _0663_ _0822_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__a221o_1
XANTENNA__5650__A2 _1648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5938__A0 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5996_ clknet_leaf_2_clk _0034_ net155 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5884__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4947_ cu.pc.pc_o\[11\] _1937_ _1814_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__mux2_1
X_4878_ _1872_ _1873_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _0871_ _0874_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5124__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3101__B1 ih.t.timer_max\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5641__A2 _1633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3652__A1 cu.reg_file.reg_l\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4601__B1 _1644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5157__A1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5823__A cu.reg_file.reg_sp\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5034__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3343__A _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3891__B2 _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5093__A0 cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap1 _2324_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5850_ _1624_ _2627_ _2115_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ _2727_ ih.ih.ih.prev_data\[0\] _2728_ ih.ih.ih.prev_data\[15\] _2731_ vssd1
+ vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__o221a_1
XANTENNA__5396__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4801_ _2923_ _2899_ _2879_ _0314_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__o311a_1
X_5781_ cu.reg_file.reg_sp\[5\] _2567_ _2539_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__mux2_1
X_4732_ cu.alu_f\[6\] alu.Cin _0359_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__mux2_1
X_4663_ _1693_ _1694_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[9\] sky130_fd_sc_hd__nor2_1
XANTENNA__5717__B _2351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3614_ cu.pc.pc_o\[3\] _0501_ _0502_ cu.reg_file.reg_b\[3\] _0536_ vssd1 vssd1 vccd1
+ vccd1 _0690_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4594_ _1329_ _1372_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__nor2_1
X_3545_ _0464_ _0487_ _0482_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__o21a_1
X_6264_ clknet_leaf_23_clk _0246_ net192 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_3476_ _0528_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__nor2_1
XANTENNA__4659__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5215_ _1075_ ih.gpio_interrupt_mask\[2\] _2127_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__mux2_1
XANTENNA__5320__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6195_ clknet_leaf_7_clk net2 net171 vssd1 vssd1 vccd1 vccd1 ih.ih.ih.prev_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5146_ _2084_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__clkbuf_1
X_5077_ _2035_ _2038_ _2951_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__o21a_4
X_4028_ _0599_ _1101_ _0610_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5979_ clknet_leaf_30_clk _0017_ net187 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5139__A1 cu.reg_file.reg_h\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4531__B _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4898__A0 cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4250__C _2923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4441__B _1496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5029__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3338__A _0293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output95_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _2889_ _2933_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__or2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5000_ cu.reg_file.reg_a\[0\] _1983_ _1985_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__mux2_1
X_3261_ _0302_ _0303_ _0317_ _0336_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__o31a_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3192_ _2926_ _2928_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__nor2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5902_ _2658_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5833_ _2611_ _2612_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2976_ net14 vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5764_ _1089_ _2552_ _2545_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__mux2_1
X_4715_ ih.t.count\[27\] _1726_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__and2_1
X_5695_ mc.cl.next_data\[12\] _2359_ _2490_ _2502_ vssd1 vssd1 vccd1 vccd1 _2503_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4646_ net220 _1679_ _1682_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[4\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4577_ _2702_ _1192_ _1209_ _2697_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__a22o_1
X_6316_ clknet_leaf_37_clk _0002_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.is_interrupted
+ sky130_fd_sc_hd__dfrtp_1
X_3528_ _0447_ _0601_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__mux2_1
X_6247_ clknet_leaf_1_clk _0229_ net152 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3459_ cu.reg_file.reg_e\[1\] _0488_ _0502_ cu.reg_file.reg_b\[1\] _0534_ vssd1 vssd1
+ vccd1 vccd1 _0535_ sky130_fd_sc_hd__a221o_1
X_6178_ clknet_leaf_21_clk _0212_ net182 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_5129_ _1226_ _1073_ _2066_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__mux2_1
XANTENNA__6073__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4807__A _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4526__B _1579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6002__RESET_B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4280__A1 cu.reg_file.reg_c\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5638__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5532__A1 _2350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output133_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5312__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5599__B2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4271__A1 cu.reg_file.reg_e\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4271__B2 cu.reg_file.reg_l\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3068__A ih.t.timer_max\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__A2 _1075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5480_ _2236_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__inv_2
X_4500_ _1296_ _1554_ _1555_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4431_ _1296_ _1487_ _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_1 _0728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4362_ cu.reg_file.reg_a\[5\] _1276_ _1287_ cu.reg_file.reg_sp\[5\] vssd1 vssd1 vccd1
+ vccd1 _1425_ sky130_fd_sc_hd__a22o_1
X_6101_ clknet_leaf_28_clk _0135_ net186 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _0374_ cu.id.cb_opcode_x\[1\] cu.id.cb_opcode_x\[0\] vssd1 vssd1 vccd1 vccd1
+ _0389_ sky130_fd_sc_hd__or3_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ cu.reg_file.reg_e\[2\] _1283_ _1285_ cu.reg_file.reg_l\[2\] _1358_ vssd1 vssd1
+ vccd1 vccd1 _1359_ sky130_fd_sc_hd__a221o_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _2884_ net151 _2934_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__and3b_2
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ clknet_leaf_4_clk _0070_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3175_ _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout164_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5211__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5816_ cu.reg_file.reg_sp\[10\] _2536_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__nand2_1
XANTENNA__5892__S _2645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2959_ mc.rw.state\[0\] mc.rw.state\[2\] _2695_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5762__A1 cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5747_ _0740_ _2116_ _2537_ _2948_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__o31a_2
XFILLER_0_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5678_ _1489_ _1631_ _1661_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__or3_2
XANTENNA__5514__A1 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4629_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5514__B2 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3706__A _0545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5132__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4971__S _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3764__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5815__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3616__A cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 ss0[6] sky130_fd_sc_hd__clkbuf_4
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 ss2[1] sky130_fd_sc_hd__clkbuf_4
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5831__A cu.reg_file.reg_sp\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5550__B _1372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5977__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5441__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4980_ _1943_ _1955_ _1967_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3931_ _0976_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
X_3862_ _0923_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5601_ net80 _1633_ _2413_ _2416_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3793_ cu.pc.pc_o\[11\] _0740_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5532_ cu.reg_file.reg_mem\[0\] _2350_ _2351_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3755__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5463_ _2289_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
X_4414_ _1463_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__or2_1
X_5394_ _1190_ net128 _2237_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__mux2_1
X_4345_ _1271_ _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4276_ _0295_ _1318_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nor2_2
XANTENNA__4483__A1 _1296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6015_ clknet_leaf_7_clk _0053_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_3227_ _2916_ _2917_ _2919_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__and3b_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3158_ cu.id.opcode\[2\] cu.id.opcode\[6\] cu.id.opcode\[7\] cu.id.opcode\[1\] vssd1
+ vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3089_ _2751_ _2825_ ih.t.count\[8\] vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5432__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5188__A _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5127__S _2069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5423__A0 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5726__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5037__S _2002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4130_ _0777_ _0949_ _1197_ _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__a22o_1
X_4061_ _1131_ _1134_ _0517_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__o21a_1
X_3012_ ih.t.timer_max\[5\] ih.t.timer_max\[6\] _2749_ vssd1 vssd1 vccd1 vccd1 _2750_
+ sky130_fd_sc_hd__or3_2
XANTENNA__4465__B2 cu.reg_file.reg_h\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4905__A cu.id.cb_opcode_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ _1952_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3914_ _2936_ _0386_ _0312_ _0323_ _0984_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a2111o_1
X_4894_ _1887_ _1888_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3845_ _0895_ _0892_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3776_ cu.reg_file.reg_b\[5\] _0426_ _0429_ cu.reg_file.reg_d\[5\] vssd1 vssd1 vccd1
+ vccd1 _0852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5515_ _1374_ _2333_ _2334_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5446_ _1640_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__buf_2
XANTENNA__4153__B1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5377_ _1192_ net121 _2226_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4328_ _1387_ _1388_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__o21a_2
Xfanout179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_4
X_4259_ cu.reg_file.reg_e\[0\] _1315_ _1317_ cu.reg_file.reg_l\[0\] _1326_ vssd1 vssd1
+ vccd1 vccd1 _1327_ sky130_fd_sc_hd__a221o_1
XANTENNA__3703__B _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4087__A _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net159 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5405__A0 _0619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A1 _2372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5708__B2 _1646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5892__A0 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__B2 cu.pc.pc_o\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__A1 cu.id.imm_i\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5320__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3630_ cu.alu_f\[2\] _0498_ _0628_ cu.reg_file.reg_mem\[2\] _0705_ vssd1 vssd1 vccd1
+ vccd1 _0706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3561_ cu.reg_file.reg_d\[6\] _0415_ _0432_ cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1
+ vccd1 _0637_ sky130_fd_sc_hd__a22o_1
XANTENNA__3076__A ih.t.timer_max\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5300_ _2187_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
X_6280_ clknet_leaf_16_clk _0262_ net178 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3492_ net143 _0532_ _0545_ _0558_ _0567_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__a221o_1
X_5231_ _1367_ _1625_ _2139_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__or3_2
XFILLER_0_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5162_ _2094_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5992__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5093_ cu.reg_file.reg_d\[5\] _2049_ _2039_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__mux2_1
X_4113_ _2946_ _2947_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__or2_2
XFILLER_0_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4044_ _1113_ _1117_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__nor2_1
XANTENNA__4635__A _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5938__A1 _2372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3949__B1 alu.Cin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5995_ clknet_leaf_2_clk _0033_ net154 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4946_ _1931_ _1936_ _1808_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__mux2_1
X_4877_ cu.pc.pc_o\[6\] _1860_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3828_ _0887_ _0901_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3759_ cu.reg_file.reg_b\[6\] _0743_ _0624_ cu.reg_file.reg_sp\[14\] vssd1 vssd1
+ vccd1 vccd1 _0835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5405__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _2022_ net70 _2262_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__mux2_1
XANTENNA__3101__A1 ih.t.timer_max\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4601__A1 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3168__A1 _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5865__A0 _2157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5823__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3340__A1 cu.reg_file.reg_sp\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3340__B2 cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output40_A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5050__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4800_ _2932_ _0330_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2992_ _2729_ ih.ih.ih.prev_data\[7\] _2730_ ih.ih.ih.prev_data\[8\] vssd1 vssd1
+ vccd1 vccd1 _2731_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5780_ _1144_ _2566_ _2545_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4731_ _2946_ _1301_ _1300_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4662_ net226 _1691_ _1687_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3613_ cu.alu_f\[3\] _0498_ _0494_ cu.reg_file.reg_mem\[3\] _0688_ vssd1 vssd1 vccd1
+ vccd1 _0689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4593_ _1434_ _1635_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__nand2_1
X_3544_ _0377_ _0393_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6263_ clknet_leaf_23_clk _0245_ net191 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3475_ _0399_ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5214_ _2129_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5856__A0 _1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6194_ clknet_leaf_35_clk net1 net162 vssd1 vssd1 vccd1 vccd1 ih.ip_ed.prev_data
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3331__B2 _2877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5145_ _2083_ cu.reg_file.reg_h\[7\] _2069_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__mux2_1
X_5076_ _0367_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4027_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__inv_2
X_5978_ clknet_leaf_30_clk _0016_ net188 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4929_ cu.pc.pc_o\[9\] cu.pc.pc_o\[8\] _1233_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5544__C1 _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5135__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4275__A cu.reg_file.reg_l\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3352__A_N _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output88_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3561__A1 cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3561__B2 cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__buf_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _2888_ _2889_ _2927_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__and3_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5066__A1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4185__A _0387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5901_ ih.t.timer_max\[19\] _1187_ _2654_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3589__C_N _0374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5832_ cu.reg_file.reg_sp\[12\] _2536_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__nand2_1
XANTENNA__3845__A_N _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6301__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5763_ _2550_ _2551_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__xor2_1
XANTENNA__4577__B1 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4714_ _1728_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[26\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2975_ _2709_ ih.ih.ih.prev_data\[1\] _2710_ net233 _2713_ vssd1 vssd1 vccd1 vccd1
+ _2714_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3529__A _0399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5694_ ih.t.timer_max\[28\] _2151_ _2320_ ih.t.timer_max\[12\] vssd1 vssd1 vccd1
+ vccd1 _2502_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4645_ ih.t.count\[4\] _1679_ _1670_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4576_ _2702_ _1190_ _1213_ _2697_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__a22o_1
X_3527_ _0548_ _0602_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nor2_2
X_6315_ clknet_leaf_37_clk _0003_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.starting_int_service
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5829__A0 cu.reg_file.reg_sp\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4079__B _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6246_ clknet_leaf_3_clk _0228_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_33_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3458_ cu.pc.pc_o\[1\] _0501_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__and2_1
X_6177_ clknet_leaf_21_clk _0211_ net182 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_3389_ _2892_ _2897_ net151 vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__and3_1
X_5128_ _2072_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4095__A _0566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5059_ _2027_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5638__B _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3791__B2 cu.reg_file.reg_sp\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3791__A1 cu.reg_file.reg_b\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2997__B net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5599__A2 _2205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output126_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4733__A _2893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3349__A _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3782__A1 cu.reg_file.reg_b\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3782__B2 cu.reg_file.reg_sp\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ cu.id.imm_i\[8\] _1294_ _1297_ cu.pc.pc_o\[8\] _1489_ vssd1 vssd1 vccd1 vccd1
+ _1490_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_2 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3084__A ih.t.timer_max\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4361_ _1415_ _1416_ _1418_ _1424_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__a211o_1
X_6100_ clknet_leaf_21_clk _0134_ net182 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ cu.id.cb_opcode_x\[1\] _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__nand2_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4292_ cu.reg_file.reg_a\[2\] _1276_ _1286_ cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1
+ vccd1 _1358_ sky130_fd_sc_hd__a22o_1
X_3243_ _2892_ _2884_ net151 _2897_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__o211a_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ clknet_leaf_2_clk _0069_ net155 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3174_ _2909_ _2910_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5739__A cu.reg_file.reg_sp\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout157_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5815_ cu.reg_file.reg_sp\[10\] _2536_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2958_ _2695_ mc.rw.state\[0\] vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__nor2_2
X_5746_ _0986_ _2532_ _2536_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5677_ ih.t.timer_max\[24\] _2151_ _2320_ ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1
+ _2489_ sky130_fd_sc_hd__a22oi_1
XANTENNA__3773__B2 cu.reg_file.reg_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3773__A1 cu.reg_file.reg_a\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4970__A0 _1209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4628_ ih.t.enable _2869_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3706__B _0600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4559_ cu.pc.pc_o\[15\] _1321_ _1314_ cu.reg_file.reg_d\[7\] _1611_ vssd1 vssd1 vccd1
+ vccd1 _1612_ sky130_fd_sc_hd__a221o_1
X_6229_ clknet_leaf_17_clk ih.t.next_count\[17\] net178 vssd1 vssd1 vccd1 vccd1 ih.t.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4818__A _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5413__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3441__B _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5450__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5450__B2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3764__B2 cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3764__A1 cu.reg_file.reg_b\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3516__A1 cu.reg_file.reg_b\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3516__B2 cu.reg_file.reg_a\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 memory_address_out[9] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 ss2[2] sky130_fd_sc_hd__clkbuf_4
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[4] sky130_fd_sc_hd__buf_2
XANTENNA__5831__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 ss0[7] sky130_fd_sc_hd__buf_2
XANTENNA__4728__A _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5550__C _1661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4492__A2 _1530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5441__A1 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4463__A cu.pc.pc_o\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3930_ _0999_ _0997_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _0887_ _0922_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ net112 _2147_ _2225_ net120 _2415_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__a221o_1
X_3792_ cu.reg_file.reg_d\[3\] _0488_ _0741_ cu.reg_file.reg_h\[3\] _0867_ vssd1 vssd1
+ vccd1 vccd1 _0868_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4952__A0 _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5531_ _1739_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5462_ net61 _2085_ _2288_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4413_ _1332_ _1473_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__xnor2_1
X_5393_ _2241_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
X_4344_ cu.reg_file.reg_c\[4\] _1281_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3542__A _0617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6014_ clknet_leaf_6_clk _0052_ net171 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_4275_ cu.reg_file.reg_l\[1\] _1317_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__and2_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _0300_ _0301_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__nor2_1
X_3157_ cu.id.opcode\[0\] vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3088_ ih.t.count\[8\] _2751_ _2825_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__and3_1
XANTENNA__5432__A1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5729_ _2518_ mc.cl.next_data\[3\] _2111_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5671__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__B2 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5423__A1 _2085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4283__A _1335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5318__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output70_A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4060_ _1120_ _0773_ _1132_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__a31o_1
X_3011_ _2748_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5662__B2 ih.t.timer_max\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3673__B1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5289__A _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4905__B cu.pc.pc_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4962_ cu.pc.pc_o\[12\] _1951_ _1814_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__mux2_1
X_4893_ _1875_ _1878_ _1876_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__o21a_1
X_3913_ _0966_ _0971_ _0987_ _0988_ _0296_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a41o_2
XFILLER_0_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3844_ _0747_ _0751_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3775_ cu.reg_file.reg_sp\[13\] _0636_ _0748_ cu.reg_file.reg_h\[5\] vssd1 vssd1
+ vccd1 vccd1 _0851_ sky130_fd_sc_hd__a22o_1
X_5514_ net63 _1638_ _2279_ net62 vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5445_ _2273_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5350__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5752__A cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5376_ _2231_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
X_4327_ cu.reg_file.reg_c\[3\] _1313_ _1389_ _1391_ vssd1 vssd1 vccd1 vccd1 _1392_
+ sky130_fd_sc_hd__a211o_1
Xfanout169 net181 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_4
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4087__B _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5102__B1 _2951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4258_ cu.reg_file.reg_sp\[0\] _0993_ _1322_ _1299_ _1325_ vssd1 vssd1 vccd1 vccd1
+ _1326_ sky130_fd_sc_hd__a221o_1
X_3209_ cu.id.state\[2\] vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__inv_2
X_4189_ _1194_ _1258_ _1027_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__mux2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5405__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4550__B _1598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__A _0373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5138__S _2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4392__A1 cu.reg_file.reg_c\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5341__A0 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__A _0412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5580__B1 _2225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ _0413_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5572__A _1649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5230_ _2138_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__buf_2
X_3491_ _0566_ _0547_ _0550_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5161_ cu.reg_file.reg_l\[5\] _1191_ _2088_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__mux2_1
XANTENNA__3477__B_N _0528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5092_ _1191_ _1209_ _2035_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__mux2_1
X_4112_ _1027_ _1075_ _1183_ _1185_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4043_ _0588_ _1059_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__or2_1
XANTENNA__3820__A _0892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5994_ clknet_leaf_2_clk _0032_ net155 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_a\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4354__C _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4945_ _1934_ _1935_ _1798_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4876_ cu.pc.pc_o\[6\] _1860_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3827_ _0902_ _0885_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__nor2_1
X_3758_ cu.reg_file.reg_d\[6\] _0488_ _0741_ cu.reg_file.reg_h\[6\] vssd1 vssd1 vccd1
+ vccd1 _0834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3689_ _0761_ _0764_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__nor2_1
XANTENNA__6067__RESET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5428_ _2139_ _2194_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__nand2_1
X_5359_ _2221_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3714__B _0632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3885__B1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5626__A1 _1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4826__A _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3101__A2 ih.t.timer_max\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__B _1598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4601__A2 _1489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5314__A0 _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3905__A _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5865__A1 ih.t.timer_max\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2999__A_N net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5617__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5331__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap3 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2991_ net16 vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4730_ _1364_ _1489_ _1644_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__a21oi_4
X_4661_ ih.t.count\[8\] ih.t.count\[9\] _1689_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3612_ cu.reg_file.reg_h\[3\] _0495_ _0499_ cu.reg_file.reg_a\[3\] vssd1 vssd1 vccd1
+ vccd1 _0688_ sky130_fd_sc_hd__a22o_1
X_4592_ _1434_ _1629_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__or3b_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3543_ _0618_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6262_ clknet_leaf_23_clk _0244_ net193 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5305__A0 _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3474_ _0392_ _0384_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__and2b_1
X_5213_ _1052_ ih.gpio_interrupt_mask\[1\] _2127_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__mux2_1
X_6193_ clknet_leaf_22_clk _0226_ net196 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5144_ _1263_ _1110_ _2066_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout187_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5075_ _0352_ _1790_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4026_ _1060_ _0588_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4292__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5977_ clknet_leaf_33_clk _0014_ net163 vssd1 vssd1 vccd1 vccd1 cu.alu_f\[7\] sky130_fd_sc_hd__dfrtp_1
X_4928_ _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4859_ _1855_ _1856_ _1799_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3725__A _0733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5326__S _2195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3635__A _0587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3190_ _2902_ cu.id.alu_opcode\[3\] vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5900_ _2657_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5831_ cu.reg_file.reg_sp\[12\] _2536_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__or2_1
X_2974_ _2711_ ih.ih.ih.prev_data\[2\] _2712_ ih.ih.ih.prev_data\[3\] vssd1 vssd1
+ vccd1 vccd1 _2713_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5762_ cu.reg_file.reg_sp\[1\] _2543_ _2541_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4577__B2 _2697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4577__A1 _2702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4713_ _1726_ _1727_ _1669_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5693_ net4 _1650_ _2488_ _2501_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__a31o_1
X_4644_ _1681_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4575_ _2702_ _1188_ _1222_ _2697_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__a22o_1
XANTENNA__5236__S _1667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3526_ _0519_ _0555_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__or2b_2
X_6314_ clknet_leaf_37_clk net201 net161 vssd1 vssd1 vccd1 vccd1 cu.id.is_halted sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6245_ clknet_leaf_3_clk _0227_ net156 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_sp\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5760__A cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3457_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[1\] vssd1 vssd1 vccd1 vccd1 _0533_
+ sky130_fd_sc_hd__o211a_1
X_6176_ clknet_leaf_21_clk _0210_ net184 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4501__A1 cu.pc.pc_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3388_ _0458_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__nor2_2
X_5127_ _2071_ cu.reg_file.reg_h\[1\] _2069_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__mux2_1
X_5058_ cu.reg_file.reg_c\[1\] _1051_ _2025_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__mux2_1
X_4009_ _0600_ _1041_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_1
XANTENNA__4095__B _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5765__A0 cu.reg_file.reg_sp\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3791__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4985__S _1808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output119_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4559__A1 cu.pc.pc_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5756__A0 _1073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3782__A2 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ _1351_ _1422_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5056__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3311_ cu.id.cb_opcode_x\[0\] vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__buf_4
X_4291_ _1350_ _1352_ _1353_ _1354_ _1357_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__a221o_4
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ clknet_leaf_5_clk _0068_ net158 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_e\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_3242_ _2938_ _2931_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nor2_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _2900_ _2899_ vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__or2b_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5747__B1 _2948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5814_ _2596_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2957_ mc.rw.state\[2\] vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5745_ _2535_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5676_ _1641_ _2344_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__nor2_2
X_4627_ _2706_ _1664_ _1668_ _1647_ _1371_ vssd1 vssd1 vccd1 vccd1 mc.rw.next_state\[2\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4558_ cu.reg_file.reg_sp\[15\] _0992_ _1343_ cu.id.imm_i\[15\] _1323_ vssd1 vssd1
+ vccd1 vccd1 _1611_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4489_ _1333_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__or2_1
X_3509_ _0582_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__nand2_1
X_6228_ clknet_leaf_17_clk ih.t.next_count\[16\] net178 vssd1 vssd1 vccd1 vccd1 ih.t.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ clknet_leaf_20_clk _0193_ net172 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4818__B _1299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3461__A1 cu.reg_file.reg_c\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3764__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3185__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 memory_data_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 memory_address_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ss1[0] sky130_fd_sc_hd__clkbuf_4
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[5] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[2] sky130_fd_sc_hd__clkbuf_4
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ss2[3] sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_28_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ _0813_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__or2b_1
X_3791_ cu.reg_file.reg_b\[3\] _0743_ _0624_ cu.reg_file.reg_sp\[11\] vssd1 vssd1
+ vccd1 vccd1 _0867_ sky130_fd_sc_hd__a22o_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _2329_ _2330_ _2343_ _2349_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__o31a_2
XANTENNA__3755__A2 _0426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5461_ _2287_ _2284_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4412_ _1467_ _1468_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__o21ai_4
X_5392_ _1188_ net127 _2237_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4343_ cu.reg_file.reg_e\[4\] _1283_ _1285_ cu.reg_file.reg_l\[4\] _1406_ vssd1 vssd1
+ vccd1 vccd1 _1407_ sky130_fd_sc_hd__a221o_1
X_4274_ _0340_ _1295_ _1298_ cu.pc.pc_o\[1\] _1305_ vssd1 vssd1 vccd1 vccd1 _1341_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3823__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5665__C1 _1660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6013_ clknet_leaf_6_clk _0051_ net170 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3225_ _2876_ _2875_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__nand2b_4
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ _2892_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__clkbuf_4
X_3087_ ih.t.timer_max\[7\] _2750_ ih.t.timer_max\[8\] vssd1 vssd1 vccd1 vccd1 _2825_
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_19_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5968__A0 cu.id.imm_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5469__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4373__B _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3708__A_N _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5728_ net20 _2519_ _2524_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__a21o_1
X_3989_ _0558_ _0694_ _0822_ _0545_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5659_ net107 _2204_ _2471_ _1401_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4829__A _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3908__A _2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4698__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4458__B _1511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output63_A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5111__A1 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3010_ ih.t.timer_max\[4\] _2747_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__or2_1
XANTENNA__3673__A1 cu.reg_file.reg_sp\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3673__B2 cu.reg_file.reg_h\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6114__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4961_ _1941_ _1950_ _1808_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__mux2_1
X_4892_ _1885_ _1886_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__and2b_1
X_3912_ _2936_ _2881_ _0469_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3843_ _0832_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3774_ cu.id.imm_i\[13\] _0739_ _0849_ _0653_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__a22oi_4
X_5513_ net60 _2277_ _2179_ net61 vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5444_ _2022_ net75 _2272_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4689__B1 _1687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5375_ _1190_ net120 _2226_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__mux2_1
X_4326_ cu.pc.pc_o\[3\] _1322_ _1315_ cu.reg_file.reg_e\[3\] _1390_ vssd1 vssd1 vccd1
+ vccd1 _1391_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout159 net197 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
XANTENNA__5102__A1 _2035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4257_ _0343_ _2950_ _1319_ _1324_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__a31o_1
X_3208_ _2907_ _2915_ _2930_ _2944_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__o211ai_1
X_4188_ cu.alu_f\[6\] _1256_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4861__A0 cu.pc.pc_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3139_ cu.id.opcode\[7\] vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5419__S _2248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3447__B cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5341__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6196__D net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4993__S _1798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output101_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4368__C1 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5580__B2 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5580__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3357__B _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3490_ _0560_ _0562_ _0564_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__o31a_4
XANTENNA__5853__A cu.reg_file.reg_sp\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5064__S _2025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _2093_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__clkbuf_1
X_5091_ _2048_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
X_4111_ cu.alu_f\[2\] _1184_ _0370_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__a21o_1
XANTENNA__5096__A0 cu.reg_file.reg_d\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4042_ _0531_ _0632_ _0566_ _0558_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__a2bb2o_1
X_5993_ clknet_leaf_29_clk _0031_ net188 vssd1 vssd1 vccd1 vccd1 cu.pc.pc_o\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ _1222_ _1931_ _1794_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__mux2_1
X_4875_ _1871_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5020__A0 _1260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3826_ _0882_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__inv_2
XANTENNA__5571__B2 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5571__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3757_ _0829_ _0832_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3688_ _0716_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5427_ _2261_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _1192_ net113 _2215_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__mux2_1
X_4309_ _1371_ _1372_ _1374_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__a21o_1
XANTENNA__5087__A0 cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5289_ _1364_ _2169_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__nor2_2
XANTENNA__4826__B cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4834__A0 _1073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6036__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4842__A cu.id.cb_opcode_y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3458__A cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5011__A0 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4565__C_N _1598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5314__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5078__A0 cu.reg_file.reg_d\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5617__A2 _2194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3628__B2 cu.reg_file.reg_e\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2990_ net15 vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4660_ _1691_ _1692_ vssd1 vssd1 vccd1 vccd1 ih.t.next_count\[8\] sky130_fd_sc_hd__nor2_1
XFILLER_0_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5002__A0 _1051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3611_ cu.reg_file.reg_c\[3\] _0485_ _0489_ cu.reg_file.reg_e\[3\] _0686_ vssd1 vssd1
+ vccd1 vccd1 _0687_ sky130_fd_sc_hd__a221o_1
X_4591_ _1455_ _1473_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3542_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__buf_4
XANTENNA__3919__A_N _0986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6261_ clknet_leaf_23_clk _0243_ net193 vssd1 vssd1 vccd1 vccd1 ih.t.timer_max\[9\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__5305__A1 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3473_ _0548_ _0393_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6192_ clknet_leaf_22_clk _0225_ net190 vssd1 vssd1 vccd1 vccd1 mc.cl.next_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_5212_ _2128_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3316__B1 _2950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5143_ _2082_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4927__A _2920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5074_ _0617_ _1622_ _2035_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4025_ _1092_ _1098_ _1069_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4292__A1 cu.reg_file.reg_a\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4292__B2 cu.reg_file.reg_sp\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5976_ clknet_leaf_36_clk _0013_ net161 vssd1 vssd1 vccd1 vccd1 cu.alu_f\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__5477__B _2284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4927_ _2920_ _1521_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4858_ _1160_ _1850_ _1795_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3809_ cu.reg_file.reg_mem\[10\] _0640_ _0883_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__5544__B2 ih.t.timer_max\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3555__B1 _0536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4789_ _0350_ _0358_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4572__A _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5535__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4338__A2 _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5299__A0 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3635__B _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4274__A1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4274__B2 cu.pc.pc_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5223__A0 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5830_ _2610_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
X_2973_ net11 vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__inv_2
X_5761_ _2548_ _2549_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__nor2_1
XANTENNA__4577__A2 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4712_ ih.t.count\[24\] ih.t.count\[25\] _1720_ ih.t.count\[26\] vssd1 vssd1 vccd1
+ vccd1 _1727_ sky130_fd_sc_hd__a31o_1
XANTENNA__3098__A ih.t.timer_max\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5692_ _2500_ _1643_ cu.reg_file.reg_mem\[11\] _1646_ vssd1 vssd1 vccd1 vccd1 _2501_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4643_ _1679_ _1680_ _1672_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5526__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4574_ _2702_ _1075_ _1226_ _2697_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__a22o_1
X_6313_ clknet_leaf_37_clk _0006_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3525_ _0575_ _0588_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__and3_1
X_6244_ clknet_leaf_37_clk _0015_ net160 vssd1 vssd1 vccd1 vccd1 cu.id.interrupt_requested
+ sky130_fd_sc_hd__dfrtp_1
X_3456_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__inv_2
X_6175_ clknet_leaf_20_clk _0209_ net182 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_mem\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4501__A2 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3387_ _0336_ _0460_ _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__a21o_1
X_5126_ _1623_ _1050_ _2066_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__mux2_1
X_5057_ _2026_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5462__A0 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4008_ _0570_ _0763_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _2689_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3776__B1 _0429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3528__A0 _0447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3471__A _0399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4559__A2 _1321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5337__S _2206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output93_A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _2877_ _2880_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__nand2_2
X_4290_ _1356_ _1354_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _2943_ _0316_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__nand2_1
XANTENNA__3381__A cu.id.starting_int_service vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5692__B1 cu.reg_file.reg_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3172_ cu.id.opcode\[6\] cu.id.opcode\[7\] vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__or2_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4196__B _1027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5444__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4643__C _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5747__A1 _0740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5813_ cu.reg_file.reg_sp\[9\] _2595_ _2539_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _2696_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__clkbuf_8
X_5744_ _2534_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5675_ _2487_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4626_ _1651_ _1667_ _1657_ _1351_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4557_ cu.pc.pc_o\[15\] _1485_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4488_ _1305_ _1541_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__o21ai_4
X_3508_ cu.id.cb_opcode_y\[2\] _0361_ _0437_ _0341_ _0583_ vssd1 vssd1 vccd1 vccd1
+ _0584_ sky130_fd_sc_hd__a221o_1
X_6227_ clknet_leaf_17_clk ih.t.next_count\[15\] net178 vssd1 vssd1 vccd1 vccd1 ih.t.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4486__A1 cu.pc.pc_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3439_ _0514_ _0400_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__or2b_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ clknet_leaf_20_clk _0192_ net172 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4486__B2 cu.reg_file.reg_d\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ cu.reg_file.reg_e\[3\] _1187_ _2056_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__mux2_1
XANTENNA__5435__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6089_ clknet_leaf_12_clk _0123_ net168 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_4
XANTENNA__5738__A1 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4410__A1 cu.pc.pc_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6199__D net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 memory_address_out[15] sky130_fd_sc_hd__clkbuf_4
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 memory_data_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 ss1[1] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 programmable_gpio_wr[6] sky130_fd_sc_hd__buf_2
XANTENNA__4297__A cu.reg_file.reg_e\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 programmable_gpio_out[3] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 ss2[4] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5426__A0 _2022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output131_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__inv_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5460_ _1369_ _2179_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4411_ cu.reg_file.reg_c\[7\] _1313_ _1469_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__4165__B1 _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5901__A1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5391_ _2240_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4342_ cu.reg_file.reg_a\[4\] _1276_ _1287_ cu.reg_file.reg_sp\[4\] vssd1 vssd1 vccd1
+ vccd1 _1406_ sky130_fd_sc_hd__a22o_1
X_4273_ _1271_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__nor2_1
XANTENNA__4000__A _1073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6012_ clknet_leaf_6_clk _0050_ net171 vssd1 vssd1 vccd1 vccd1 cu.reg_file.reg_c\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4468__A1 _1521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3224_ _0298_ _0299_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__nand2_1
.ends

