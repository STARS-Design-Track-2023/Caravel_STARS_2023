magic
tech sky130A
magscale 1 2
timestamp 1694284114
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 14 2128 19214 17456
<< metal2 >>
rect 1306 19200 1362 20000
rect 4526 19200 4582 20000
rect 7746 19200 7802 20000
rect 10322 19200 10378 20000
rect 13542 19200 13598 20000
rect 16762 19200 16818 20000
rect 19338 19200 19394 20000
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 9034 0 9090 800
rect 11610 0 11666 800
rect 14830 0 14886 800
rect 18050 0 18106 800
<< obsm2 >>
rect 20 19144 1250 19200
rect 1418 19144 4470 19200
rect 4638 19144 7690 19200
rect 7858 19144 10266 19200
rect 10434 19144 13486 19200
rect 13654 19144 16706 19200
rect 16874 19144 19210 19200
rect 20 856 19210 19144
rect 130 711 2538 856
rect 2706 711 5758 856
rect 5926 711 8978 856
rect 9146 711 11554 856
rect 11722 711 14774 856
rect 14942 711 17994 856
rect 18162 711 19210 856
<< metal3 >>
rect 0 19048 800 19168
rect 19200 17008 20000 17128
rect 0 15648 800 15768
rect 19200 13608 20000 13728
rect 0 12248 800 12368
rect 19200 10208 20000 10328
rect 0 9528 800 9648
rect 19200 7488 20000 7608
rect 0 6128 800 6248
rect 19200 4088 20000 4208
rect 0 2728 800 2848
rect 19200 688 20000 808
<< obsm3 >>
rect 800 17208 19200 17441
rect 800 16928 19120 17208
rect 800 15848 19200 16928
rect 880 15568 19200 15848
rect 800 13808 19200 15568
rect 800 13528 19120 13808
rect 800 12448 19200 13528
rect 880 12168 19200 12448
rect 800 10408 19200 12168
rect 800 10128 19120 10408
rect 800 9728 19200 10128
rect 880 9448 19200 9728
rect 800 7688 19200 9448
rect 800 7408 19120 7688
rect 800 6328 19200 7408
rect 880 6048 19200 6328
rect 800 4288 19200 6048
rect 800 4008 19120 4288
rect 800 2928 19200 4008
rect 880 2648 19200 2928
rect 800 888 19200 2648
rect 800 715 19120 888
<< metal4 >>
rect 3163 2128 3483 17456
rect 5382 2128 5702 17456
rect 7602 2128 7922 17456
rect 9821 2128 10141 17456
rect 12041 2128 12361 17456
rect 14260 2128 14580 17456
rect 16480 2128 16800 17456
rect 18699 2128 19019 17456
<< labels >>
rlabel metal3 s 0 2728 800 2848 6 clk
port 1 nsew signal input
rlabel metal3 s 19200 4088 20000 4208 6 in[0]
port 2 nsew signal input
rlabel metal2 s 13542 19200 13598 20000 6 in[1]
port 3 nsew signal input
rlabel metal2 s 4526 19200 4582 20000 6 in[2]
port 4 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 in[3]
port 5 nsew signal input
rlabel metal2 s 19338 19200 19394 20000 6 in[4]
port 6 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 in[5]
port 7 nsew signal input
rlabel metal3 s 19200 17008 20000 17128 6 in[6]
port 8 nsew signal input
rlabel metal2 s 16762 19200 16818 20000 6 in[7]
port 9 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 in[8]
port 10 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 in[9]
port 11 nsew signal input
rlabel metal3 s 19200 10208 20000 10328 6 nrst
port 12 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 out[0]
port 13 nsew signal output
rlabel metal2 s 18 0 74 800 6 out[10]
port 14 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 out[11]
port 15 nsew signal output
rlabel metal2 s 7746 19200 7802 20000 6 out[12]
port 16 nsew signal output
rlabel metal3 s 19200 688 20000 808 6 out[13]
port 17 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 out[1]
port 18 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 out[2]
port 19 nsew signal output
rlabel metal3 s 19200 13608 20000 13728 6 out[3]
port 20 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 out[4]
port 21 nsew signal output
rlabel metal2 s 10322 19200 10378 20000 6 out[5]
port 22 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 out[6]
port 23 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 out[7]
port 24 nsew signal output
rlabel metal2 s 1306 19200 1362 20000 6 out[8]
port 25 nsew signal output
rlabel metal3 s 19200 7488 20000 7608 6 out[9]
port 26 nsew signal output
rlabel metal4 s 3163 2128 3483 17456 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 17456 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 17456 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 17456 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 17456 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 17456 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 17456 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 17456 6 vssd1
port 28 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 212514
string GDS_FILE /home/designer-05/Caravel_STARS_2023/openlane/ReducedMacro/runs/23_09_09_11_27/results/signoff/reducedMacroMain.magic.gds
string GDS_START 23764
<< end >>

