* NGSPICE file created from silly_synthesizer.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt silly_synthesizer clk cs gpio[0] gpio[10] gpio[11] gpio[12] gpio[13] gpio[14]
+ gpio[15] gpio[16] gpio[1] gpio[2] gpio[3] gpio[4] gpio[5] gpio[6] gpio[7] gpio[8]
+ gpio[9] nrst pwm vccd1 vssd1
XFILLER_0_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2037_ _0467_ _0472_ _0474_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__o21a_1
X_2106_ _0543_ _0528_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1270_ _0917_ net18 vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2655_ clknet_leaf_18_clk inputs.keypad\[16\] net55 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ clknet_leaf_18_clk net155 net56 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1606_ outputs.scaled_buffer\[5\] _1187_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1537_ _1115_ _1116_ _1117_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__or4_1
X_1468_ _1041_ _1063_ _1065_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__and3_1
X_1399_ _1003_ outputs.sig_gen.count\[1\] outputs.divider_buffer\[13\] _1004_ vssd1
+ vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__a2bb2o_1
X_2586_ clknet_leaf_36_clk net77 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold181 outputs.div.a\[22\] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold170 outputs.div.divisor\[16\] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 inputs.mode_edge.det_edge vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2440_ _0847_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1253_ _0918_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1322_ _0959_ _0960_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[9\]
+ sky130_fd_sc_hd__nor2_1
X_2371_ _0572_ _0791_ _0794_ _0796_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2707_ clknet_leaf_13_clk net97 net58 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_2569_ clknet_leaf_27_clk outputs.sample_rate.next_count\[5\] net30 vssd1 vssd1 vccd1
+ vccd1 outputs.sample_rate.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_2638_ clknet_leaf_26_clk net89 net31 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.octave_key_up
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1940_ outputs.div.q\[25\] _0915_ _0996_ net204 _0418_ vssd1 vssd1 vccd1 vccd1 _0054_
+ sky130_fd_sc_hd__a221o_1
X_1871_ outputs.div.a\[22\] _0355_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2423_ _0838_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1305_ inputs.random_update_clock.count\[16\] inputs.random_update_clock.count\[19\]
+ inputs.random_update_clock.count\[18\] inputs.random_update_clock.count\[17\] vssd1
+ vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__and4bb_1
X_2285_ _0541_ _0689_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__or2_1
X_2354_ _0541_ _0556_ _0754_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1854_ _0359_ _0362_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nand2_1
X_1923_ outputs.div.q\[17\] _0400_ _0405_ net137 _0409_ vssd1 vssd1 vccd1 vccd1 _0046_
+ sky130_fd_sc_hd__a221o_1
X_1785_ _0300_ _0301_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2406_ net232 _0827_ _0798_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2199_ _0585_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__inv_2
X_2337_ _0481_ _0581_ _0748_ _0615_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__a31o_1
X_2268_ _0699_ _0489_ _0494_ _0583_ _0508_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__a41o_1
XFILLER_0_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold52 outputs.signal_buffer2\[13\] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 outputs.signal_buffer2\[12\] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 _0146_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 outputs.signal_buffer2\[1\] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold30 inputs.key_encoder.octave_key_up vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold96 outputs.sample_rate.next_count\[2\] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 inputs.key_encoder.mode_key vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dlygate4sd3_1
X_1570_ _1131_ _1134_ _1139_ _1123_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__and4b_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2053_ _0481_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__buf_2
X_2122_ _0527_ _0557_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1906_ _0914_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_4
X_1837_ _0330_ _0346_ _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1768_ _0248_ _0285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1699_ outputs.div.a\[5\] vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 pwm sky130_fd_sc_hd__buf_2
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2671_ clknet_leaf_20_clk _0017_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2740_ clknet_leaf_22_clk outputs.output_gen.next_count\[7\] net34 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1622_ _1196_ _1197_ _1198_ _1203_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__and4b_1
XFILLER_0_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1484_ _1077_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
X_1553_ _1019_ outputs.shaper.count\[4\] vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nand2_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2036_ _0473_ _0465_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__nand2_1
X_2105_ inputs.key_encoder.sync_keys\[12\] _0526_ _0516_ vssd1 vssd1 vccd1 vccd1 _0543_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2869_ clknet_leaf_34_clk _0187_ net22 vssd1 vssd1 vccd1 vccd1 inputs.frequency_lut.rng\[2\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2723_ clknet_leaf_17_clk net165 net56 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2654_ clknet_leaf_5_clk inputs.keypad\[15\] net44 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1536_ outputs.divider_buffer\[13\] _1110_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__nor2_1
X_1605_ outputs.scaled_buffer\[4\] _1099_ net21 vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__o21ai_1
X_2585_ clknet_leaf_36_clk net93 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1398_ outputs.sig_gen.count\[13\] vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__inv_2
X_1467_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2019_ outputs.div.m\[15\] net239 _0453_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold182 outputs.div.q\[1\] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 outputs.div.q\[2\] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 outputs.div.divisor\[2\] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 inputs.wavetype_fsm.next_state\[1\] vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1252_ _0917_ net2 vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1321_ net213 _0958_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__nor2_1
X_2370_ _1224_ _0737_ _0795_ _0463_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2706_ clknet_leaf_8_clk _0052_ net49 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1519_ outputs.shaper.count\[14\] vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__inv_2
X_2499_ net284 outputs.sig_gen.count\[14\] _0861_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2637_ clknet_leaf_30_clk net134 net32 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2568_ clknet_leaf_28_clk outputs.sample_rate.next_count\[4\] net30 vssd1 vssd1 vccd1
+ vccd1 outputs.sample_rate.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1870_ _0995_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2422_ outputs.divider_buffer\[4\] outputs.div.m\[4\] _0798_ vssd1 vssd1 vccd1 vccd1
+ _0838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2353_ _0774_ _0776_ _0778_ _0779_ _0506_ _0508_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__mux4_1
X_1304_ _0945_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nor2_1
X_2284_ _1199_ _0522_ _0557_ _0566_ _0558_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__a311o_1
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1999_ _0449_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ outputs.div.oscillator_out\[9\] _0398_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1853_ _0359_ _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__or2_1
X_1784_ _0290_ _0292_ _0288_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2336_ _0470_ _0471_ _0731_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a31o_1
X_2405_ _1208_ _0464_ _0556_ _0760_ _0826_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__a41o_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2198_ _0630_ _0632_ _1207_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__mux2_1
X_2267_ _0615_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold42 _0143_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _0144_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 outputs.signal_buffer2\[16\] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 outputs.div.q\[16\] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 inputs.random_note_generator.out\[10\] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 outputs.div.divisor\[6\] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 inputs.keypad_synchronizer.half_sync\[1\] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 outputs.sample_rate.count\[1\] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2052_ _0485_ _0487_ _0489_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__o21ai_1
X_2121_ _0526_ _0522_ _0557_ _0549_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__a311o_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1905_ net189 _0333_ _0377_ net195 _0399_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1836_ _0335_ _0338_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__a21oi_1
X_1767_ outputs.div.m\[11\] outputs.div.m\[10\] _0249_ _0264_ vssd1 vssd1 vccd1 vccd1
+ _0285_ sky130_fd_sc_hd__or4_2
X_1698_ _0205_ _0221_ _0222_ _1228_ net191 vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2319_ _0653_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1552_ outputs.divider_buffer\[4\] _1124_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__or2_1
X_2670_ clknet_leaf_19_clk _0016_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1621_ inputs.key_encoder.sync_keys\[12\] _1199_ _1201_ _1202_ vssd1 vssd1 vccd1
+ vccd1 _1203_ sky130_fd_sc_hd__or4_1
X_1483_ _1041_ _1074_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2104_ _0532_ _0540_ _0541_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2035_ inputs.frequency_lut.rng\[1\] vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__clkbuf_4
X_2868_ clknet_leaf_34_clk _0186_ net22 vssd1 vssd1 vccd1 vccd1 inputs.frequency_lut.rng\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1819_ _0914_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__clkbuf_4
X_2799_ clknet_leaf_1_clk _0117_ net29 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2722_ clknet_leaf_22_clk _0068_ net36 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1535_ outputs.divider_buffer\[12\] _1112_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__nor2_1
X_1604_ outputs.output_gen.count\[5\] _1167_ _1180_ _1184_ _1185_ vssd1 vssd1 vccd1
+ vccd1 _1186_ sky130_fd_sc_hd__o221a_1
X_2584_ clknet_leaf_36_clk net80 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2653_ clknet_leaf_26_clk inputs.keypad\[14\] net31 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1466_ outputs.sig_gen.count\[8\] _1061_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__and2_1
X_1397_ outputs.divider_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2018_ _0459_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold150 inputs.random_update_clock.count\[3\] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _0032_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 outputs.div.divisor\[12\] vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 outputs.output_gen.count\[4\] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 outputs.sample_rate.count\[6\] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1320_ inputs.random_update_clock.count\[9\] inputs.random_update_clock.count\[8\]
+ _0954_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1251_ net1 vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2705_ clknet_leaf_8_clk net179 net49 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2636_ clknet_leaf_25_clk net67 net30 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2498_ _0868_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1518_ _1022_ outputs.shaper.count\[13\] vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__and2_1
X_1449_ _1041_ _1050_ _1051_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__and3_1
X_2567_ clknet_leaf_27_clk outputs.sample_rate.next_count\[3\] net30 vssd1 vssd1 vccd1
+ vccd1 outputs.sample_rate.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1303_ inputs.random_update_clock.count\[9\] inputs.random_update_clock.count\[11\]
+ inputs.random_update_clock.count\[10\] inputs.random_update_clock.count\[8\] vssd1
+ vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__or4bb_1
X_2421_ _0837_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkbuf_1
X_2283_ _0708_ _0710_ _0712_ _0713_ _0616_ _0508_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__mux4_1
X_2352_ _0492_ _0470_ _0467_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1998_ outputs.div.m\[5\] net294 _0436_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__mux2_1
X_2619_ clknet_leaf_28_clk inputs.down.ff_in net32 vssd1 vssd1 vccd1 vccd1 inputs.down.det_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1921_ net137 _0400_ _0405_ net150 _0408_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__a221o_1
X_1852_ _0360_ _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1783_ _0298_ _0299_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2335_ _0586_ _0695_ inputs.frequency_lut.rng\[3\] vssd1 vssd1 vccd1 vccd1 _0763_
+ sky130_fd_sc_hd__o21a_1
X_2266_ _0472_ _0697_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__or2_1
X_2404_ _0603_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__nor2_1
X_2197_ _0599_ _0631_ _0556_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold65 _0147_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _0046_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 outputs.signal_buffer2\[9\] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 outputs.div.q_out\[2\] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 inputs.keypad_synchronizer.half_sync\[0\] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 outputs.signal_buffer2\[4\] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 inputs.random_note_generator.out\[6\] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 inputs.keypad_synchronizer.half_sync\[2\] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 inputs.mode_edge.ff_out vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2120_ _0534_ _0535_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__nor2_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2051_ _0467_ _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1835_ _0335_ _0338_ _0326_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__o21a_1
X_1904_ outputs.div.oscillator_out\[1\] _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1766_ outputs.div.a\[11\] vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__inv_2
X_1697_ _0216_ _0213_ _0220_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__nand3_1
X_2249_ _0548_ _0662_ _1215_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__mux2_1
X_2318_ _0699_ _0744_ _0746_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1482_ _1075_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__inv_2
X_1551_ _1126_ _1132_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1620_ inputs.key_encoder.sync_keys\[4\] inputs.key_encoder.sync_keys\[5\] inputs.key_encoder.sync_keys\[6\]
+ inputs.key_encoder.sync_keys\[7\] vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__or4_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2103_ _1214_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2034_ _0470_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__nand2_2
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1818_ _0328_ _0330_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__nand2_1
X_2798_ clknet_leaf_1_clk _0116_ net29 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2867_ clknet_leaf_34_clk _0185_ net22 vssd1 vssd1 vccd1 vccd1 inputs.frequency_lut.rng\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1749_ _0252_ _0259_ _0260_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__o21ai_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2721_ clknet_leaf_23_clk _0067_ net36 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2652_ clknet_leaf_34_clk inputs.keypad\[13\] net22 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1534_ outputs.divider_buffer\[11\] _1113_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nor2_1
X_1465_ outputs.sig_gen.count\[8\] _1061_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__or2_1
X_1603_ outputs.output_gen.count\[4\] _1183_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__or2_1
X_2583_ clknet_leaf_36_clk net70 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2017_ outputs.div.m\[14\] net230 _0453_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__mux2_1
X_1396_ _1001_ _1002_ vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold140 inputs.random_update_clock.count\[2\] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold151 inputs.random_update_clock.count\[9\] vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 outputs.div.a\[13\] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold184 outputs.div.count\[1\] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 outputs.div.count\[4\] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 outputs.div.q\[0\] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1250_ _0916_ vssd1 vssd1 vccd1 vccd1 outputs.div.next_start sky130_fd_sc_hd__inv_2
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2704_ clknet_leaf_8_clk net142 net48 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2635_ clknet_leaf_33_clk net86 net23 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_2497_ net306 outputs.sig_gen.count\[13\] _0861_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__mux2_1
X_1448_ _1010_ _1047_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__nand2_1
X_1517_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] outputs.scaled_buffer\[3\]
+ outputs.scaled_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__or4_2
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2566_ clknet_leaf_27_clk net158 net31 vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1379_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2420_ outputs.divider_buffer\[3\] outputs.div.m\[3\] _0798_ vssd1 vssd1 vccd1 vccd1
+ _0837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1302_ inputs.random_update_clock.count\[12\] inputs.random_update_clock.count\[15\]
+ inputs.random_update_clock.count\[14\] inputs.random_update_clock.count\[13\] vssd1
+ vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__or4b_1
X_2282_ _0482_ _0472_ _0591_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o21ba_1
X_2351_ _0749_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__nand2_1
X_1997_ _0448_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2549_ _0896_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
X_2618_ clknet_leaf_27_clk inputs.down.in net31 vssd1 vssd1 vccd1 vccd1 inputs.down.ff_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1920_ outputs.div.oscillator_out\[8\] _0398_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__and2_1
X_1851_ outputs.div.a\[19\] _0342_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1782_ _0295_ _0297_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2403_ _0650_ _0823_ _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__mux2_1
X_2334_ _0692_ _0761_ _1224_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__mux2_1
X_2196_ _0532_ _0559_ _1215_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__mux2_1
X_2265_ _0498_ _0467_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold22 inputs.random_note_generator.out\[4\] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 inputs.keypad_synchronizer.half_sync\[11\] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 outputs.signal_buffer2\[14\] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 outputs.div.q\[15\] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 _0140_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 _0071_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 inputs.keypad_synchronizer.half_sync\[10\] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 outputs.signal_buffer2\[0\] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 outputs.sample_rate.count\[5\] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _0486_ _0473_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nor2_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1903_ _0994_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__buf_2
X_1834_ _0328_ _0339_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__or2_1
X_1765_ net225 _0916_ outputs.div.next_div _0283_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1696_ _0216_ _0213_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2248_ _1208_ _0600_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nand2_1
X_2179_ inputs.frequency_lut.rng\[4\] vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__clkbuf_4
X_2317_ _0492_ _0581_ _0731_ _0745_ _0650_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1481_ outputs.sig_gen.count\[12\] _1073_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__and2_1
X_1550_ _1127_ _1130_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2033_ _0468_ inputs.frequency_lut.rng\[1\] vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__nand2_2
X_2102_ _0537_ _0538_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2866_ clknet_leaf_9_clk _0184_ net47 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1817_ _0328_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__or2_1
X_2797_ clknet_leaf_1_clk _0115_ net28 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_1748_ _0261_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1679_ _0996_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2720_ clknet_leaf_23_clk _0066_ net54 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2651_ clknet_leaf_37_clk inputs.keypad\[12\] net25 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1602_ outputs.output_gen.count\[4\] _1183_ _1170_ outputs.output_gen.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__a22o_1
X_2582_ clknet_leaf_0_clk net68 net25 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1533_ outputs.divider_buffer\[10\] _1107_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nor2_1
X_1464_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[7\] sky130_fd_sc_hd__nor2_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1395_ net303 _0909_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2016_ _0458_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold152 inputs.random_update_clock.count\[1\] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _0937_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold185 inputs.random_update_clock.count\[7\] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 outputs.div.a\[20\] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlygate4sd3_1
X_2849_ clknet_leaf_11_clk _0167_ net42 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold163 outputs.div.a\[11\] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 outputs.div.a\[8\] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 outputs.div.q\[5\] vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2703_ clknet_leaf_7_clk _0049_ net48 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2634_ clknet_leaf_0_clk net63 net25 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2565_ clknet_leaf_26_clk outputs.sample_rate.next_count\[1\] net31 vssd1 vssd1 vccd1
+ vccd1 outputs.sample_rate.count\[1\] sky130_fd_sc_hd__dfrtp_1
X_1516_ _1098_ vssd1 vssd1 vccd1 vccd1 inputs.up.ff_in sky130_fd_sc_hd__clkbuf_1
X_2496_ _0867_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_1447_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__inv_2
X_1378_ outputs.sample_rate.count\[6\] outputs.sample_rate.count\[7\] _0908_ vssd1
+ vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1301_ _0942_ _0943_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2281_ _0637_ _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__or2_1
X_2350_ _0479_ _0591_ _0492_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1996_ outputs.div.m\[4\] net273 _0436_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2617_ clknet_leaf_25_clk inputs.mode_edge.ff_in net30 vssd1 vssd1 vccd1 vccd1 inputs.mode_edge.det_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2548_ _0894_ _0486_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__mux2_1
X_2479_ _0858_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1850_ outputs.div.a\[19\] _0342_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1781_ _0295_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2402_ _0485_ _0586_ _0809_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__a21o_1
X_2333_ _0736_ _0760_ _0554_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2195_ _0598_ _0629_ _0553_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__mux2_1
X_2264_ _0498_ _0653_ _0695_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1979_ _0439_ _0442_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold45 _0145_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 outputs.div.q\[23\] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 inputs.random_update_clock.count\[22\] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 inputs.random_note_generator.out\[2\] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 inputs.random_note_generator.out\[14\] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _0045_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 outputs.signal_buffer2\[8\] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 _0999_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1902_ net195 _0333_ _0377_ net271 _0397_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1833_ _0343_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__nand2_1
X_1764_ _0279_ _0282_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1695_ _0217_ _0219_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2316_ _0579_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2178_ _0489_ _0587_ _0506_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__a21o_1
X_2247_ _0658_ _0671_ _0673_ _0679_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1480_ outputs.sig_gen.count\[12\] _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2032_ _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__clkbuf_4
X_2101_ _0524_ _0515_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__nand2b_2
X_2865_ clknet_leaf_8_clk _0183_ net49 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1816_ _0308_ _0311_ _0320_ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__o31a_2
XFILLER_0_40_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2796_ clknet_leaf_1_clk _0114_ net29 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1747_ outputs.div.a\[9\] _0266_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__xnor2_2
X_1678_ net278 _0916_ _0203_ _0204_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1532_ outputs.divider_buffer\[12\] _1112_ _1113_ outputs.divider_buffer\[11\] vssd1
+ vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1601_ outputs.scaled_buffer\[4\] _1161_ _1182_ _1157_ _1165_ vssd1 vssd1 vccd1 vccd1
+ _1183_ sky130_fd_sc_hd__a221oi_2
X_2581_ clknet_leaf_36_clk net83 net25 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2650_ clknet_leaf_35_clk inputs.keypad\[11\] net22 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1394_ _0994_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__buf_4
X_1463_ outputs.sig_gen.count\[7\] _1058_ _1042_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2015_ outputs.div.m\[13\] net286 _0453_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2848_ clknet_leaf_9_clk _0166_ net46 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold131 outputs.div.q\[18\] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 outputs.div.q\[24\] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 inputs.random_update_clock.count\[6\] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 inputs.random_update_clock.count\[20\] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 outputs.div.a\[24\] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _0035_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 outputs.sig_gen.count\[0\] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__dlygate4sd3_1
X_2779_ clknet_leaf_32_clk _0097_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold120 outputs.div.a\[4\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2702_ clknet_leaf_7_clk net194 net48 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2495_ net289 outputs.sig_gen.count\[12\] _0861_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2564_ clknet_leaf_27_clk outputs.sample_rate.next_count\[0\] net31 vssd1 vssd1 vccd1
+ vccd1 outputs.sample_rate.count\[0\] sky130_fd_sc_hd__dfrtp_1
X_1515_ inputs.up.ff_out inputs.key_encoder.octave_key_up vssd1 vssd1 vccd1 vccd1
+ _1098_ sky130_fd_sc_hd__and2b_1
X_2633_ clknet_leaf_35_clk net73 net22 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1446_ _1010_ _1047_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__nor2_1
X_1377_ net177 _0990_ vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[7\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1300_ inputs.random_update_clock.count\[1\] inputs.random_update_clock.count\[0\]
+ inputs.random_update_clock.count\[3\] inputs.random_update_clock.count\[2\] vssd1
+ vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__or4_1
X_2280_ _0493_ _0634_ _0498_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1995_ _0447_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2616_ clknet_leaf_25_clk net147 net30 vssd1 vssd1 vccd1 vccd1 inputs.mode_edge.ff_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1429_ _1033_ outputs.sig_gen.count\[0\] _1019_ outputs.sig_gen.count\[5\] vssd1
+ vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__a2bb2o_1
X_2478_ net274 outputs.sig_gen.count\[4\] _0850_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__mux2_1
X_2547_ _0951_ _0572_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__nand2_4
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1780_ outputs.div.m\[13\] _0296_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__xnor2_1
X_2401_ _0650_ _0639_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__nand2_1
X_2332_ _1215_ _0754_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2263_ inputs.frequency_lut.rng\[0\] inputs.frequency_lut.rng\[2\] vssd1 vssd1 vccd1
+ vccd1 _0695_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2194_ _0608_ _0628_ _1214_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1978_ outputs.div.q\[1\] outputs.div.q\[0\] _0440_ _0441_ vssd1 vssd1 vccd1 vccd1
+ _0442_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold79 outputs.div.q\[20\] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 _0053_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 inputs.random_update_clock.next_count\[22\] vssd1 vssd1 vccd1 vccd1 net119
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0139_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 outputs.signal_buffer2\[3\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 outputs.output_gen.pwm_ff vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 inputs.keypad_synchronizer.half_sync\[13\] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1832_ outputs.div.a\[17\] _0342_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__or2_1
X_1901_ outputs.div.oscillator_out\[0\] _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1763_ _0281_ _0271_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__nand2_1
X_1694_ outputs.div.m\[5\] _0218_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2246_ _0616_ _0675_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__o21ba_1
X_2315_ _0741_ _0743_ _0507_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2177_ _0485_ _0475_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2100_ _0525_ _0515_ _0522_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__or3b_1
X_2031_ _0468_ inputs.frequency_lut.rng\[1\] vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2864_ clknet_leaf_8_clk _0182_ net47 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1815_ _0306_ _0318_ _0319_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__a21bo_1
X_2795_ clknet_leaf_1_clk _0113_ net28 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1746_ outputs.div.m\[10\] _0265_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__xnor2_2
X_1677_ _0197_ _0202_ _0996_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _0628_ _0662_ _0541_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1531_ outputs.shaper.count\[10\] vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__inv_2
X_1462_ outputs.sig_gen.count\[6\] outputs.sig_gen.count\[7\] _1055_ vssd1 vssd1 vccd1
+ vccd1 _1061_ sky130_fd_sc_hd__and3_1
X_1600_ outputs.scaled_buffer\[3\] _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__xor2_1
X_2580_ clknet_leaf_0_clk net69 net26 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1393_ _0909_ _1000_ vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2014_ _0457_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2847_ clknet_leaf_7_clk _0165_ net48 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold110 outputs.div.a\[16\] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ clknet_leaf_31_clk _0096_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold132 _0048_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 inputs.random_update_clock.count\[15\] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 outputs.div.a\[21\] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _0054_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 outputs.div.q\[10\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 outputs.div.q\[4\] vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 outputs.div.q\[26\] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ outputs.div.m\[8\] _0250_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__xor2_1
Xhold187 outputs.output_gen.count\[5\] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2701_ clknet_leaf_7_clk net144 net45 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2632_ clknet_leaf_30_clk net95 net33 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_2494_ _0866_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__clkbuf_1
X_1445_ _1048_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1514_ _1097_ vssd1 vssd1 vccd1 vccd1 inputs.down.ff_in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2563_ _0905_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
X_1376_ _0992_ vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout60 net61 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1994_ outputs.div.m\[3\] net240 _0436_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2615_ clknet_leaf_16_clk net119 net61 vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2477_ _0857_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
X_1428_ outputs.divider_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2546_ _0892_ _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1359_ inputs.key_encoder.octave_key_up inputs.key_encoder.sync_keys\[15\] vssd1
+ vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2400_ _0822_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2331_ _0759_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
X_2262_ _1208_ _0692_ _0693_ _0464_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__o211a_1
X_2193_ _0565_ _0550_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1977_ outputs.div.q\[3\] outputs.div.q\[2\] outputs.div.q\[5\] outputs.div.q\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2529_ _0884_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold69 outputs.signal_buffer2\[10\] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 outputs.signal_buffer2\[7\] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _0134_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 outputs.div.q\[11\] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 inputs.random_note_generator.out\[0\] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 inputs.keypad_synchronizer.half_sync\[8\] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1831_ outputs.div.a\[17\] _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__nand2_1
X_1900_ _0994_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1762_ _0280_ _0266_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__or2_1
X_1693_ outputs.div.m\[4\] _0209_ _1229_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2245_ _0615_ _0494_ _0677_ _0650_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__a31o_1
X_2176_ _0610_ _0611_ _1207_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__mux2_1
X_2314_ _0477_ _0742_ _0499_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2030_ inputs.frequency_lut.rng\[0\] vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2863_ clknet_leaf_8_clk _0181_ net49 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1814_ _0326_ _0327_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nand2_1
X_2794_ clknet_leaf_11_clk _0112_ net41 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1745_ _0249_ _0264_ _0248_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1676_ _0197_ _0202_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__nand2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _0528_ _0529_ _0546_ _0562_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__a31o_1
X_2228_ _0660_ _0661_ _0534_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1530_ outputs.shaper.count\[11\] vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__inv_2
X_1461_ _1060_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1392_ net223 _0908_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2013_ outputs.div.m\[12\] net256 _0453_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2846_ clknet_leaf_7_clk _0164_ net48 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold144 inputs.random_update_clock.count\[16\] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _0040_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 outputs.div.q\[8\] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 outputs.div.q_out\[5\] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 outputs.div.a\[0\] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _0248_ _0249_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__nand2_1
X_2777_ clknet_leaf_1_clk _0095_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold166 outputs.div.a\[15\] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _0055_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold177 outputs.div.divisor\[15\] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ net210 _0916_ outputs.div.next_div _1235_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a22o_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 _0989_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 outputs.output_gen.count\[3\] vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2700_ clknet_leaf_6_clk net138 net44 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2631_ clknet_leaf_36_clk net71 net25 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2562_ _0904_ _0658_ _0895_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__mux2_1
X_2493_ net275 outputs.sig_gen.count\[11\] _0861_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1444_ _1041_ _1046_ _1047_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__and3_1
X_1375_ _0990_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1513_ inputs.down.ff_out inputs.down.in vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2829_ clknet_leaf_13_clk net127 net49 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout50 net19 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_4
Xfanout61 net62 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _0446_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2614_ clknet_leaf_16_clk inputs.random_update_clock.next_count\[21\] net61 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2545_ _0492_ _1093_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2476_ net267 outputs.sig_gen.count\[3\] _0850_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__mux2_1
X_1427_ outputs.divider_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__inv_2
X_1358_ net146 net92 inputs.key_encoder.sync_keys\[14\] vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.mode_key
+ sky130_fd_sc_hd__nor3b_1
X_1289_ net214 net169 vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ net295 _0758_ _0606_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__mux2_1
X_2261_ _1208_ _0610_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__nand2_1
X_2192_ inputs.key_encoder.sync_keys\[12\] _1199_ _0526_ _0523_ _0516_ vssd1 vssd1
+ vccd1 vccd1 _0627_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1976_ outputs.div.q\[7\] outputs.div.q\[6\] outputs.div.q\[8\] vssd1 vssd1 vccd1
+ vccd1 _0440_ sky130_fd_sc_hd__or3b_1
XFILLER_0_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2528_ outputs.shaper.count\[10\] net131 _0396_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold59 _0138_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ net120 _0829_ _0407_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__a21o_1
Xhold37 _0041_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 outputs.signal_buffer2\[2\] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 inputs.random_note_generator.out\[11\] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 inputs.random_note_generator.out\[12\] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1830_ outputs.div.m\[17\] _0336_ _0248_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__o21a_2
X_1761_ outputs.div.a\[9\] vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__inv_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1692_ outputs.div.a\[4\] vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
X_2313_ _0468_ _0466_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2175_ _0542_ _0564_ _0556_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__mux2_1
X_2244_ _0577_ _0676_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__nand2_1
X_1959_ outputs.scaled_buffer\[1\] net154 _1001_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2862_ clknet_leaf_8_clk _0180_ net48 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1813_ _0323_ _0325_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__nand2_1
X_2793_ clknet_leaf_31_clk _0111_ net37 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1744_ outputs.div.m\[9\] outputs.div.m\[8\] vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ _0200_ _0201_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__nor2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2158_ _0578_ _0584_ _0590_ _0594_ _0506_ _0508_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__mux4_1
X_2227_ _0515_ _0527_ _0546_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__o21a_1
X_2089_ _0526_ _0522_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1460_ _1041_ _1057_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__and3_1
X_1391_ _0908_ net140 vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2012_ _0456_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__clkbuf_1
X_2845_ clknet_leaf_7_clk _0163_ net48 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold123 inputs.random_update_clock.count\[14\] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 outputs.div.q\[14\] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 inputs.random_update_clock.count\[19\] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 outputs.sig_gen.count\[17\] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold167 outputs.div.a\[17\] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 outputs.div.q_out\[4\] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ clknet_leaf_11_clk _0094_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[17\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold101 _0074_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _1226_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__xor2_1
X_1727_ outputs.div.m\[7\] outputs.div.m\[6\] _0209_ _0224_ vssd1 vssd1 vccd1 vccd1
+ _0249_ sky130_fd_sc_hd__or4_2
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold189 outputs.div.a\[19\] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ outputs.scaled_buffer\[0\] net21 outputs.scaled_buffer\[1\] vssd1 vssd1 vccd1
+ vccd1 _1171_ sky130_fd_sc_hd__a21oi_1
Xhold178 outputs.div.divisor\[3\] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2492_ _0865_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2630_ clknet_leaf_29_clk net76 net32 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1512_ _1096_ vssd1 vssd1 vccd1 vccd1 inputs.mode_edge.ff_in sky130_fd_sc_hd__inv_2
X_2561_ _0699_ _1093_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__xor2_1
X_1443_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] outputs.sig_gen.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__nand3_1
X_1374_ outputs.output_gen.count\[6\] _0988_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2828_ clknet_leaf_8_clk net136 net49 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2759_ clknet_leaf_1_clk _0077_ net28 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout62 net19 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_2
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout51 net62 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_4
Xfanout40 net43 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ outputs.div.m\[2\] net222 _0436_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2613_ clknet_leaf_16_clk inputs.random_update_clock.next_count\[20\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[20\] sky130_fd_sc_hd__dfrtp_1
X_2475_ _0856_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2544_ _0658_ _0699_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1288_ net169 vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[0\]
+ sky130_fd_sc_hd__inv_2
X_1357_ net118 _0981_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[22\]
+ sky130_fd_sc_hd__xnor2_1
X_1426_ outputs.divider_buffer\[13\] _1004_ _1022_ outputs.sig_gen.count\[14\] _1031_
+ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2191_ _0626_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_1
X_2260_ _0556_ _0690_ _0691_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1975_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold16 inputs.keypad_synchronizer.half_sync\[4\] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dlygate4sd3_1
X_2527_ _0883_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
X_2458_ net101 _0829_ _0406_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1409_ _1014_ outputs.sig_gen.count\[10\] _1003_ outputs.sig_gen.count\[1\] vssd1
+ vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__a2bb2o_1
Xhold27 inputs.keypad_synchronizer.half_sync\[16\] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 outputs.output_gen.count\[0\] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_1
Xhold49 outputs.signal_buffer2\[17\] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _0616_ _0499_ _0467_ _0476_ _0507_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__a41o_1
XFILLER_0_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1760_ _0276_ _0278_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1691_ _0215_ _0211_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__or2_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ _0498_ _0479_ _0591_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__or3_1
X_2243_ inputs.frequency_lut.rng\[3\] _0585_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__or2_1
X_2174_ _0552_ _0609_ _0554_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1958_ _0429_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
X_1889_ _0377_ _0392_ _0393_ _0333_ net302 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2861_ clknet_leaf_7_clk _0179_ net48 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1812_ _0323_ _0325_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__or2_1
X_1743_ net268 _0916_ _0262_ _0263_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a22o_1
X_2792_ clknet_leaf_31_clk _0110_ net37 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1674_ outputs.div.a\[2\] _0199_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _0521_ _0527_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__nor2_1
X_2157_ _0495_ _0592_ _0593_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2088_ _0525_ _1202_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1390_ outputs.sample_rate.count\[4\] _0907_ net139 vssd1 vssd1 vccd1 vccd1 _0999_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2011_ outputs.div.m\[11\] net288 _0453_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__mux2_1
X_2844_ clknet_leaf_6_clk _0162_ net50 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold124 _0971_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _0044_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 outputs.div.q\[12\] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 outputs.div.q_out\[0\] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlygate4sd3_1
X_2775_ clknet_leaf_11_clk _0093_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold113 _0073_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 outputs.div.q_out\[7\] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 outputs.div.divisor\[14\] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__or2_1
X_1588_ outputs.scaled_buffer\[3\] _1161_ _1169_ _1157_ _1165_ vssd1 vssd1 vccd1 vccd1
+ _1170_ sky130_fd_sc_hd__a221oi_2
X_1726_ _1229_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__buf_2
Xhold179 outputs.output_gen.count\[2\] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _0572_ _0633_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2491_ net276 outputs.sig_gen.count\[10\] _0861_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1442_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] outputs.sig_gen.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__a21o_1
X_2560_ _0895_ _0893_ _0903_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__o21ai_1
X_1511_ net149 inputs.key_encoder.mode_key vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1373_ outputs.output_gen.count\[6\] _0988_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2827_ clknet_leaf_8_clk net107 net49 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2758_ clknet_leaf_5_clk outputs.sig_gen.next_count\[17\] net44 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2689_ clknet_leaf_19_clk net259 net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1709_ _0217_ _0219_ _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__a21o_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout52 net62 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_2
XFILLER_0_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout41 net42 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_4
Xfanout30 net31 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2612_ clknet_leaf_18_clk inputs.random_update_clock.next_count\[19\] net55 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1991_ _0445_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2543_ _0891_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
X_1425_ _1030_ outputs.sig_gen.count\[6\] outputs.divider_buffer\[16\] _1023_ vssd1
+ vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__o22a_1
X_2474_ net279 outputs.sig_gen.count\[2\] _0850_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__mux2_1
X_1356_ _0982_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[21\]
+ sky130_fd_sc_hd__clkbuf_1
X_1287_ _0935_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2190_ net222 _0625_ _0606_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1974_ outputs.div.div _0910_ _0913_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2526_ outputs.shaper.count\[9\] net116 _0396_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__mux2_1
X_2457_ net123 _0829_ _0404_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__a21o_1
Xhold39 outputs.signal_buffer2\[6\] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ outputs.divider_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__inv_2
Xhold28 inputs.keypad_synchronizer.half_sync\[6\] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 inputs.random_note_generator.out\[3\] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _0696_ _0810_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1339_ inputs.random_update_clock.count\[15\] _0970_ vssd1 vssd1 vccd1 vccd1 _0972_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1690_ outputs.div.a\[3\] vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _0740_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
X_2242_ _0495_ _0674_ _0485_ _0591_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_20_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2173_ _0597_ _0608_ _1214_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ outputs.scaled_buffer\[0\] net164 _1001_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__mux2_1
X_1888_ _0383_ _0387_ _0391_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__nand3_1
X_2509_ _0874_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_36_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2860_ clknet_leaf_6_clk _0178_ net50 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1811_ outputs.div.m\[16\] _0324_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__xnor2_1
X_2791_ clknet_leaf_1_clk _0109_ net28 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1742_ _0252_ _0255_ _0261_ _0996_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__o31a_1
X_1673_ outputs.div.a\[2\] _0199_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2225_ _0506_ _0654_ _0655_ _0657_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__o311a_1
XFILLER_0_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2156_ _0494_ _0497_ _0485_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2087_ _1199_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2010_ _0455_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__clkbuf_1
X_2843_ clknet_leaf_6_clk _0161_ net50 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2774_ clknet_leaf_11_clk _0092_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_1725_ outputs.div.a\[7\] vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold125 outputs.div.q\[19\] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold114 outputs.div.count\[2\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _0042_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _0069_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 outputs.div.q_out\[6\] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _0076_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ outputs.scaled_buffer\[2\] _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__xnor2_1
X_1656_ _1230_ _1231_ outputs.div.a\[0\] vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__a21oi_1
Xhold169 outputs.div.a\[2\] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _0484_ _0488_ _0470_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__o21ai_1
X_2208_ _0603_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2490_ _0864_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1441_ _1045_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_1510_ _1094_ _1095_ vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.feedback
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1372_ _0988_ net250 vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2826_ clknet_leaf_8_clk net115 net48 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2757_ clknet_leaf_5_clk outputs.sig_gen.next_count\[16\] net44 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[16\] sky130_fd_sc_hd__dfrtp_1
X_2688_ clknet_leaf_19_clk _0034_ net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1708_ _0215_ _0211_ _0219_ _0217_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__o22a_1
X_1639_ inputs.octave_fsm.state\[1\] inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__a21o_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout42 net43 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_4
Xfanout53 net56 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_4
Xfanout31 net32 vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1990_ outputs.div.m\[1\] net280 _0436_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__mux2_1
X_2542_ net305 net111 _0396_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__mux2_1
X_2611_ clknet_leaf_17_clk inputs.random_update_clock.next_count\[18\] net55 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[18\] sky130_fd_sc_hd__dfrtp_1
X_1355_ _0955_ _0980_ _0981_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__and3_1
X_2473_ _0855_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
X_1424_ outputs.divider_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__inv_2
X_1286_ net1 outputs.pwm_output vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2809_ clknet_leaf_2_clk _0127_ net41 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1973_ _0437_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2525_ _0882_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1338_ _0970_ net186 vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
X_1407_ outputs.divider_buffer\[3\] _1010_ outputs.divider_buffer\[9\] _1011_ _1012_
+ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__a221o_1
X_2456_ net105 _0829_ _0403_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold18 inputs.random_note_generator.out\[9\] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 inputs.random_note_generator.out\[13\] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ _0482_ _0467_ _0803_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1269_ _0926_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ net292 _0739_ _0606_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__mux2_1
X_2241_ _0481_ _0477_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__nor2_1
X_2172_ _0531_ _0528_ _0539_ _0547_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1956_ _0428_ _0425_ _1001_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__a21oi_1
X_1887_ _0383_ _0387_ _0391_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2508_ outputs.shaper.count\[0\] net128 _0872_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__mux2_1
X_2439_ outputs.divider_buffer\[12\] outputs.div.m\[12\] _0839_ vssd1 vssd1 vccd1
+ vccd1 _0847_ sky130_fd_sc_hd__mux2_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810_ outputs.div.m\[15\] _0314_ _0248_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__o21a_1
X_1741_ _0252_ _0255_ _0261_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__o21ai_1
X_2790_ clknet_leaf_1_clk _0108_ net28 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1672_ outputs.div.m\[3\] _0198_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _0481_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__nor2_1
X_2224_ _0650_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2086_ _0517_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__or2_1
X_1939_ outputs.div.oscillator_out\[17\] _0411_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2842_ clknet_leaf_6_clk _0160_ net50 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold126 outputs.div.a\[23\] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold104 outputs.div.a\[14\] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dlygate4sd3_1
X_2773_ clknet_leaf_11_clk _0091_ net41 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[14\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold115 outputs.output_gen.count\[7\] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ _0229_ _0234_ _0242_ _0245_ _0241_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__o32a_2
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold159 inputs.random_update_clock.count\[11\] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _0075_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] net21 vssd1 vssd1 vccd1
+ vccd1 _1168_ sky130_fd_sc_hd__o21ai_1
Xhold148 outputs.div.a\[1\] vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ outputs.div.a\[0\] _1230_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__and3_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ _0575_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2207_ _0635_ _0638_ _0640_ _0641_ _0615_ _0507_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__mux4_1
X_2069_ inputs.frequency_lut.rng\[5\] vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1440_ _1042_ _1043_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__and3_1
X_1371_ outputs.output_gen.count\[4\] _0986_ net249 vssd1 vssd1 vccd1 vccd1 _0989_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2825_ clknet_leaf_7_clk net104 net48 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2756_ clknet_leaf_5_clk outputs.sig_gen.next_count\[15\] net44 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[15\] sky130_fd_sc_hd__dfrtp_2
X_2687_ clknet_leaf_19_clk net253 net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1707_ _0216_ _0230_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1638_ _1213_ _1218_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1569_ _1007_ outputs.shaper.count\[16\] outputs.shaper.count\[0\] _1003_ vssd1 vssd1
+ vccd1 vccd1 _1151_ sky130_fd_sc_hd__o22a_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout43 net19 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout54 net56 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout32 net38 vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2541_ _0890_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
X_2610_ clknet_leaf_17_clk inputs.random_update_clock.next_count\[17\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[17\] sky130_fd_sc_hd__dfrtp_1
X_2472_ net281 outputs.sig_gen.count\[1\] _0850_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1354_ inputs.random_update_clock.count\[21\] _0978_ vssd1 vssd1 vccd1 vccd1 _0981_
+ sky130_fd_sc_hd__nand2_1
X_1285_ _0934_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[16\] sky130_fd_sc_hd__clkbuf_1
X_1423_ outputs.divider_buffer\[7\] _1026_ outputs.divider_buffer\[11\] _1027_ _1028_
+ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2808_ clknet_leaf_2_clk _0126_ net41 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2739_ clknet_leaf_22_clk outputs.output_gen.next_count\[6\] net34 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1972_ net308 net219 _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2524_ net301 net129 _0872_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__mux2_1
X_2455_ net108 _0829_ _0402_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1337_ inputs.random_update_clock.count\[13\] _0964_ net185 vssd1 vssd1 vccd1 vccd1
+ _0971_ sky130_fd_sc_hd__a21oi_1
X_1406_ outputs.divider_buffer\[4\] outputs.sig_gen.count\[4\] vssd1 vssd1 vccd1 vccd1
+ _1012_ sky130_fd_sc_hd__xor2_1
Xhold19 inputs.random_note_generator.out\[1\] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dlygate4sd3_1
X_1268_ _0917_ net17 vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__and2b_1
X_2386_ _0482_ _0586_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2171_ _0607_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
X_2240_ _0499_ _0496_ _0672_ _0616_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1955_ net235 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
X_1886_ _0389_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2507_ _0873_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2438_ _0846_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2369_ _1206_ _0754_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__or2_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1671_ outputs.div.m\[2\] _1229_ _1238_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__a21o_1
X_1740_ _0259_ _0260_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0486_ _0465_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__nor2_2
X_2223_ _0497_ _0587_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__a21bo_1
X_2085_ _0521_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1938_ outputs.div.q\[24\] _0915_ _0996_ net96 _0417_ vssd1 vssd1 vccd1 vccd1 _0053_
+ sky130_fd_sc_hd__a221o_1
X_1869_ _0205_ _0375_ _0376_ _0333_ net243 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2841_ clknet_leaf_6_clk _0159_ net45 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold116 outputs.div.q\[21\] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 inputs.random_update_clock.count\[4\] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 outputs.div.q\[13\] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 outputs.div.q\[9\] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ outputs.div.m\[0\] outputs.div.m\[1\] _1229_ vssd1 vssd1 vccd1 vccd1 _1231_
+ sky130_fd_sc_hd__nand3_1
X_2772_ clknet_leaf_1_clk _0090_ net28 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[13\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold149 outputs.div.a\[7\] vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dlygate4sd3_1
X_1723_ _0237_ _0239_ _0227_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _1156_ _1159_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__o21a_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2206_ _0503_ _0577_ _0582_ _0491_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2137_ net283 _0574_ _0453_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__mux2_1
X_2068_ _0505_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1370_ outputs.output_gen.count\[5\] outputs.output_gen.count\[4\] _0986_ vssd1 vssd1
+ vccd1 vccd1 _0988_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2824_ clknet_leaf_6_clk net113 net45 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2755_ clknet_leaf_5_clk outputs.sig_gen.next_count\[14\] net44 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2686_ clknet_leaf_19_clk net234 net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1706_ _0215_ _0211_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__nand2_1
X_1637_ inputs.octave_fsm.state\[1\] _1212_ _1215_ _1217_ vssd1 vssd1 vccd1 vccd1
+ _1218_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1499_ _1023_ _1085_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__nor2_1
X_1568_ _1140_ _1136_ _1126_ _1149_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__or4b_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout44 net45 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_4
Xfanout55 net56 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout33 net37 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout22 net23 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2540_ outputs.shaper.count\[16\] net126 _0396_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__mux2_1
X_1422_ outputs.divider_buffer\[8\] outputs.sig_gen.count\[8\] vssd1 vssd1 vccd1 vccd1
+ _1028_ sky130_fd_sc_hd__xor2_1
X_2471_ _0854_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1353_ inputs.random_update_clock.count\[21\] _0978_ vssd1 vssd1 vccd1 vccd1 _0980_
+ sky130_fd_sc_hd__or2_1
X_1284_ net1 net8 vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2807_ clknet_leaf_3_clk _0125_ net39 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2738_ clknet_leaf_24_clk outputs.output_gen.next_count\[5\] net35 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2669_ clknet_leaf_20_clk _0015_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1971_ _0411_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2523_ _0881_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
X_1405_ outputs.sig_gen.count\[9\] vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__inv_2
X_2454_ net110 _0829_ _0401_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2385_ _0481_ _0486_ _0473_ _0466_ _0615_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a41o_1
X_1267_ _0925_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[7\] sky130_fd_sc_hd__clkbuf_1
Xinput1 cs vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_8
X_1336_ inputs.random_update_clock.count\[13\] inputs.random_update_clock.count\[14\]
+ _0964_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2170_ net280 _0605_ _0606_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1954_ _0427_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1885_ outputs.div.a\[24\] _0355_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2506_ net290 outputs.sig_gen.count\[17\] _0872_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2437_ outputs.divider_buffer\[11\] outputs.div.m\[11\] _0839_ vssd1 vssd1 vccd1
+ vccd1 _0846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2368_ _0699_ _0727_ _0792_ _0793_ _0508_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1319_ _0951_ _0957_ _0958_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2299_ _0482_ _0477_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a21o_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1670_ _0192_ _0196_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _0491_ _0588_ _0615_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__a21oi_1
X_2153_ _0579_ _0585_ _0587_ _0589_ _0468_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__o32a_1
X_2084_ inputs.key_encoder.sync_keys\[12\] _0516_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1937_ outputs.div.oscillator_out\[16\] _0411_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1868_ _0360_ _0365_ _0374_ _0371_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__nand4_1
X_1799_ outputs.div.m\[14\] outputs.div.m\[13\] outputs.div.m\[12\] _0285_ vssd1 vssd1
+ vccd1 vccd1 _0314_ sky130_fd_sc_hd__or4_2
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2840_ clknet_leaf_5_clk _0158_ net44 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2771_ clknet_leaf_1_clk _0089_ net28 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold139 outputs.div.q\[22\] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _0051_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 _0043_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1653_ outputs.div.m\[0\] _1229_ outputs.div.m\[1\] vssd1 vssd1 vccd1 vccd1 _1230_
+ sky130_fd_sc_hd__a21o_1
X_1584_ outputs.scaled_buffer\[5\] _1161_ _1165_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__a21oi_1
X_1722_ net211 _0916_ outputs.div.next_div _0244_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold128 outputs.div.a\[6\] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2205_ _0579_ _0585_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2136_ _0464_ _0509_ _0573_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__o21ai_1
X_2067_ inputs.frequency_lut.rng\[4\] vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2823_ clknet_leaf_6_clk net132 net45 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2754_ clknet_leaf_5_clk outputs.sig_gen.next_count\[13\] net44 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1705_ _0227_ _0228_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1567_ _1007_ outputs.shaper.count\[16\] outputs.shaper.count\[17\] vssd1 vssd1 vccd1
+ vccd1 _1149_ sky130_fd_sc_hd__a21oi_1
X_2685_ clknet_leaf_17_clk _0031_ net55 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1636_ inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\] _1216_ _1208_ _1210_
+ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__o32a_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1023_ _1085_ _1087_ _1042_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[16\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ _0530_ _0521_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__or2b_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout45 net50 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout56 net62 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_2
Xfanout34 net36 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout23 net38 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_2
XFILLER_0_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1421_ outputs.sig_gen.count\[11\] vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2470_ net265 outputs.sig_gen.count\[0\] _0850_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1283_ _0933_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[15\] sky130_fd_sc_hd__clkbuf_1
X_1352_ _0978_ _0979_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[20\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2668_ clknet_leaf_19_clk _0014_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2806_ clknet_leaf_37_clk _0124_ net26 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_2737_ clknet_leaf_24_clk outputs.output_gen.next_count\[4\] net35 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2599_ clknet_leaf_17_clk inputs.random_update_clock.next_count\[6\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[6\] sky130_fd_sc_hd__dfrtp_1
X_1619_ inputs.key_encoder.sync_keys\[13\] inputs.key_encoder.sync_keys\[1\] inputs.key_encoder.sync_keys\[0\]
+ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1970_ _0435_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__clkbuf_1
X_2522_ net304 net120 _0872_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1335_ _0969_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[13\]
+ sky130_fd_sc_hd__clkbuf_1
X_1404_ outputs.sig_gen.count\[3\] vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__inv_2
X_2453_ net125 _0829_ _0399_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__a21o_1
X_2384_ _0808_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_1
Xinput2 gpio[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_1266_ _0917_ net16 vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1953_ _0910_ _0425_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__and3_1
X_1884_ outputs.div.a\[24\] _0355_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2505_ _0994_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1318_ inputs.random_update_clock.count\[8\] _0954_ vssd1 vssd1 vccd1 vccd1 _0958_
+ sky130_fd_sc_hd__and2_1
X_2436_ _0845_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2298_ _0589_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__nand2_1
X_2367_ _0482_ _0586_ _0585_ _0697_ _0505_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__o311a_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ _0915_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__clkbuf_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ _0484_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__nand2_1
X_2221_ _0502_ _0647_ _0484_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2083_ _0518_ _0520_ inputs.key_encoder.sync_keys\[11\] inputs.key_encoder.sync_keys\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__a211o_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1936_ net96 _0915_ _0405_ net201 _0416_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a221o_1
X_1867_ _0360_ _0365_ _0371_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1798_ _0205_ _0312_ _0313_ _1228_ net166 vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2419_ _0836_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2770_ clknet_leaf_0_clk _0088_ net26 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1721_ _0242_ _0243_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 inputs.random_update_clock.count\[0\] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_1
Xhold118 outputs.div.a\[10\] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ outputs.div.a\[25\] vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__inv_2
X_1583_ net21 _1162_ _1164_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__o21ai_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold129 outputs.div.a\[5\] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _0468_ _0637_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__and2_1
X_2135_ _1224_ _0555_ _0571_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2066_ _0492_ _0477_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__a21oi_1
X_1919_ net150 _0400_ _0405_ net196 _0407_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2822_ clknet_leaf_6_clk net117 net45 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2753_ clknet_leaf_4_clk outputs.sig_gen.next_count\[12\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[12\] sky130_fd_sc_hd__dfrtp_2
X_2684_ clknet_leaf_17_clk _0030_ net55 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1704_ _0223_ _0226_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1497_ _1023_ _1085_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__nand2_1
X_1566_ _1100_ _1106_ _1146_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__o31ai_2
X_1635_ inputs.octave_fsm.state\[1\] _1210_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__nor2_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2118_ inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__a21oi_4
X_2049_ _0486_ _0473_ _0466_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__a21o_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout57 net62 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_4
Xfanout46 net50 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout35 net36 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
Xfanout24 net25 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1351_ net218 _0977_ net226 vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__a21oi_1
X_1420_ outputs.sig_gen.count\[7\] vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1282_ net1 net7 vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2805_ clknet_leaf_3_clk _0123_ net39 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2667_ clknet_leaf_21_clk _0013_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2736_ clknet_leaf_24_clk outputs.output_gen.next_count\[3\] net35 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1618_ inputs.key_encoder.sync_keys\[2\] inputs.key_encoder.sync_keys\[3\] vssd1
+ vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2598_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[5\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_1549_ outputs.divider_buffer\[3\] _1125_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2521_ _0880_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1265_ _0924_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[6\] sky130_fd_sc_hd__clkbuf_1
X_1334_ _0955_ _0967_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__and3_1
X_1403_ _1006_ outputs.sig_gen.count\[9\] _1007_ outputs.sig_gen.count\[17\] _1008_
+ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__a221o_1
X_2452_ net128 _0829_ _0397_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__a21o_1
X_2383_ net286 _0807_ _0798_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__mux2_1
Xinput3 gpio[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2719_ clknet_leaf_19_clk _0065_ net54 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1952_ outputs.div.start _0422_ outputs.div.count\[3\] vssd1 vssd1 vccd1 vccd1 _0426_
+ sky130_fd_sc_hd__a21o_1
X_1883_ _0386_ _0388_ net215 _0916_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2504_ _0871_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
X_2435_ outputs.divider_buffer\[10\] outputs.div.m\[10\] _0839_ vssd1 vssd1 vccd1
+ vccd1 _0845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1317_ inputs.random_update_clock.count\[8\] _0954_ vssd1 vssd1 vccd1 vccd1 _0957_
+ sky130_fd_sc_hd__nor2_1
X_1248_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2297_ _0481_ _0466_ _0470_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__nand3_1
X_2366_ _0485_ _0586_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2082_ _1200_ _0519_ inputs.key_encoder.sync_keys\[6\] inputs.key_encoder.sync_keys\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__a211o_1
X_2151_ _0465_ _0473_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__and2b_1
X_2220_ _0479_ _0653_ _0499_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__o21a_1
X_1935_ net313 _0411_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__and2_1
X_1866_ _0372_ _0373_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1797_ _0308_ _0311_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2418_ outputs.divider_buffer\[2\] outputs.div.m\[2\] _0798_ vssd1 vssd1 vccd1 vccd1
+ _0836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2349_ _0499_ _0480_ _0775_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 outputs.div.q_out\[3\] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ _1225_ _1226_ _1227_ _1228_ net173 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a32o_1
X_1720_ _0229_ _0234_ _0227_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold119 outputs.div.a\[12\] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ outputs.scaled_buffer\[6\] _1158_ _1163_ outputs.scaled_buffer\[7\] vssd1
+ vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or4b_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _0580_ _0592_ _0636_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__a31oi_1
X_2065_ _0486_ _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__nor2_1
X_2134_ _0533_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1918_ outputs.div.oscillator_out\[7\] _0398_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__and2_1
X_1849_ _0330_ _0354_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ clknet_leaf_7_clk net130 net44 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2683_ clknet_leaf_17_clk _0029_ net55 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2752_ clknet_leaf_4_clk outputs.sig_gen.next_count\[11\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[11\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1703_ _0223_ _0226_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__or2_1
X_1634_ _1214_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__inv_2
X_1496_ _1086_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
X_1565_ _1104_ _1105_ _1007_ outputs.shaper.count\[16\] vssd1 vssd1 vccd1 vccd1 _1147_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2048_ inputs.frequency_lut.rng\[0\] vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__clkbuf_4
X_2117_ _0542_ _0552_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__mux2_1
Xfanout58 net62 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_2
Xfanout47 net50 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout36 net37 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_2
Xfanout25 net26 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1350_ inputs.random_update_clock.count\[19\] inputs.random_update_clock.count\[20\]
+ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1281_ _0932_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[14\] sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2804_ clknet_leaf_0_clk _0122_ net26 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2597_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[4\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[4\] sky130_fd_sc_hd__dfrtp_1
X_2666_ clknet_leaf_21_clk _0012_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_2735_ clknet_leaf_24_clk outputs.output_gen.next_count\[2\] net35 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_1617_ inputs.key_encoder.sync_keys\[11\] inputs.key_encoder.sync_keys\[8\] inputs.key_encoder.sync_keys\[9\]
+ inputs.key_encoder.sync_keys\[10\] vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__or4_4
X_1479_ _1027_ _1070_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__nor2_1
X_1548_ outputs.divider_buffer\[1\] _1128_ _1127_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2520_ outputs.shaper.count\[6\] net101 _0872_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__mux2_1
X_1402_ outputs.divider_buffer\[12\] outputs.sig_gen.count\[12\] vssd1 vssd1 vccd1
+ vccd1 _1008_ sky130_fd_sc_hd__xor2_1
X_2451_ _0853_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1264_ _0917_ net15 vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__and2b_1
X_1333_ inputs.random_update_clock.count\[13\] _0964_ vssd1 vssd1 vccd1 vccd1 _0968_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2382_ _0572_ _0800_ _0806_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__o21ai_1
Xinput4 gpio[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2718_ clknet_leaf_18_clk _0064_ net54 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2649_ clknet_leaf_13_clk inputs.keypad\[10\] net58 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1951_ _0424_ _0913_ _0423_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__or3_1
X_1882_ _0996_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2503_ net291 outputs.sig_gen.count\[16\] _0861_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2434_ _0844_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2365_ _0699_ _0788_ _0790_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__a21o_1
X_1316_ _0954_ _0956_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[7\]
+ sky130_fd_sc_hd__nor2_1
X_1247_ _0910_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2296_ _0482_ _0489_ _0494_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2081_ inputs.key_encoder.sync_keys\[4\] inputs.key_encoder.sync_keys\[5\] vssd1
+ vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__nor2_1
X_2150_ _0481_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1934_ outputs.div.q\[22\] _0915_ _0405_ net178 _0415_ vssd1 vssd1 vccd1 vccd1 _0051_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1865_ outputs.div.a\[21\] _0355_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__or2_1
X_1796_ _0308_ _0311_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2417_ _0835_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__clkbuf_1
X_2348_ _0484_ _0579_ _0585_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2279_ _0482_ _0695_ _0709_ _0581_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1650_ _0915_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__clkbuf_4
Xhold109 _0072_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dlygate4sd3_1
X_1581_ outputs.scaled_buffer\[5\] outputs.scaled_buffer\[4\] _1099_ vssd1 vssd1 vccd1
+ vccd1 _1163_ sky130_fd_sc_hd__or3_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2202_ _0484_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2064_ _0473_ _0466_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nor2_2
X_2133_ _0556_ _0564_ _0570_ _1207_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__o211a_1
X_1917_ outputs.div.q\[14\] _0400_ _0405_ net167 _0406_ vssd1 vssd1 vccd1 vccd1 _0043_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1848_ outputs.div.a\[18\] _0355_ _0348_ _0356_ _0357_ vssd1 vssd1 vccd1 vccd1 _0358_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1779_ outputs.div.m\[12\] _0285_ _0248_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2820_ clknet_leaf_9_clk net121 net46 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2751_ clknet_leaf_4_clk outputs.sig_gen.next_count\[10\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1564_ _1117_ _1118_ _1144_ _1145_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__o31a_1
X_2682_ clknet_leaf_12_clk _0028_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1702_ outputs.div.m\[6\] _0225_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__xnor2_1
X_1633_ inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _1214_ sky130_fd_sc_hd__nor2b_2
X_1495_ _1041_ _1084_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout37 net38 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_2
Xfanout26 net38 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_4
X_2047_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__clkbuf_4
X_2116_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__clkbuf_4
Xfanout48 net50 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_4
Xfanout59 net61 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1280_ net1 net6 vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2803_ clknet_leaf_1_clk _0121_ net29 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2734_ clknet_leaf_24_clk outputs.output_gen.next_count\[1\] net34 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2596_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[3\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1547_ outputs.divider_buffer\[2\] outputs.shaper.count\[1\] vssd1 vssd1 vccd1 vccd1
+ _1129_ sky130_fd_sc_hd__or2b_1
X_2665_ clknet_leaf_31_clk _0011_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1616_ inputs.key_encoder.sync_keys\[14\] inputs.key_encoder.sync_keys\[15\] inputs.key_encoder.octave_key_up
+ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__nor3_2
X_1478_ _1027_ _1070_ _1072_ _1042_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[11\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2450_ net312 outputs.div.m\[17\] _0850_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__mux2_1
X_1401_ outputs.divider_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
X_2381_ _0658_ _0801_ _0805_ _0603_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__a211o_1
X_1332_ inputs.random_update_clock.count\[13\] _0964_ vssd1 vssd1 vccd1 vccd1 _0967_
+ sky130_fd_sc_hd__or2_1
X_1263_ _0923_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 gpio[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2717_ clknet_leaf_18_clk _0063_ net54 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2648_ clknet_leaf_3_clk inputs.keypad\[9\] net39 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2579_ clknet_leaf_36_clk net84 net26 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1950_ outputs.div.count\[3\] vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
X_2502_ _0870_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
X_1881_ _0381_ _0382_ _0385_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1315_ net247 _0952_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__o21ai_1
X_2433_ outputs.divider_buffer\[9\] outputs.div.m\[9\] _0839_ vssd1 vssd1 vccd1 vccd1
+ _0844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2364_ _0506_ _0499_ _0730_ _0789_ _0650_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1246_ outputs.div.count\[3\] outputs.div.count\[4\] _0911_ _0912_ vssd1 vssd1 vccd1
+ vccd1 _0913_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2295_ _0498_ _0479_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ inputs.key_encoder.sync_keys\[8\] inputs.key_encoder.sync_keys\[9\] vssd1
+ vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__nor2_1
X_1933_ outputs.div.oscillator_out\[14\] _0411_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1864_ outputs.div.a\[21\] _0355_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__nand2_1
X_1795_ _0290_ _0292_ _0300_ _0310_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2416_ outputs.divider_buffer\[1\] outputs.div.m\[1\] _0798_ vssd1 vssd1 vccd1 vccd1
+ _0835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2278_ _0491_ _0470_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__nand2_1
X_2347_ _0587_ _0742_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1580_ inputs.wavetype_fsm.state\[0\] inputs.wavetype_fsm.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _1162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ inputs.frequency_lut.rng\[1\] inputs.frequency_lut.rng\[2\] vssd1 vssd1 vccd1
+ vccd1 _0636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2132_ _0541_ _0568_ _0569_ _0554_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2063_ _0492_ _0496_ _0500_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1916_ outputs.div.oscillator_out\[6\] _0398_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1847_ _0343_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1778_ outputs.div.a\[12\] vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2681_ clknet_leaf_12_clk _0027_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2750_ clknet_leaf_4_clk outputs.sig_gen.next_count\[9\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1701_ _0209_ _0224_ _1229_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1494_ outputs.sig_gen.count\[15\] _1083_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nand2_1
X_1563_ _1111_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__inv_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1632_ _1208_ _1209_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__a21oi_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a21o_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout49 net50 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_2
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout38 net19 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_2
Xfanout27 net29 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_4
X_2046_ inputs.frequency_lut.rng\[3\] vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2802_ clknet_leaf_0_clk _0120_ net26 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2664_ clknet_leaf_21_clk _0010_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2733_ clknet_leaf_25_clk outputs.output_gen.next_count\[0\] net34 vssd1 vssd1 vccd1
+ vccd1 outputs.output_gen.count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2595_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[2\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_1477_ _1027_ _1070_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nand2_1
X_1546_ outputs.shaper.count\[0\] vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1615_ outputs.output_gen.count\[7\] _1194_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2029_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1331_ _0966_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[12\]
+ sky130_fd_sc_hd__clkbuf_1
X_1400_ outputs.divider_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2380_ _0802_ _0804_ _0658_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1262_ _0917_ net14 vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput6 gpio[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2716_ clknet_leaf_18_clk _0062_ net56 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_2647_ clknet_leaf_29_clk inputs.keypad\[8\] net32 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1529_ _1022_ outputs.shaper.count\[13\] _1110_ outputs.divider_buffer\[13\] vssd1
+ vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a2bb2o_1
X_2578_ clknet_leaf_36_clk net79 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1880_ _0381_ _0382_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__and3_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2501_ net287 outputs.sig_gen.count\[15\] _0861_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1314_ _0944_ _0947_ _0948_ _0949_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__nand4_2
XFILLER_0_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2432_ _0843_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
X_2294_ _0655_ _0723_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__or2_1
X_2363_ _0615_ _0676_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1245_ outputs.div.start vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ outputs.div.q\[21\] _0915_ _0405_ net141 _0414_ vssd1 vssd1 vccd1 vccd1 _0050_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1863_ _0359_ _0370_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1794_ _0288_ _0309_ _0299_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a21o_1
X_2415_ _0834_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2346_ _0773_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
X_2277_ _0491_ _0707_ _0653_ _0579_ _0577_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_32_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _0491_ _0494_ _0634_ _0592_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__a31o_1
X_2131_ _0537_ _0539_ _0544_ _0541_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__a31oi_1
X_2062_ _0494_ _0497_ _0499_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1915_ _0995_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__clkbuf_4
X_1846_ _0345_ _0351_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1777_ _0205_ _0293_ _0294_ _1228_ net181 vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2329_ _0747_ _0753_ _0757_ _0572_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2680_ clknet_leaf_12_clk _0026_ net57 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1700_ outputs.div.m\[5\] outputs.div.m\[4\] vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1631_ _1210_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__or2b_1
X_1493_ outputs.sig_gen.count\[15\] _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_1
X_1562_ _1108_ _1143_ _1114_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_3_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ _0475_ _0480_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _0545_ _0551_ _1215_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__mux2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout39 net43 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout28 net29 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1829_ net229 _0334_ outputs.div.next_div _0341_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2801_ clknet_leaf_2_clk _0119_ net41 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2594_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[1\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[1\] sky130_fd_sc_hd__dfrtp_1
X_2732_ clknet_leaf_12_clk outputs.div.next_start net52 vssd1 vssd1 vccd1 vccd1 outputs.div.start
+ sky130_fd_sc_hd__dfrtp_1
X_1614_ _1186_ _1190_ _1194_ outputs.output_gen.count\[7\] _1195_ vssd1 vssd1 vccd1
+ vccd1 _1196_ sky130_fd_sc_hd__o221a_1
X_2663_ clknet_leaf_30_clk _0009_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1476_ _1071_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
X_1545_ outputs.shaper.count\[1\] outputs.divider_buffer\[2\] vssd1 vssd1 vccd1 vccd1
+ _1127_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2028_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold250 outputs.divider_buffer\[17\] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1261_ _0922_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[4\] sky130_fd_sc_hd__clkbuf_1
X_1330_ _0964_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__and2b_1
Xinput7 gpio[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2646_ clknet_leaf_14_clk inputs.keypad\[7\] net58 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2715_ clknet_leaf_18_clk _0061_ net55 vssd1 vssd1 vccd1 vccd1 outputs.scaled_buffer\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2577_ clknet_leaf_36_clk net85 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1528_ outputs.shaper.count\[12\] vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1459_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2500_ _0869_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
X_2431_ outputs.divider_buffer\[8\] outputs.div.m\[8\] _0839_ vssd1 vssd1 vccd1 vccd1
+ _0843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1313_ inputs.random_update_clock.count\[6\] inputs.random_update_clock.count\[7\]
+ _0941_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__and3_1
X_1244_ outputs.div.count\[1\] outputs.div.count\[0\] outputs.div.count\[2\] vssd1
+ vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__a21o_1
X_2293_ _0653_ _0695_ _0481_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__o21a_1
X_2362_ _0472_ _0577_ _0787_ _0492_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2629_ clknet_leaf_15_clk net64 net58 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1931_ outputs.div.oscillator_out\[13\] _0411_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__and2_1
X_1862_ _0362_ _0367_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1793_ _0298_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 gpio[1] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_2414_ net311 outputs.div.m\[0\] _0798_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2345_ net285 _0772_ _0606_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__mux2_1
X_2276_ _0466_ _0470_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2130_ _0565_ _0567_ _0546_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__or3b_1
X_2061_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__buf_2
X_1914_ net167 _0400_ _0377_ net208 _0404_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1845_ _0342_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__buf_2
X_1776_ _0290_ _0292_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2328_ _0683_ _0756_ _1224_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2259_ _0556_ _0663_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1630_ inputs.octave_fsm.octave_key_up inputs.down.det_edge vssd1 vssd1 vccd1 vccd1
+ _1211_ sky130_fd_sc_hd__or2b_1
X_1492_ _1081_ _1079_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_1
X_1561_ _1115_ _1116_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2044_ _0481_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__clkbuf_4
X_2113_ _0548_ _0549_ _0550_ _0534_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__or4b_1
Xfanout29 net38 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_2
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1828_ _0339_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__xnor2_1
X_1759_ _0277_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2731_ clknet_leaf_17_clk outputs.div.next_div net59 vssd1 vssd1 vccd1 vccd1 outputs.div.div
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2800_ clknet_leaf_1_clk _0118_ net28 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2593_ clknet_leaf_14_clk inputs.random_update_clock.next_count\[0\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[0\] sky130_fd_sc_hd__dfstp_1
X_1544_ outputs.divider_buffer\[4\] _1124_ _1125_ outputs.divider_buffer\[3\] vssd1
+ vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__a22o_1
X_1613_ outputs.output_gen.count\[6\] _1189_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__or2_1
X_2662_ clknet_leaf_22_clk _0008_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1475_ _1041_ _1069_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2027_ inputs.frequency_lut.rng\[2\] vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold251 outputs.div.oscillator_out\[15\] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 outputs.div.a\[25\] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1260_ _0917_ net13 vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__and2b_1
Xinput8 gpio[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ clknet_leaf_12_clk _0060_ net52 vssd1 vssd1 vccd1 vccd1 outputs.div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2645_ clknet_leaf_6_clk inputs.keypad\[6\] net45 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1527_ _1006_ outputs.shaper.count\[8\] _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__a21o_1
X_2576_ clknet_leaf_36_clk net81 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1458_ outputs.sig_gen.count\[6\] _1055_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__and2_1
X_1389_ net145 _0907_ vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2430_ _0842_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2361_ _0581_ _0748_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__and2_1
X_1312_ _0952_ _0953_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
X_2292_ _0722_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
X_1243_ outputs.sample_rate.count\[7\] _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__nand2_4
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2628_ clknet_leaf_36_clk net90 net25 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2559_ _0699_ _0895_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1930_ net141 _0915_ _0405_ net187 _0413_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1861_ _0205_ _0368_ _0369_ _0333_ net238 vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a32o_1
X_1792_ _0306_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 gpio[2] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_2413_ net122 _0829_ _0833_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__a21o_1
X_2344_ _0464_ _0762_ _0771_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__a21o_1
X_2275_ net159 _1001_ _0694_ _0706_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2060_ inputs.frequency_lut.rng\[3\] vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__buf_2
X_1913_ outputs.div.oscillator_out\[5\] _0398_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1844_ _0345_ _0346_ _0351_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__or3_1
X_1775_ _0290_ _0292_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2258_ _0547_ _0689_ _0541_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__mux2_1
X_2327_ _0717_ _0755_ _0554_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2189_ _0464_ _0612_ _0618_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_62_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ _1121_ _1123_ _1141_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__and3b_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1491_ _1081_ _1079_ _1082_ _1042_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[14\]
+ sky130_fd_sc_hd__o211a_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2112_ _0515_ _0528_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2043_ inputs.frequency_lut.rng\[3\] vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1827_ _0328_ _0330_ _0326_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1758_ outputs.div.a\[10\] _0275_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1689_ _0205_ _0213_ _0214_ _1228_ net182 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a32o_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ clknet_leaf_19_clk net220 net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2661_ clknet_leaf_22_clk _0007_ net34 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1474_ outputs.sig_gen.count\[10\] _1068_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand2_1
X_1543_ outputs.shaper.count\[2\] vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__inv_2
X_1612_ _1191_ _1192_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2592_ clknet_leaf_29_clk _0002_ net32 vssd1 vssd1 vccd1 vccd1 inputs.octave_fsm.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2026_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2859_ clknet_leaf_6_clk _0177_ net45 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold252 outputs.div.oscillator_out\[12\] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 outputs.div.divisor\[8\] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 outputs.sample_rate.count\[7\] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 gpio[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2713_ clknet_leaf_13_clk _0059_ net57 vssd1 vssd1 vccd1 vccd1 outputs.div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2644_ clknet_leaf_23_clk inputs.keypad\[5\] net36 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1526_ _1006_ outputs.shaper.count\[8\] outputs.divider_buffer\[10\] _1107_ vssd1
+ vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a2bb2o_1
X_1457_ outputs.sig_gen.count\[6\] _1055_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__or2_1
X_2575_ clknet_leaf_36_clk net87 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1388_ _0907_ _0998_ vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
X_2009_ outputs.div.m\[10\] net285 _0453_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1311_ net237 _0941_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2291_ net282 _0721_ _0606_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__mux2_1
X_2360_ _0786_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1242_ outputs.sample_rate.count\[6\] _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2627_ clknet_leaf_24_clk net65 net34 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2489_ net272 outputs.sig_gen.count\[9\] _0861_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__mux2_1
X_1509_ net88 inputs.random_note_generator.out\[10\] vssd1 vssd1 vccd1 vccd1 _1095_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2558_ _0902_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_35_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1860_ _0360_ _0363_ _0367_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1791_ _0303_ _0305_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 gpio[3] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_2412_ _0830_ _0831_ _0832_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__a21oi_1
X_2274_ _0572_ _0701_ _0705_ _0910_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a31o_1
X_2343_ _0603_ _0770_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ _0444_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1843_ net251 _0334_ outputs.div.next_div _0353_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__a22o_1
X_1912_ outputs.div.q\[12\] _0400_ _0377_ net98 _0403_ vssd1 vssd1 vccd1 vccd1 _0041_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1774_ _0267_ _0270_ _0276_ _0278_ _0291_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2257_ _0536_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__and2_1
X_2326_ _0541_ _0735_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__o21ai_1
X_2188_ _0508_ _0623_ _0533_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1490_ _1081_ _1079_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1 inputs.keypad_synchronizer.half_sync\[12\] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ _0521_ _0538_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__nor2_1
X_2042_ _0477_ _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1826_ _0335_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1757_ outputs.div.a\[10\] _0275_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__nand2_2
X_1688_ _0208_ _0212_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__or2_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _0572_ _0733_ _0734_ _0738_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1611_ outputs.scaled_buffer\[7\] _1161_ _1165_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__a21oi_1
X_2660_ clknet_leaf_22_clk _0006_ net34 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1542_ outputs.shaper.count\[3\] vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__inv_2
X_1473_ outputs.sig_gen.count\[10\] _1068_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2591_ clknet_leaf_33_clk _0001_ net23 vssd1 vssd1 vccd1 vccd1 inputs.octave_fsm.state\[1\]
+ sky130_fd_sc_hd__dfstp_2
X_2025_ inputs.key_encoder.sync_keys\[13\] _1198_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold242 outputs.shaper.count\[7\] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
X_2858_ clknet_leaf_5_clk _0176_ net45 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold231 inputs.random_update_clock.count\[17\] vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1809_ outputs.div.a\[15\] vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__inv_2
Xhold253 outputs.div.oscillator_out\[2\] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlygate4sd3_1
X_2789_ clknet_leaf_0_clk _0107_ net26 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold220 outputs.div.divisor\[7\] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2643_ clknet_leaf_8_clk inputs.keypad\[4\] net49 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2712_ clknet_leaf_13_clk _0058_ net57 vssd1 vssd1 vccd1 vccd1 outputs.div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2574_ clknet_leaf_36_clk inputs.random_note_generator.feedback net24 vssd1 vssd1
+ vccd1 vccd1 inputs.random_note_generator.out\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1525_ outputs.shaper.count\[9\] vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__inv_2
X_1456_ _1055_ _1056_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_22_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1387_ net152 _0906_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__nor2_1
X_2008_ _0454_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1310_ inputs.random_update_clock.count\[6\] _0941_ vssd1 vssd1 vccd1 vccd1 _0952_
+ sky130_fd_sc_hd__and2_1
X_2290_ _0714_ _0720_ _0603_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__mux2_1
X_1241_ outputs.sample_rate.count\[4\] outputs.sample_rate.count\[5\] _0907_ vssd1
+ vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2626_ clknet_leaf_14_clk net78 net58 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2557_ _0901_ _0492_ _0895_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ _0863_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__clkbuf_1
X_1439_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] vssd1 vssd1 vccd1 vccd1
+ _1044_ sky130_fd_sc_hd__nand2_1
X_1508_ _1093_ inputs.random_note_generator.out\[13\] vssd1 vssd1 vccd1 vccd1 _1094_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 gpio[4] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1790_ _0303_ _0305_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__or2_1
X_2411_ _0910_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2342_ _0767_ _0769_ _0508_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__mux2_1
X_2273_ _0703_ _0704_ _0658_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1988_ outputs.div.m\[0\] net283 _0436_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2609_ clknet_leaf_17_clk inputs.random_update_clock.next_count\[16\] net55 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1842_ _0351_ _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1911_ outputs.div.oscillator_out\[4\] _0398_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__and2_1
X_1773_ _0281_ _0276_ _0277_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2187_ _0586_ _0585_ _0619_ _0622_ _0616_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__o32a_1
X_2325_ _0515_ _0524_ _0536_ _0531_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__o211a_2
X_2256_ _0543_ _0535_ _0557_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 inputs.keypad_synchronizer.half_sync\[7\] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2041_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__buf_2
X_2110_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1825_ outputs.div.m\[17\] _0337_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__xnor2_2
X_1756_ _0274_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1687_ _0208_ _0212_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2308_ _1207_ _0737_ _0603_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__o21a_1
X_2239_ _0491_ _0636_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1610_ outputs.scaled_buffer\[6\] net21 _1163_ _1158_ vssd1 vssd1 vccd1 vccd1 _1192_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ clknet_leaf_29_clk _0000_ net32 vssd1 vssd1 vccd1 vccd1 inputs.octave_fsm.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1541_ outputs.divider_buffer\[8\] _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__or2_1
X_1472_ _1011_ _1065_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2024_ _0462_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
X_2857_ clknet_leaf_7_clk _0175_ net45 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold243 outputs.shaper.count\[17\] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold210 outputs.div.oscillator_out\[9\] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1808_ net228 _0916_ outputs.div.next_div _0322_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1739_ outputs.div.a\[8\] _0258_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__or2_1
Xhold221 outputs.div.divisor\[0\] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 outputs.div.divisor\[5\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
X_2788_ clknet_leaf_36_clk _0106_ net26 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2711_ clknet_leaf_13_clk _0057_ net57 vssd1 vssd1 vccd1 vccd1 outputs.div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1524_ _1102_ _1104_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__or3b_1
X_2573_ clknet_leaf_24_clk net255 net34 vssd1 vssd1 vccd1 vccd1 inputs.wavetype_fsm.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2642_ clknet_leaf_33_clk inputs.keypad\[3\] net23 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1455_ net307 _1053_ _1042_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__o21ai_1
X_1386_ _0906_ net157 vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
X_2007_ outputs.div.m\[9\] net295 _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1240_ outputs.sample_rate.count\[3\] _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2487_ net269 outputs.sig_gen.count\[8\] _0861_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1507_ inputs.random_note_generator.out\[15\] vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__buf_2
X_2625_ clknet_leaf_29_clk net66 net32 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2556_ _0467_ _1093_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1438_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] vssd1 vssd1 vccd1 vccd1
+ _1043_ sky130_fd_sc_hd__or2_1
X_1369_ net245 _0986_ vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[4\] sky130_fd_sc_hd__xor2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput14 gpio[5] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2410_ _0658_ _0699_ _0464_ _0792_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__or4_1
X_2341_ _0615_ _0577_ _0768_ _0656_ _0648_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__a32o_1
X_2272_ _0492_ _0487_ _0497_ _0647_ _0699_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a311o_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1987_ net219 _0439_ _0443_ outputs.div.q\[7\] vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__o22a_1
X_2608_ clknet_leaf_16_clk inputs.random_update_clock.next_count\[15\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[15\] sky130_fd_sc_hd__dfrtp_1
X_2539_ _0889_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1910_ net98 _0400_ _0377_ net183 _0402_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1841_ _0345_ _0349_ _0343_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1772_ _0288_ _0289_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2324_ _0506_ _0750_ _0752_ _0603_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2186_ _0482_ _0494_ _0620_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__a31o_1
X_2255_ _0515_ _0523_ _0527_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 inputs.keypad_synchronizer.half_sync\[5\] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ inputs.frequency_lut.rng\[2\] _0469_ _0471_ vssd1 vssd1 vccd1 vccd1 _0478_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ clknet_leaf_24_clk net75 net35 vssd1 vssd1 vccd1 vccd1 outputs.pwm_output
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1824_ _0248_ _0336_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__and2_1
X_1755_ outputs.div.m\[11\] _0273_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__xnor2_1
X_1686_ outputs.div.a\[3\] _0211_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__xnor2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2238_ _0669_ _0582_ _0670_ _0505_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__a211o_1
X_2307_ _0690_ _0736_ _0554_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2169_ _0411_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1540_ outputs.shaper.count\[7\] vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1471_ _1011_ _1065_ _1067_ _1042_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[9\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2023_ outputs.div.m\[17\] net122 _0453_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__mux2_1
X_2856_ clknet_leaf_9_clk _0174_ net47 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1807_ _0320_ _0321_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold244 outputs.div.oscillator_out\[13\] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 outputs.div.oscillator_out\[14\] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 outputs.div.q\[6\] vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _1225_ _0195_ _0196_ _1228_ net231 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a32o_1
X_1738_ outputs.div.a\[8\] _0258_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__and2_1
Xhold233 outputs.div.divisor\[9\] vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
X_2787_ clknet_leaf_0_clk _0105_ net25 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold211 outputs.div.divisor\[4\] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2710_ clknet_leaf_13_clk _0056_ net58 vssd1 vssd1 vccd1 vccd1 outputs.div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1523_ _1103_ outputs.shaper.count\[15\] vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__nand2_1
X_1454_ outputs.sig_gen.count\[4\] outputs.sig_gen.count\[5\] _1049_ vssd1 vssd1 vccd1
+ vccd1 _1055_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2572_ clknet_leaf_24_clk inputs.wavetype_fsm.next_state\[0\] net30 vssd1 vssd1 vccd1
+ vccd1 inputs.wavetype_fsm.state\[0\] sky130_fd_sc_hd__dfrtp_1
X_2641_ clknet_leaf_27_clk inputs.keypad\[2\] net31 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1385_ net148 outputs.sample_rate.count\[0\] net156 vssd1 vssd1 vccd1 vccd1 _0997_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2006_ _0411_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2839_ clknet_leaf_5_clk _0157_ net44 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2624_ clknet_leaf_28_clk net72 net32 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2486_ _0862_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__clkbuf_1
X_1437_ net248 _1042_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[0\] sky130_fd_sc_hd__nand2_1
X_1506_ inputs.wavetype_fsm.state\[1\] _1090_ vssd1 vssd1 vccd1 vccd1 inputs.wavetype_fsm.next_state\[1\]
+ sky130_fd_sc_hd__xnor2_1
X_2555_ _0900_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1299_ inputs.random_update_clock.count\[4\] inputs.random_update_clock.count\[6\]
+ inputs.random_update_clock.count\[7\] inputs.random_update_clock.count\[5\] vssd1
+ vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1368_ _0986_ _0987_ vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_53_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 gpio[6] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2340_ _0477_ _0707_ _0485_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__o21ai_1
X_2271_ _0702_ _0506_ _0589_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1986_ net198 _0439_ _0443_ outputs.div.q\[6\] vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2607_ clknet_leaf_16_clk inputs.random_update_clock.next_count\[14\] net61 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2469_ net111 _0832_ _0418_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__a21o_1
X_2538_ outputs.shaper.count\[15\] net135 _0396_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1840_ outputs.div.a\[18\] _0342_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1771_ _0284_ _0287_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2254_ _0686_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
X_2323_ _0492_ _0494_ _0751_ _0658_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__o211ai_1
X_2185_ _0498_ _0471_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ outputs.scaled_buffer\[6\] outputs.div.q_out\[6\] _1001_ vssd1 vssd1 vccd1
+ vccd1 _0435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 inputs.keypad_synchronizer.half_sync\[3\] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1823_ outputs.div.m\[16\] outputs.div.m\[15\] _0314_ vssd1 vssd1 vccd1 vccd1 _0336_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_29_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2872_ clknet_leaf_35_clk _0190_ net23 vssd1 vssd1 vccd1 vccd1 inputs.frequency_lut.rng\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_1754_ outputs.div.m\[10\] _0249_ _0264_ _0248_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__o31a_1
X_1685_ outputs.div.m\[4\] _0210_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__xor2_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2237_ _0498_ _0468_ _0588_ _0592_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__a31o_1
X_2306_ _0715_ _0735_ _0541_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2099_ _0530_ _0528_ _0536_ _0531_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__o211a_1
X_2168_ _0464_ _0595_ _0601_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1470_ outputs.sig_gen.count\[9\] _1064_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2022_ _0461_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2855_ clknet_leaf_9_clk _0173_ net47 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1806_ _0308_ _0311_ _0306_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 _0036_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2786_ clknet_leaf_0_clk _0104_ net25 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold234 inputs.random_update_clock.count\[5\] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 outputs.div.oscillator_out\[4\] vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold245 outputs.sig_gen.count\[5\] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
X_1599_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] outputs.scaled_buffer\[2\]
+ net21 vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__o31a_1
X_1668_ _1236_ _0194_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__or2_1
X_1737_ outputs.div.m\[9\] _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__xor2_1
Xhold223 outputs.div.divisor\[10\] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ clknet_leaf_34_clk inputs.keypad\[1\] net22 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1522_ _1103_ outputs.shaper.count\[15\] _1101_ outputs.divider_buffer\[15\] vssd1
+ vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1453_ _1053_ _1054_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[4\] sky130_fd_sc_hd__nor2_1
X_2571_ clknet_leaf_22_clk outputs.sample_rate.next_count\[7\] net34 vssd1 vssd1 vccd1
+ vccd1 outputs.sample_rate.count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ _0452_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1384_ net148 net133 vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2838_ clknet_leaf_7_clk _0156_ net46 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2769_ clknet_leaf_0_clk _0087_ net25 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2623_ clknet_leaf_29_clk net82 net32 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2554_ _0899_ _0467_ _0895_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2485_ net277 outputs.sig_gen.count\[7\] _0861_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__mux2_1
X_1436_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__buf_2
X_1367_ net261 _0984_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__nor2_1
X_1505_ _1092_ vssd1 vssd1 vccd1 vccd1 inputs.wavetype_fsm.next_state\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1298_ inputs.random_update_clock.count\[4\] inputs.random_update_clock.count\[5\]
+ _0938_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 gpio[7] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2270_ _0502_ _0647_ _0499_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ net162 _0439_ _0443_ outputs.div.q\[5\] vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2537_ _0888_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
X_2606_ clknet_leaf_16_clk inputs.random_update_clock.next_count\[13\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2468_ net126 _0832_ _0417_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1419_ _1022_ outputs.sig_gen.count\[14\] outputs.divider_buffer\[16\] _1023_ _1024_
+ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__a221o_1
X_2399_ net239 _0821_ _0798_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ _0284_ _0287_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__or2_1
X_2253_ net294 _0685_ _0606_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__mux2_1
X_2184_ _0468_ _0466_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__nand2_1
X_2322_ _0485_ _0479_ _0502_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1899_ outputs.div.q\[7\] _1228_ _1225_ net262 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__a22o_1
X_1968_ _0434_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 inputs.keypad_synchronizer.half_sync\[14\] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1822_ outputs.div.a\[16\] vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1753_ _0205_ _0271_ _0272_ _1228_ net180 vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2871_ clknet_leaf_35_clk _0189_ net23 vssd1 vssd1 vccd1 vccd1 inputs.frequency_lut.rng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1684_ _1229_ _0209_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _0486_ _0467_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__or2_1
X_2167_ _1224_ _0602_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__o21ai_1
X_2305_ _0527_ _0539_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2098_ _0534_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2021_ outputs.div.m\[16\] net232 _0453_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold213 outputs.div.oscillator_out\[11\] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
X_2854_ clknet_leaf_13_clk _0172_ net47 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold202 outputs.div.oscillator_out\[6\] vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__dlygate4sd3_1
X_1805_ _0318_ _0319_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1736_ outputs.div.m\[8\] _0249_ _1229_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__o21a_1
Xhold224 outputs.div.divisor\[13\] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2785_ clknet_leaf_31_clk _0103_ net29 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold235 outputs.div.m\[6\] vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ _1236_ _0194_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__nand2_1
Xhold246 outputs.scaled_buffer\[7\] vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlygate4sd3_1
X_1598_ outputs.output_gen.count\[3\] _1170_ _1174_ outputs.output_gen.count\[2\]
+ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__o221a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _0469_ _0471_ _0465_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2570_ clknet_leaf_25_clk outputs.sample_rate.next_count\[6\] net30 vssd1 vssd1 vccd1
+ vccd1 outputs.sample_rate.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1521_ outputs.divider_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__inv_2
X_1452_ outputs.sig_gen.count\[4\] _1049_ _1042_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1383_ net133 vssd1 vssd1 vccd1 vccd1 outputs.sample_rate.next_count\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2004_ outputs.div.m\[8\] net292 _0436_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2699_ clknet_leaf_7_clk net151 net46 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2837_ clknet_leaf_10_clk _0155_ net42 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2768_ clknet_leaf_0_clk _0086_ net26 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_1719_ _0240_ _0241_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__or2_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1504_ _1090_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__and2_1
X_2622_ clknet_leaf_25_clk net94 net30 vssd1 vssd1 vccd1 vccd1 inputs.key_encoder.sync_keys\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2553_ _0473_ _1093_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__xor2_1
X_2484_ _0994_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__clkbuf_4
X_1435_ _1016_ _1021_ _1025_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__or4_4
X_1366_ outputs.output_gen.count\[3\] _0984_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1297_ inputs.random_update_clock.count\[4\] _0938_ net296 vssd1 vssd1 vccd1 vccd1
+ _0940_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput17 gpio[8] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1984_ net174 _0439_ _0443_ outputs.div.q\[4\] vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2536_ outputs.shaper.count\[14\] net106 _0396_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__mux2_1
X_2605_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[12\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[12\] sky130_fd_sc_hd__dfrtp_1
X_2467_ net135 _0832_ _0416_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1349_ net218 _0977_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[19\]
+ sky130_fd_sc_hd__xor2_1
X_1418_ outputs.divider_buffer\[2\] outputs.sig_gen.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1024_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _1208_ _0464_ _0782_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2321_ _0497_ _0748_ _0749_ _0621_ _0650_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__a311o_1
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2183_ _0616_ _0576_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__nand2_1
X_2252_ _0572_ _0680_ _0681_ _0684_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1898_ outputs.div.q\[6\] _0334_ _1225_ net258 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__a22o_1
X_1967_ outputs.scaled_buffer\[5\] net162 _1001_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__mux2_1
X_2519_ _0879_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 inputs.random_note_generator.out\[7\] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2870_ clknet_leaf_34_clk _0188_ net22 vssd1 vssd1 vccd1 vccd1 inputs.frequency_lut.rng\[3\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1821_ _0915_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1752_ _0267_ _0270_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__or2_1
X_1683_ outputs.div.m\[3\] outputs.div.m\[2\] outputs.div.m\[0\] outputs.div.m\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__or4_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2304_ _1208_ _0664_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _0668_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__clkbuf_1
X_2097_ _0530_ _0523_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__nand2_1
X_2166_ _0463_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2020_ _0460_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2853_ clknet_leaf_2_clk _0171_ net43 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold236 outputs.shaper.count\[11\] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 outputs.div.oscillator_out\[10\] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 outputs.div.oscillator_out\[15\] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
X_1804_ outputs.div.a\[14\] _0317_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__or2_1
Xhold203 outputs.div.oscillator_out\[0\] vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 outputs.divider_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1666_ _0192_ _0193_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__nand2_1
X_1735_ _0255_ _0256_ net192 _0916_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a2bb2o_1
X_2784_ clknet_leaf_0_clk _0102_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ outputs.output_gen.count\[2\] _1174_ _1176_ _1178_ vssd1 vssd1 vccd1 vccd1
+ _1179_ sky130_fd_sc_hd__a22o_1
X_2149_ _0486_ inputs.frequency_lut.rng\[1\] inputs.frequency_lut.rng\[2\] vssd1 vssd1
+ vccd1 vccd1 _0586_ sky130_fd_sc_hd__a21oi_4
X_2218_ _0646_ _0649_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1520_ outputs.divider_buffer\[15\] _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1451_ outputs.sig_gen.count\[4\] _1049_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__and2_1
X_1382_ _0996_ vssd1 vssd1 vccd1 vccd1 outputs.div.next_div sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2003_ _0451_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2836_ clknet_leaf_10_clk _0154_ net46 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2698_ clknet_leaf_9_clk net197 net46 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1649_ outputs.div.m\[0\] outputs.div.q\[26\] vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__or2_1
X_2767_ clknet_leaf_31_clk _0085_ net37 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_1718_ _0237_ _0239_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__and2_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2483_ _0860_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1503_ inputs.wavetype_fsm.state\[0\] inputs.mode_edge.det_edge vssd1 vssd1 vccd1
+ vccd1 _1091_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2621_ clknet_leaf_28_clk inputs.up.ff_in net31 vssd1 vssd1 vccd1 vccd1 inputs.octave_fsm.octave_key_up
+ sky130_fd_sc_hd__dfrtp_1
X_2552_ _0898_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1296_ net200 _0938_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
X_1434_ _1029_ _1032_ _1036_ _1039_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1365_ _0984_ net242 vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_0_65_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2819_ clknet_leaf_9_clk net102 net46 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 gpio[9] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2604_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[11\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1983_ net170 _0439_ _0443_ outputs.div.q\[3\] vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2535_ _0887_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
X_2466_ net106 _0832_ _0415_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1417_ outputs.sig_gen.count\[16\] vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1348_ _0951_ _0976_ _0977_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[18\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1279_ _0931_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[13\] sky130_fd_sc_hd__clkbuf_1
X_2397_ _0817_ _0819_ _0533_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2320_ _0498_ _0479_ _0502_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__or3_1
X_2251_ _1224_ _0683_ _0533_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2182_ _0613_ _0614_ _0617_ _0508_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1966_ _0433_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1897_ net258 _0334_ _1225_ net260 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2518_ outputs.shaper.count\[5\] net123 _0872_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__mux2_1
X_2449_ _0852_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7 inputs.random_note_generator.out\[5\] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ _0205_ _0331_ _0332_ _0333_ net172 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1751_ _0267_ _0270_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__nand2_1
X_1682_ _0201_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ net273 _0667_ _0606_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2303_ _0724_ _0726_ _0729_ _0732_ _0616_ _0650_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2165_ _0532_ _0559_ _0563_ _0568_ _1215_ _0556_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__mux4_1
X_2096_ _0533_ _0517_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1949_ _0911_ _0377_ _0423_ _0333_ net176 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2852_ clknet_leaf_11_clk _0170_ net43 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1803_ outputs.div.a\[14\] _0317_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2783_ clknet_leaf_30_clk _0101_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold237 outputs.shaper.count\[12\] vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 outputs.div.oscillator_out\[7\] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 outputs.div.a\[18\] vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 outputs.divider_buffer\[14\] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1665_ _1237_ _0191_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__nand2_1
X_1734_ _0246_ _0254_ _0996_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__a21bo_1
X_1596_ outputs.output_gen.count\[1\] _1175_ _1177_ outputs.output_gen.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a211o_1
Xhold226 outputs.div.divisor\[11\] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2217_ _0646_ _0649_ _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2148_ inputs.frequency_lut.rng\[0\] inputs.frequency_lut.rng\[1\] inputs.frequency_lut.rng\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__and3_4
X_2079_ inputs.key_encoder.sync_keys\[12\] _1199_ _1202_ _0516_ vssd1 vssd1 vccd1
+ vccd1 _0517_ sky130_fd_sc_hd__o31a_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1450_ _1052_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1381_ _0995_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2002_ outputs.div.m\[7\] net282 _0436_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2835_ clknet_leaf_3_clk _0153_ net39 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2766_ clknet_leaf_0_clk _0084_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2697_ clknet_leaf_9_clk net168 net46 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1648_ outputs.div.m\[0\] outputs.div.q\[26\] vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__nand2_1
X_1579_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__buf_2
X_1717_ _0237_ _0239_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__nor2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2620_ clknet_leaf_28_clk net92 net30 vssd1 vssd1 vccd1 vccd1 inputs.up.ff_out sky130_fd_sc_hd__dfrtp_1
X_2482_ net264 outputs.sig_gen.count\[6\] _0850_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__mux2_1
X_1433_ _1037_ outputs.sig_gen.count\[7\] _1014_ outputs.sig_gen.count\[10\] _1038_
+ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__a221o_1
X_1502_ inputs.wavetype_fsm.state\[0\] net254 vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__nand2_1
X_2551_ _0897_ _0473_ _0895_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__mux2_1
X_1295_ _0938_ _0939_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
X_1364_ outputs.output_gen.count\[1\] net100 net241 vssd1 vssd1 vccd1 vccd1 _0985_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2818_ clknet_leaf_13_clk net124 net46 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2749_ clknet_leaf_4_clk outputs.sig_gen.next_count\[8\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 nrst vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_2
XFILLER_0_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1982_ net160 _0439_ _0443_ outputs.div.q\[2\] vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__o22a_1
X_2534_ outputs.shaper.count\[13\] net114 _0396_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__mux2_1
X_2603_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[10\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2465_ net114 _0832_ _0414_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__a21o_1
X_1347_ inputs.random_update_clock.count\[18\] _0975_ vssd1 vssd1 vccd1 vccd1 _0977_
+ sky130_fd_sc_hd__and2_1
X_1416_ outputs.divider_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__inv_2
X_2396_ _0803_ _0818_ _0508_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire21 _1155_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_4
X_1278_ net1 net9 vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ _0629_ _0682_ _0554_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2181_ _0499_ _0489_ _0496_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1965_ outputs.scaled_buffer\[4\] net174 _1001_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2517_ _0878_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
X_1896_ outputs.div.q\[4\] _0334_ _1225_ net252 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2448_ outputs.divider_buffer\[16\] outputs.div.m\[16\] _0850_ vssd1 vssd1 vccd1
+ vccd1 _0852_ sky130_fd_sc_hd__mux2_1
X_2379_ _0579_ _0676_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 inputs.random_note_generator.out\[8\] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1750_ _0246_ _0254_ _0268_ _0269_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1681_ _1236_ _0194_ _0206_ _0192_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _1207_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__nor2_1
X_2233_ _0603_ _0652_ _0659_ _0665_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__o32a_1
X_2302_ _0482_ _0730_ _0731_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2095_ inputs.key_encoder.sync_keys\[13\] _1198_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__and2_2
XFILLER_0_75_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1948_ _0422_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1879_ _0383_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1802_ _0316_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
X_2851_ clknet_leaf_11_clk _0169_ net42 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1733_ _0246_ _0254_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2782_ clknet_leaf_31_clk _0100_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold227 outputs.div.oscillator_out\[12\] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 outputs.div.oscillator_out\[3\] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold238 outputs.shaper.count\[1\] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold249 outputs.divider_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1595_ outputs.scaled_buffer\[0\] _1161_ _1165_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__a21oi_1
X_1664_ _1237_ _0191_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__or2_1
Xhold216 outputs.div.a\[3\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2147_ _0491_ _0479_ _0579_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2216_ inputs.frequency_lut.rng\[5\] vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2078_ inputs.key_encoder.sync_keys\[13\] _1198_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1380_ _0994_ _0913_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2001_ _0450_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2696_ clknet_leaf_13_clk net209 net57 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2834_ clknet_leaf_10_clk _0152_ net42 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1716_ outputs.div.m\[7\] _0238_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__xnor2_1
X_2765_ clknet_leaf_30_clk _0083_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1647_ _0996_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__clkbuf_4
X_1578_ inputs.wavetype_fsm.state\[0\] inputs.wavetype_fsm.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _1160_ sky130_fd_sc_hd__and2b_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2550_ _0486_ _1093_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__xor2_1
X_2481_ _0859_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
X_1501_ net207 _1088_ _1089_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[17\]
+ sky130_fd_sc_hd__a21oi_1
X_1432_ _1018_ outputs.sig_gen.count\[15\] _1030_ outputs.sig_gen.count\[6\] vssd1
+ vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1363_ outputs.output_gen.count\[2\] outputs.output_gen.count\[1\] outputs.output_gen.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1294_ net212 _0936_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2679_ clknet_leaf_13_clk _0025_ net57 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_2748_ clknet_leaf_4_clk outputs.sig_gen.next_count\[7\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[7\] sky130_fd_sc_hd__dfrtp_4
X_2817_ clknet_leaf_2_clk _0135_ net42 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1981_ net154 _0439_ _0443_ outputs.div.q\[1\] vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__o22a_1
X_2533_ _0886_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2602_ clknet_leaf_15_clk inputs.random_update_clock.next_count\[9\] net60 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2464_ net103 _0832_ _0413_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__a21o_1
X_1346_ inputs.random_update_clock.count\[18\] _0975_ vssd1 vssd1 vccd1 vccd1 _0976_
+ sky130_fd_sc_hd__nor2_1
X_1415_ _1017_ outputs.sig_gen.count\[3\] _1018_ outputs.sig_gen.count\[15\] _1020_
+ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2395_ _0585_ _0731_ _0505_ _0487_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1277_ _0930_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2180_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1895_ outputs.div.q\[3\] _0334_ _1225_ net233 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__a22o_1
X_1964_ _0432_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2447_ _0851_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__clkbuf_1
X_2516_ outputs.shaper.count\[4\] net105 _0872_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1329_ inputs.random_update_clock.count\[11\] inputs.random_update_clock.count\[10\]
+ _0959_ inputs.random_update_clock.count\[12\] vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2378_ _0498_ _0487_ _0505_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold9 inputs.keypad_synchronizer.half_sync\[9\] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1680_ outputs.div.a\[2\] _0199_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2301_ _0484_ _0474_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__and2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2163_ _0598_ _0599_ _0556_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__mux2_1
X_2232_ _1224_ _0555_ _0603_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2094_ _0515_ _0524_ _0528_ _0529_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1947_ outputs.div.count\[2\] outputs.div.count\[1\] outputs.div.count\[0\] vssd1
+ vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1878_ outputs.div.a\[23\] _0355_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2850_ clknet_leaf_2_clk _0168_ net41 vssd1 vssd1 vccd1 vccd1 outputs.shaper.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1801_ outputs.div.m\[15\] _0315_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__xor2_1
Xhold217 outputs.div.oscillator_out\[2\] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 outputs.div.a\[9\] vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlygate4sd3_1
X_1663_ outputs.div.m\[2\] _1238_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__xnor2_1
X_1732_ _0252_ _0253_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2781_ clknet_leaf_32_clk _0099_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold228 outputs.div.oscillator_out\[17\] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 outputs.shaper.count\[8\] vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ outputs.output_gen.count\[1\] _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2077_ inputs.key_encoder.sync_keys\[10\] _0514_ inputs.key_encoder.sync_keys\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__o21bai_4
X_2146_ _0491_ _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__nand2_1
X_2215_ _0485_ _0647_ _0648_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2000_ outputs.div.m\[6\] net159 _0436_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__mux2_1
X_2833_ clknet_leaf_2_clk _0151_ net41 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2695_ clknet_leaf_13_clk net99 net57 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1715_ outputs.div.m\[6\] _0209_ _0224_ _1229_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__o31a_1
X_2764_ clknet_leaf_31_clk _0082_ net33 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_1646_ _1211_ _1224_ _1220_ _1210_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1577_ outputs.scaled_buffer\[4\] _1099_ net21 _1158_ vssd1 vssd1 vccd1 vccd1 _1159_
+ sky130_fd_sc_hd__a31o_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2129_ _0526_ _0521_ _0522_ _0566_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__a31o_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1500_ net207 _1088_ _1042_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__o21ai_1
X_2480_ net270 outputs.sig_gen.count\[5\] _0850_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1293_ inputs.random_update_clock.count\[3\] _0936_ vssd1 vssd1 vccd1 vccd1 _0938_
+ sky130_fd_sc_hd__and2_1
X_1431_ outputs.divider_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__inv_2
X_1362_ net153 net100 vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2816_ clknet_leaf_12_clk net109 net42 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2678_ clknet_leaf_14_clk _0024_ net57 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_2747_ clknet_leaf_4_clk outputs.sig_gen.next_count\[6\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1629_ inputs.down.det_edge inputs.octave_fsm.octave_key_up vssd1 vssd1 vccd1 vccd1
+ _1210_ sky130_fd_sc_hd__and2b_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ net164 _0439_ _0443_ outputs.div.q\[0\] vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2532_ net299 net103 _0396_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__mux2_1
X_2463_ net112 _0832_ _0412_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__a21o_1
X_2601_ clknet_leaf_17_clk inputs.random_update_clock.next_count\[8\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1345_ _0951_ _0974_ _0975_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[17\]
+ sky130_fd_sc_hd__nor3_1
X_1414_ _1019_ outputs.sig_gen.count\[5\] _1007_ outputs.sig_gen.count\[17\] vssd1
+ vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1276_ net1 net5 vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2394_ _0650_ _0616_ _0499_ _0647_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1894_ net233 _0334_ _1225_ net244 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__a22o_1
X_1963_ outputs.scaled_buffer\[3\] net170 _1001_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2515_ _0877_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
X_2446_ outputs.divider_buffer\[15\] outputs.div.m\[15\] _0850_ vssd1 vssd1 vccd1
+ vccd1 _0851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1328_ inputs.random_update_clock.count\[11\] inputs.random_update_clock.count\[10\]
+ inputs.random_update_clock.count\[12\] _0959_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1259_ _0921_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[3\] sky130_fd_sc_hd__clkbuf_1
X_2377_ _0485_ _0480_ _0741_ _0506_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2300_ _0470_ _0477_ _0695_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a21o_1
X_2231_ _1207_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__nor2_1
X_2162_ _0540_ _0551_ _0541_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__mux2_1
X_2093_ _0517_ _0521_ _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__or3_4
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1946_ _0420_ _0377_ _0421_ _0333_ net246 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__a32o_1
X_1877_ outputs.div.a\[23\] _0355_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__nand2_1
X_2429_ outputs.divider_buffer\[7\] outputs.div.m\[7\] _0839_ vssd1 vssd1 vccd1 vccd1
+ _0842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1800_ _0248_ _0314_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__nand2_1
Xhold229 outputs.div.oscillator_out\[16\] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold207 outputs.div.oscillator_out\[8\] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__dlygate4sd3_1
X_1731_ _0247_ _0251_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__and2_1
X_1662_ outputs.div.m\[0\] outputs.div.m\[1\] outputs.div.a\[25\] vssd1 vssd1 vccd1
+ vccd1 _1238_ sky130_fd_sc_hd__o21ba_1
Xhold218 outputs.div.divisor\[1\] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
X_2780_ clknet_leaf_32_clk _0098_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.divisor\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ outputs.scaled_buffer\[0\] _1157_ _1161_ outputs.scaled_buffer\[1\] _1165_
+ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2214_ _0484_ _0494_ _0620_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nand3_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2076_ inputs.key_encoder.sync_keys\[8\] _0513_ inputs.key_encoder.sync_keys\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__o21ba_1
X_2145_ _0580_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__and2_1
X_1929_ net314 _0411_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 outputs.sample_rate.count\[3\] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dlygate4sd3_1
X_2832_ clknet_leaf_2_clk _0150_ net41 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2763_ clknet_leaf_32_clk _0081_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_2694_ clknet_leaf_12_clk net184 net52 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1576_ _1157_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__inv_2
X_1714_ outputs.div.a\[6\] vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__inv_2
X_1645_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _0467_ _0470_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2128_ _0539_ _0561_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__nand2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1430_ _1033_ outputs.sig_gen.count\[0\] _1034_ outputs.sig_gen.count\[11\] _1035_
+ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1292_ _0936_ net203 vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1361_ net100 vssd1 vssd1 vccd1 vccd1 outputs.output_gen.next_count\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_73_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2815_ clknet_leaf_11_clk _0133_ net42 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2746_ clknet_leaf_4_clk outputs.sig_gen.next_count\[5\] net39 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2677_ clknet_leaf_14_clk _0023_ net57 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1559_ _1137_ _1138_ _1139_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1628_ inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _1209_ sky130_fd_sc_hd__or2b_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2600_ clknet_leaf_17_clk inputs.random_update_clock.next_count\[7\] net59 vssd1
+ vssd1 vccd1 vccd1 inputs.random_update_clock.count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2531_ _0885_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
X_2462_ net131 _0832_ _0410_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__a21o_1
X_1413_ outputs.divider_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__inv_2
X_2393_ _0816_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1344_ inputs.random_update_clock.count\[16\] inputs.random_update_clock.count\[17\]
+ _0972_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__and3_1
X_1275_ _0929_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2729_ clknet_leaf_19_clk net199 net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1962_ _0431_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1893_ net244 _0334_ _1225_ net257 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2514_ outputs.shaper.count\[3\] net108 _0872_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__mux2_1
X_2445_ _0994_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__buf_4
X_2376_ _0699_ _0698_ _0792_ _0789_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__a31o_1
X_1327_ net221 _0961_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[11\]
+ sky130_fd_sc_hd__xnor2_1
X_1258_ _0917_ net12 vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2230_ _0609_ _0663_ _0554_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2161_ _0545_ _0597_ _1214_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__mux2_1
X_2092_ _0515_ _0522_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1945_ outputs.div.count\[1\] outputs.div.count\[0\] vssd1 vssd1 vccd1 vccd1 _0421_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_61_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1876_ outputs.div.a\[22\] outputs.div.a\[21\] outputs.div.a\[20\] outputs.div.a\[19\]
+ _0355_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o41ai_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2428_ _0841_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
X_2359_ net288 _0785_ _0606_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold208 outputs.div.oscillator_out\[5\] vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 outputs.div.oscillator_out\[1\] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1661_ outputs.div.a\[1\] vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__inv_2
X_1592_ _1171_ _1172_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__o21a_1
X_1730_ _0247_ _0251_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _0465_ _0471_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__nand2_2
X_2213_ _0473_ _0465_ _0486_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__and3b_2
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2075_ inputs.key_encoder.sync_keys\[6\] _0512_ inputs.key_encoder.sync_keys\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__o21ba_1
X_1928_ net187 _0400_ _0405_ net193 _0412_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1859_ _0360_ _0363_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold80 _0050_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 outputs.output_gen.count\[1\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2831_ clknet_leaf_3_clk _0149_ net39 vssd1 vssd1 vccd1 vccd1 outputs.div.oscillator_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2762_ clknet_leaf_31_clk _0080_ net28 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1713_ _0205_ _0235_ _0236_ _1228_ net190 vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2693_ clknet_leaf_12_clk _0039_ net52 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1575_ inputs.wavetype_fsm.state\[1\] inputs.wavetype_fsm.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _1157_ sky130_fd_sc_hd__nor2b_2
X_1644_ inputs.octave_fsm.state\[2\] _1205_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__and2_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _0531_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _0494_ _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__nand2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1360_ _0983_ vssd1 vssd1 vccd1 vccd1 inputs.down.in sky130_fd_sc_hd__clkbuf_1
X_1291_ inputs.random_update_clock.count\[1\] inputs.random_update_clock.count\[0\]
+ net202 vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2676_ clknet_leaf_17_clk _0022_ net59 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_2745_ clknet_leaf_3_clk outputs.sig_gen.next_count\[4\] net39 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[4\] sky130_fd_sc_hd__dfrtp_2
X_2814_ clknet_leaf_2_clk _0132_ net41 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1489_ outputs.sig_gen.count\[14\] vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__inv_2
X_1558_ _1037_ outputs.shaper.count\[6\] outputs.divider_buffer\[8\] _1122_ vssd1
+ vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__a2bb2o_1
X_1627_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__buf_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2530_ net298 net112 _0396_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2461_ net116 _0832_ _0409_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__a21o_1
X_1343_ inputs.random_update_clock.count\[16\] _0972_ net293 vssd1 vssd1 vccd1 vccd1
+ _0974_ sky130_fd_sc_hd__a21oi_1
X_1412_ outputs.divider_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__inv_2
X_2392_ net230 _0815_ _0798_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1274_ net1 net4 vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2728_ clknet_leaf_19_clk net163 net54 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2659_ clknet_leaf_22_clk _0005_ net36 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1892_ net257 _0334_ outputs.div.next_div _0395_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__a22o_1
X_1961_ outputs.scaled_buffer\[2\] net160 _1001_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2513_ _0876_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
X_1326_ _0963_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[10\]
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2444_ _0849_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__clkbuf_1
X_2375_ _0754_ _0756_ _1207_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__mux2_1
X_1257_ _0920_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2160_ _0531_ _0536_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__and3_1
X_2091_ _0525_ _0515_ _0523_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1944_ outputs.div.count\[1\] outputs.div.count\[0\] vssd1 vssd1 vccd1 vccd1 _0420_
+ sky130_fd_sc_hd__nand2_1
X_1875_ _0359_ _0374_ _0370_ _0378_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2427_ net309 net297 _0839_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1309_ _0940_ _0941_ _0951_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2289_ _1224_ _0718_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a21oi_1
X_2358_ _0464_ _0780_ _0784_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold209 outputs.div.q\[7\] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _1226_ _1233_ _1232_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__o21ba_1
X_1591_ outputs.scaled_buffer\[2\] _1161_ _1165_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _0465_ _0473_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__or2b_1
X_2212_ _0616_ _0480_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2074_ inputs.key_encoder.sync_keys\[4\] _0511_ inputs.key_encoder.sync_keys\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__o21ba_1
X_1927_ outputs.div.oscillator_out\[11\] _0411_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__and2_1
X_1858_ _0365_ _0366_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1789_ outputs.div.m\[14\] _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold81 outputs.div.q\[17\] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 _0141_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 outputs.div.q_out\[1\] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ clknet_leaf_9_clk _0148_ net46 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2692_ clknet_leaf_12_clk _0038_ net52 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2761_ clknet_leaf_1_clk _0079_ net27 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_1712_ _0229_ _0234_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__nand2_1
X_1643_ _1212_ _1208_ _1213_ _1222_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1574_ _1099_ net21 outputs.scaled_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__a21oi_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ _0466_ _0472_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__nand2_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2126_ _0559_ _0563_ _1215_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__mux2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1290_ inputs.random_update_clock.count\[1\] inputs.random_update_clock.count\[0\]
+ inputs.random_update_clock.count\[2\] vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2813_ clknet_leaf_2_clk _0131_ net41 vssd1 vssd1 vccd1 vccd1 outputs.signal_buffer2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2675_ clknet_leaf_17_clk _0021_ net55 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_2744_ clknet_leaf_3_clk outputs.sig_gen.next_count\[3\] net40 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1626_ _1206_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1488_ _1080_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
X_1557_ _1037_ outputs.shaper.count\[6\] vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nand2_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2109_ _0529_ _0544_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2460_ net129 _0829_ _0408_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1273_ _0928_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[10\] sky130_fd_sc_hd__clkbuf_1
X_1342_ net206 _0972_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[16\]
+ sky130_fd_sc_hd__xor2_1
X_1411_ outputs.divider_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__inv_2
X_2391_ _1208_ _0464_ _0761_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2727_ clknet_leaf_19_clk net175 net54 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2658_ clknet_leaf_23_clk _0004_ net36 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1609_ net21 _1163_ outputs.scaled_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2589_ clknet_leaf_35_clk net74 net22 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1891_ _0387_ _0391_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1960_ _0430_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2512_ outputs.shaper.count\[2\] net110 _0872_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__mux2_1
X_2443_ net310 outputs.div.m\[14\] _0839_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1325_ _0955_ _0961_ _0962_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__and3_1
X_2374_ _0799_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
X_1256_ _0917_ net11 vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2090_ _0521_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__or2_2
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1943_ _0419_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
X_1874_ _0377_ _0379_ _0380_ _0333_ net188 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2426_ _0840_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1308_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1239_ outputs.sample_rate.count\[1\] outputs.sample_rate.count\[0\] outputs.sample_rate.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__and3_1
X_2288_ _1206_ _0630_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__and2_1
X_2357_ _1207_ _0718_ _0783_ _0572_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] net21 _1158_ vssd1 vssd1
+ vccd1 vccd1 _1172_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _0645_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__clkbuf_1
X_2142_ _0466_ _0488_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nor2_4
X_2073_ inputs.key_encoder.sync_keys\[1\] _0510_ inputs.key_encoder.sync_keys\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1857_ outputs.div.a\[20\] _0342_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or2_1
X_1788_ outputs.div.m\[13\] outputs.div.m\[12\] _0285_ _0248_ vssd1 vssd1 vccd1 vccd1
+ _0304_ sky130_fd_sc_hd__o31a_1
X_1926_ _0994_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2409_ inputs.octave_fsm.state\[2\] _0754_ _1205_ vssd1 vssd1 vccd1 vccd1 _0830_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_79_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold82 _0047_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 _0070_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 outputs.div.divisor\[17\] vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold71 outputs.sample_rate.count\[0\] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_1
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2691_ clknet_leaf_12_clk _0037_ net52 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2760_ clknet_leaf_31_clk _0078_ net28 vssd1 vssd1 vccd1 vccd1 outputs.div.m\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_1711_ _0229_ _0234_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__or2_1
X_1642_ _1219_ _1221_ _1210_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1573_ _1142_ _1148_ _1149_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o211ai_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2056_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__clkbuf_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2125_ _0558_ _0560_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__or3_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1909_ outputs.div.oscillator_out\[3\] _0398_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2812_ clknet_leaf_11_clk _0130_ net42 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2743_ clknet_leaf_3_clk outputs.sig_gen.next_count\[2\] net39 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2674_ clknet_leaf_19_clk _0020_ net55 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1556_ _1030_ outputs.shaper.count\[5\] vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1625_ inputs.octave_fsm.state\[2\] _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__nand2_1
X_1487_ _1041_ _1078_ _1079_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__and3_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2039_ _0465_ _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nor2_4
X_2108_ _0525_ _0521_ _0530_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1410_ _1005_ _1009_ _1013_ _1015_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1272_ net1 net3 vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__and2b_1
X_1341_ _0972_ _0973_ vssd1 vssd1 vccd1 vccd1 inputs.random_update_clock.next_count\[15\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2390_ _0658_ _0812_ _0813_ _0789_ _0533_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2726_ clknet_leaf_18_clk net171 net54 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1539_ _1100_ _1106_ _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__or3_1
X_2657_ clknet_leaf_20_clk _0003_ net53 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1608_ outputs.output_gen.count\[5\] _1167_ _1189_ outputs.output_gen.count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2588_ clknet_leaf_35_clk net91 net22 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 outputs.div.q\[3\] vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1890_ outputs.div.m\[17\] outputs.div.a\[25\] _0336_ _0383_ _0389_ vssd1 vssd1 vccd1
+ vccd1 _0394_ sky130_fd_sc_hd__o311a_1
XFILLER_0_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2511_ _0875_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
X_2442_ _0848_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
X_2373_ net256 _0797_ _0798_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1324_ inputs.random_update_clock.count\[10\] _0959_ vssd1 vssd1 vccd1 vccd1 _0962_
+ sky130_fd_sc_hd__or2_1
X_1255_ _0919_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2709_ clknet_leaf_20_clk net217 net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1942_ _0996_ _0915_ outputs.div.count\[0\] vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1873_ _0372_ _0375_ _0378_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand3_1
XFILLER_0_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2425_ outputs.divider_buffer\[5\] outputs.div.m\[5\] _0839_ vssd1 vssd1 vccd1 vccd1
+ _0840_ sky130_fd_sc_hd__mux2_1
X_2356_ _1207_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__nor2_1
X_1307_ _0944_ _0947_ _0948_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2287_ _0682_ _0717_ _0554_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ net240 _0644_ _0606_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2072_ inputs.key_encoder.sync_keys\[2\] vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__inv_2
X_2141_ _0477_ _0576_ _0577_ _0468_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1925_ outputs.div.q\[18\] _0400_ _0405_ net143 _0410_ vssd1 vssd1 vccd1 vccd1 _0047_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1856_ outputs.div.a\[20\] _0355_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__nand2_1
X_1787_ outputs.div.a\[13\] vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2408_ _0910_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__clkbuf_4
X_2339_ _0615_ _0764_ _0765_ _0766_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold50 outputs.signal_buffer2\[11\] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 outputs.signal_buffer2\[5\] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 inputs.keypad_synchronizer.half_sync\[15\] vssd1 vssd1 vccd1 vccd1 net134
+ sky130_fd_sc_hd__buf_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 outputs.sample_rate.count\[2\] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 outputs.sample_rate.count\[4\] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1572_ _1130_ _1121_ _1150_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__or4b_1
X_2690_ clknet_leaf_19_clk net263 net53 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1710_ _0201_ _0207_ _0231_ _0220_ _0233_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__o41a_1
X_1641_ _1205_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _0524_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__nand2_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ _0465_ _0470_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__or2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1839_ net266 _0334_ outputs.div.next_div _0350_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__a22o_1
X_1908_ net183 _0400_ _0377_ net189 _0401_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2811_ clknet_leaf_11_clk _0129_ net52 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_2742_ clknet_leaf_3_clk outputs.sig_gen.next_count\[1\] net39 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2673_ clknet_leaf_20_clk _0019_ net51 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1555_ _1133_ _1134_ _1135_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__a31o_1
X_1624_ inputs.octave_fsm.state\[1\] inputs.octave_fsm.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _1205_ sky130_fd_sc_hd__nor2_1
X_1486_ outputs.sig_gen.count\[13\] _1075_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2107_ _0531_ _0544_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2038_ _0468_ inputs.frequency_lut.rng\[1\] vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1340_ net227 _0970_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1271_ _0927_ vssd1 vssd1 vccd1 vccd1 inputs.keypad\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2725_ clknet_leaf_18_clk net161 net54 vssd1 vssd1 vccd1 vccd1 outputs.div.q_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2656_ clknet_leaf_24_clk outputs.output_gen.pwm_unff net34 vssd1 vssd1 vccd1 vccd1
+ outputs.output_gen.pwm_ff sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1538_ _1109_ _1111_ _1114_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__or4_1
X_1469_ _1066_ vssd1 vssd1 vccd1 vccd1 outputs.sig_gen.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_1607_ outputs.scaled_buffer\[6\] _1161_ _1188_ _1157_ _1165_ vssd1 vssd1 vccd1 vccd1
+ _1189_ sky130_fd_sc_hd__a221oi_1
X_2587_ clknet_leaf_35_clk net88 net24 vssd1 vssd1 vccd1 vccd1 inputs.random_note_generator.out\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold180 _0985_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _0033_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2510_ net300 net125 _0872_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1323_ inputs.random_update_clock.count\[10\] _0959_ vssd1 vssd1 vccd1 vccd1 _0961_
+ sky130_fd_sc_hd__nand2_1
X_2441_ outputs.divider_buffer\[13\] outputs.div.m\[13\] _0839_ vssd1 vssd1 vccd1
+ vccd1 _0848_ sky130_fd_sc_hd__mux2_1
X_2372_ _0994_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1254_ _0917_ net10 vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2639_ clknet_leaf_15_clk inputs.keypad\[0\] net60 vssd1 vssd1 vccd1 vccd1 inputs.keypad_synchronizer.half_sync\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2708_ clknet_leaf_13_clk net205 net57 vssd1 vssd1 vccd1 vccd1 outputs.div.q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1872_ _0372_ _0375_ _0378_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__a21o_1
X_1941_ net216 _1228_ _1225_ outputs.div.q\[25\] vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1306_ inputs.random_update_clock.count\[20\] inputs.random_update_clock.count\[22\]
+ inputs.random_update_clock.count\[21\] vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__nor3b_1
X_2424_ _0994_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__clkbuf_4
X_2286_ _1215_ _0715_ _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__o21ai_1
X_2355_ _0554_ _0755_ _0781_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2140_ _0481_ _0474_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2071_ _0483_ _0490_ _0501_ _0504_ _0506_ _0508_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__mux4_1
X_1924_ outputs.div.oscillator_out\[10\] _0398_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__and2_1
X_1855_ _0205_ _0363_ _0364_ _0333_ net236 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1786_ net224 _0916_ outputs.div.next_div _0302_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2407_ _0828_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_1
X_2338_ _0491_ _0730_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__nor2_1
X_2269_ _0506_ _0696_ _0698_ _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold40 _0137_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold51 _0142_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 outputs.signal_buffer2\[15\] vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0136_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _0997_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 inputs.key_encoder.sync_keys\[15\] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1571_ _1135_ _1138_ _1151_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__and4_1
X_1640_ inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _0515_ _0528_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__or2_1
X_2054_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1838_ _0345_ _0349_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__xor2_1
X_1907_ net315 _0398_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1769_ outputs.div.m\[12\] _0286_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2810_ clknet_leaf_11_clk _0128_ net42 vssd1 vssd1 vccd1 vccd1 outputs.divider_buffer\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_2672_ clknet_leaf_19_clk _0018_ net53 vssd1 vssd1 vccd1 vccd1 outputs.div.a\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2741_ clknet_leaf_3_clk outputs.sig_gen.next_count\[0\] net39 vssd1 vssd1 vccd1
+ vccd1 outputs.sig_gen.count\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1485_ outputs.sig_gen.count\[13\] _1075_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__or2_1
X_1554_ _1030_ outputs.shaper.count\[5\] outputs.shaper.count\[4\] _1019_ vssd1 vssd1
+ vccd1 vccd1 _1136_ sky130_fd_sc_hd__o22ai_2
X_1623_ _1204_ vssd1 vssd1 vccd1 vccd1 outputs.output_gen.pwm_unff sky130_fd_sc_hd__clkbuf_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

