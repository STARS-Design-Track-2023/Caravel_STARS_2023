magic
tech sky130A
magscale 1 2
timestamp 1693854964
<< obsli1 >>
rect 1104 2159 72404 73457
<< obsm1 >>
rect 14 2048 72574 73488
<< metal2 >>
rect 4526 74901 4582 75701
rect 10322 74901 10378 75701
rect 16118 74901 16174 75701
rect 21270 74901 21326 75701
rect 27066 74901 27122 75701
rect 32218 74901 32274 75701
rect 38014 74901 38070 75701
rect 43166 74901 43222 75701
rect 48962 74901 49018 75701
rect 54758 74901 54814 75701
rect 59910 74901 59966 75701
rect 65706 74901 65762 75701
rect 70858 74901 70914 75701
rect 18 0 74 800
rect 5170 0 5226 800
rect 10966 0 11022 800
rect 16118 0 16174 800
rect 21914 0 21970 800
rect 27066 0 27122 800
rect 32862 0 32918 800
rect 38014 0 38070 800
rect 43810 0 43866 800
rect 49606 0 49662 800
rect 54758 0 54814 800
rect 60554 0 60610 800
rect 65706 0 65762 800
rect 71502 0 71558 800
<< obsm2 >>
rect 20 74845 4470 75449
rect 4638 74845 10266 75449
rect 10434 74845 16062 75449
rect 16230 74845 21214 75449
rect 21382 74845 27010 75449
rect 27178 74845 32162 75449
rect 32330 74845 37958 75449
rect 38126 74845 43110 75449
rect 43278 74845 48906 75449
rect 49074 74845 54702 75449
rect 54870 74845 59854 75449
rect 60022 74845 65650 75449
rect 65818 74845 70802 75449
rect 70970 74845 72570 75449
rect 20 856 72570 74845
rect 130 734 5114 856
rect 5282 734 10910 856
rect 11078 734 16062 856
rect 16230 734 21858 856
rect 22026 734 27010 856
rect 27178 734 32806 856
rect 32974 734 37958 856
rect 38126 734 43754 856
rect 43922 734 49550 856
rect 49718 734 54702 856
rect 54870 734 60498 856
rect 60666 734 65650 856
rect 65818 734 71446 856
rect 71614 734 72570 856
<< metal3 >>
rect 0 75488 800 75608
rect 72757 72768 73557 72888
rect 0 69368 800 69488
rect 72757 67328 73557 67448
rect 0 63928 800 64048
rect 72757 61208 73557 61328
rect 0 57808 800 57928
rect 72757 55768 73557 55888
rect 0 52368 800 52488
rect 72757 49648 73557 49768
rect 0 46248 800 46368
rect 72757 43528 73557 43648
rect 0 40128 800 40248
rect 72757 38088 73557 38208
rect 0 34688 800 34808
rect 72757 31968 73557 32088
rect 0 28568 800 28688
rect 72757 26528 73557 26648
rect 0 23128 800 23248
rect 72757 20408 73557 20528
rect 0 17008 800 17128
rect 72757 14968 73557 15088
rect 0 11568 800 11688
rect 72757 8848 73557 8968
rect 0 5448 800 5568
rect 72757 2728 73557 2848
<< obsm3 >>
rect 880 75408 72757 75578
rect 798 72968 72757 75408
rect 798 72688 72677 72968
rect 798 69568 72757 72688
rect 880 69288 72757 69568
rect 798 67528 72757 69288
rect 798 67248 72677 67528
rect 798 64128 72757 67248
rect 880 63848 72757 64128
rect 798 61408 72757 63848
rect 798 61128 72677 61408
rect 798 58008 72757 61128
rect 880 57728 72757 58008
rect 798 55968 72757 57728
rect 798 55688 72677 55968
rect 798 52568 72757 55688
rect 880 52288 72757 52568
rect 798 49848 72757 52288
rect 798 49568 72677 49848
rect 798 46448 72757 49568
rect 880 46168 72757 46448
rect 798 43728 72757 46168
rect 798 43448 72677 43728
rect 798 40328 72757 43448
rect 880 40048 72757 40328
rect 798 38288 72757 40048
rect 798 38008 72677 38288
rect 798 34888 72757 38008
rect 880 34608 72757 34888
rect 798 32168 72757 34608
rect 798 31888 72677 32168
rect 798 28768 72757 31888
rect 880 28488 72757 28768
rect 798 26728 72757 28488
rect 798 26448 72677 26728
rect 798 23328 72757 26448
rect 880 23048 72757 23328
rect 798 20608 72757 23048
rect 798 20328 72677 20608
rect 798 17208 72757 20328
rect 880 16928 72757 17208
rect 798 15168 72757 16928
rect 798 14888 72677 15168
rect 798 11768 72757 14888
rect 880 11488 72757 11768
rect 798 9048 72757 11488
rect 798 8768 72677 9048
rect 798 5648 72757 8768
rect 880 5368 72757 5648
rect 798 2928 72757 5368
rect 798 2648 72677 2928
rect 798 2143 72757 2648
<< metal4 >>
rect 4208 2128 4528 73488
rect 19568 2128 19888 73488
rect 34928 2128 35248 73488
rect 50288 2128 50608 73488
rect 65648 2128 65968 73488
<< obsm4 >>
rect 15515 10235 19488 71909
rect 19968 10235 34848 71909
rect 35328 10235 50208 71909
rect 50688 10235 59373 71909
<< obsm5 >>
rect 19068 32140 45700 35180
<< labels >>
rlabel metal4 s 19568 2128 19888 73488 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 73488 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 73488 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 73488 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 73488 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 16118 0 16174 800 6 beat_led[0]
port 3 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 beat_led[1]
port 4 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 beat_led[2]
port 5 nsew signal output
rlabel metal2 s 4526 74901 4582 75701 6 beat_led[3]
port 6 nsew signal output
rlabel metal3 s 72757 38088 73557 38208 6 beat_led[4]
port 7 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 beat_led[5]
port 8 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 beat_led[6]
port 9 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 beat_led[7]
port 10 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 cs
port 11 nsew signal input
rlabel metal3 s 72757 8848 73557 8968 6 hwclk
port 12 nsew signal input
rlabel metal2 s 48962 74901 49018 75701 6 mode_out[0]
port 13 nsew signal output
rlabel metal3 s 72757 2728 73557 2848 6 mode_out[1]
port 14 nsew signal output
rlabel metal2 s 59910 74901 59966 75701 6 multi[0]
port 15 nsew signal output
rlabel metal3 s 72757 14968 73557 15088 6 multi[1]
port 16 nsew signal output
rlabel metal2 s 10322 74901 10378 75701 6 multi[2]
port 17 nsew signal output
rlabel metal3 s 72757 20408 73557 20528 6 multi[3]
port 18 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 n_rst
port 19 nsew signal input
rlabel metal3 s 72757 67328 73557 67448 6 note1[0]
port 20 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 note1[1]
port 21 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 note1[2]
port 22 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 note1[3]
port 23 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 note2[0]
port 24 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 note2[1]
port 25 nsew signal output
rlabel metal3 s 72757 55768 73557 55888 6 note2[2]
port 26 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 note2[3]
port 27 nsew signal output
rlabel metal2 s 43166 74901 43222 75701 6 note3[0]
port 28 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 note3[1]
port 29 nsew signal output
rlabel metal3 s 72757 72768 73557 72888 6 note3[2]
port 30 nsew signal output
rlabel metal2 s 32218 74901 32274 75701 6 note3[3]
port 31 nsew signal output
rlabel metal3 s 72757 43528 73557 43648 6 note4[0]
port 32 nsew signal output
rlabel metal2 s 54758 74901 54814 75701 6 note4[1]
port 33 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 note4[2]
port 34 nsew signal output
rlabel metal2 s 18 0 74 800 6 note4[3]
port 35 nsew signal output
rlabel metal2 s 21270 74901 21326 75701 6 piano_keys[0]
port 36 nsew signal input
rlabel metal3 s 72757 61208 73557 61328 6 piano_keys[10]
port 37 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 piano_keys[11]
port 38 nsew signal input
rlabel metal3 s 72757 49648 73557 49768 6 piano_keys[12]
port 39 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 piano_keys[13]
port 40 nsew signal input
rlabel metal2 s 38014 74901 38070 75701 6 piano_keys[14]
port 41 nsew signal input
rlabel metal3 s 72757 26528 73557 26648 6 piano_keys[1]
port 42 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 piano_keys[2]
port 43 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 piano_keys[3]
port 44 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 piano_keys[4]
port 45 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 piano_keys[5]
port 46 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 piano_keys[6]
port 47 nsew signal input
rlabel metal2 s 70858 74901 70914 75701 6 piano_keys[7]
port 48 nsew signal input
rlabel metal2 s 65706 74901 65762 75701 6 piano_keys[8]
port 49 nsew signal input
rlabel metal2 s 16118 74901 16174 75701 6 piano_keys[9]
port 50 nsew signal input
rlabel metal2 s 27066 74901 27122 75701 6 pwm_o
port 51 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 seq_led_on
port 52 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 seq_play
port 53 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 seq_power
port 54 nsew signal input
rlabel metal3 s 72757 31968 73557 32088 6 tempo_select
port 55 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 73557 75701
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13720450
string GDS_FILE /home/designer-25/CUP/openlane/SaSS/runs/23_09_04_12_07/results/signoff/sass_synth.magic.gds
string GDS_START 1144644
<< end >>

