magic
tech sky130A
magscale 1 2
timestamp 1691545472
<< obsli1 >>
rect 1104 2159 38272 39185
<< obsm1 >>
rect 14 2128 38350 39216
<< metal2 >>
rect 662 40765 718 41565
rect 2594 40765 2650 41565
rect 5170 40765 5226 41565
rect 7102 40765 7158 41565
rect 9678 40765 9734 41565
rect 11610 40765 11666 41565
rect 14186 40765 14242 41565
rect 16118 40765 16174 41565
rect 18694 40765 18750 41565
rect 20626 40765 20682 41565
rect 23202 40765 23258 41565
rect 25134 40765 25190 41565
rect 27066 40765 27122 41565
rect 29642 40765 29698 41565
rect 31574 40765 31630 41565
rect 34150 40765 34206 41565
rect 36082 40765 36138 41565
rect 38658 40765 38714 41565
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 15474 0 15530 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 21914 0 21970 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28998 0 29054 800
rect 30930 0 30986 800
rect 32862 0 32918 800
rect 35438 0 35494 800
rect 37370 0 37426 800
<< obsm2 >>
rect 20 40709 606 40882
rect 774 40709 2538 40882
rect 2706 40709 5114 40882
rect 5282 40709 7046 40882
rect 7214 40709 9622 40882
rect 9790 40709 11554 40882
rect 11722 40709 14130 40882
rect 14298 40709 16062 40882
rect 16230 40709 18638 40882
rect 18806 40709 20570 40882
rect 20738 40709 23146 40882
rect 23314 40709 25078 40882
rect 25246 40709 27010 40882
rect 27178 40709 29586 40882
rect 29754 40709 31518 40882
rect 31686 40709 34094 40882
rect 34262 40709 36026 40882
rect 36194 40709 38346 40882
rect 20 856 38346 40709
rect 130 31 1894 856
rect 2062 31 3826 856
rect 3994 31 6402 856
rect 6570 31 8334 856
rect 8502 31 10910 856
rect 11078 31 12842 856
rect 13010 31 15418 856
rect 15586 31 17350 856
rect 17518 31 19926 856
rect 20094 31 21858 856
rect 22026 31 24434 856
rect 24602 31 26366 856
rect 26534 31 28942 856
rect 29110 31 30874 856
rect 31042 31 32806 856
rect 32974 31 35382 856
rect 35550 31 37314 856
rect 37482 31 38346 856
<< metal3 >>
rect 38621 40128 39421 40248
rect 0 39448 800 39568
rect 0 37408 800 37528
rect 38621 37408 39421 37528
rect 38621 35368 39421 35488
rect 0 34688 800 34808
rect 0 32648 800 32768
rect 38621 32648 39421 32768
rect 0 30608 800 30728
rect 38621 30608 39421 30728
rect 0 27888 800 28008
rect 38621 27888 39421 28008
rect 0 25848 800 25968
rect 38621 25848 39421 25968
rect 38621 23808 39421 23928
rect 0 23128 800 23248
rect 0 21088 800 21208
rect 38621 21088 39421 21208
rect 38621 19048 39421 19168
rect 0 18368 800 18488
rect 0 16328 800 16448
rect 38621 16328 39421 16448
rect 38621 14288 39421 14408
rect 0 13608 800 13728
rect 0 11568 800 11688
rect 38621 11568 39421 11688
rect 38621 9528 39421 9648
rect 0 8848 800 8968
rect 0 6808 800 6928
rect 38621 6808 39421 6928
rect 38621 4768 39421 4888
rect 0 4088 800 4208
rect 0 2048 800 2168
rect 38621 2048 39421 2168
rect 38621 8 39421 128
<< obsm3 >>
rect 800 40048 38541 40221
rect 800 39648 38621 40048
rect 880 39368 38621 39648
rect 800 37608 38621 39368
rect 880 37328 38541 37608
rect 800 35568 38621 37328
rect 800 35288 38541 35568
rect 800 34888 38621 35288
rect 880 34608 38621 34888
rect 800 32848 38621 34608
rect 880 32568 38541 32848
rect 800 30808 38621 32568
rect 880 30528 38541 30808
rect 800 28088 38621 30528
rect 880 27808 38541 28088
rect 800 26048 38621 27808
rect 880 25768 38541 26048
rect 800 24008 38621 25768
rect 800 23728 38541 24008
rect 800 23328 38621 23728
rect 880 23048 38621 23328
rect 800 21288 38621 23048
rect 880 21008 38541 21288
rect 800 19248 38621 21008
rect 800 18968 38541 19248
rect 800 18568 38621 18968
rect 880 18288 38621 18568
rect 800 16528 38621 18288
rect 880 16248 38541 16528
rect 800 14488 38621 16248
rect 800 14208 38541 14488
rect 800 13808 38621 14208
rect 880 13528 38621 13808
rect 800 11768 38621 13528
rect 880 11488 38541 11768
rect 800 9728 38621 11488
rect 800 9448 38541 9728
rect 800 9048 38621 9448
rect 880 8768 38621 9048
rect 800 7008 38621 8768
rect 880 6728 38541 7008
rect 800 4968 38621 6728
rect 800 4688 38541 4968
rect 800 4288 38621 4688
rect 880 4008 38621 4288
rect 800 2248 38621 4008
rect 880 1968 38541 2248
rect 800 208 38621 1968
rect 800 35 38541 208
<< metal4 >>
rect 4208 2128 4528 39216
rect 4868 2128 5188 39216
rect 34928 2128 35248 39216
rect 35588 2128 35908 39216
<< obsm4 >>
rect 11467 2347 31037 35869
<< metal5 >>
rect 1056 36642 38320 36962
rect 1056 35982 38320 36302
rect 1056 6006 38320 6326
rect 1056 5346 38320 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 39216 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 39216 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 38320 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 38320 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 39216 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 39216 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 38320 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 38320 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 2594 40765 2650 41565 6 clk
port 3 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 cs
port 4 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 gpi[0]
port 5 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 gpi[10]
port 6 nsew signal input
rlabel metal3 s 38621 23808 39421 23928 6 gpi[11]
port 7 nsew signal input
rlabel metal2 s 16118 40765 16174 41565 6 gpi[12]
port 8 nsew signal input
rlabel metal2 s 38658 40765 38714 41565 6 gpi[13]
port 9 nsew signal input
rlabel metal3 s 38621 27888 39421 28008 6 gpi[14]
port 10 nsew signal input
rlabel metal3 s 38621 6808 39421 6928 6 gpi[15]
port 11 nsew signal input
rlabel metal3 s 38621 25848 39421 25968 6 gpi[16]
port 12 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 gpi[17]
port 13 nsew signal input
rlabel metal3 s 38621 9528 39421 9648 6 gpi[18]
port 14 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 gpi[19]
port 15 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 gpi[1]
port 16 nsew signal input
rlabel metal3 s 38621 4768 39421 4888 6 gpi[20]
port 17 nsew signal input
rlabel metal2 s 11610 40765 11666 41565 6 gpi[21]
port 18 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 gpi[22]
port 19 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 gpi[23]
port 20 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 gpi[24]
port 21 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 gpi[25]
port 22 nsew signal input
rlabel metal3 s 38621 30608 39421 30728 6 gpi[26]
port 23 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 gpi[27]
port 24 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 gpi[28]
port 25 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 gpi[29]
port 26 nsew signal input
rlabel metal3 s 38621 32648 39421 32768 6 gpi[2]
port 27 nsew signal input
rlabel metal3 s 38621 16328 39421 16448 6 gpi[30]
port 28 nsew signal input
rlabel metal2 s 29642 40765 29698 41565 6 gpi[31]
port 29 nsew signal input
rlabel metal2 s 7102 40765 7158 41565 6 gpi[32]
port 30 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 gpi[33]
port 31 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 gpi[3]
port 32 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 gpi[4]
port 33 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 gpi[5]
port 34 nsew signal input
rlabel metal2 s 20626 40765 20682 41565 6 gpi[6]
port 35 nsew signal input
rlabel metal3 s 38621 40128 39421 40248 6 gpi[7]
port 36 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 gpi[8]
port 37 nsew signal input
rlabel metal2 s 18694 40765 18750 41565 6 gpi[9]
port 38 nsew signal input
rlabel metal3 s 38621 2048 39421 2168 6 gpo[0]
port 39 nsew signal output
rlabel metal3 s 38621 11568 39421 11688 6 gpo[10]
port 40 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 gpo[11]
port 41 nsew signal output
rlabel metal3 s 38621 14288 39421 14408 6 gpo[12]
port 42 nsew signal output
rlabel metal2 s 25134 40765 25190 41565 6 gpo[13]
port 43 nsew signal output
rlabel metal2 s 27066 40765 27122 41565 6 gpo[14]
port 44 nsew signal output
rlabel metal2 s 662 40765 718 41565 6 gpo[15]
port 45 nsew signal output
rlabel metal2 s 18 0 74 800 6 gpo[16]
port 46 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 gpo[17]
port 47 nsew signal output
rlabel metal2 s 23202 40765 23258 41565 6 gpo[18]
port 48 nsew signal output
rlabel metal2 s 31574 40765 31630 41565 6 gpo[19]
port 49 nsew signal output
rlabel metal3 s 38621 37408 39421 37528 6 gpo[1]
port 50 nsew signal output
rlabel metal2 s 14186 40765 14242 41565 6 gpo[20]
port 51 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 gpo[21]
port 52 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 gpo[22]
port 53 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 gpo[23]
port 54 nsew signal output
rlabel metal2 s 36082 40765 36138 41565 6 gpo[24]
port 55 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 gpo[25]
port 56 nsew signal output
rlabel metal3 s 38621 35368 39421 35488 6 gpo[26]
port 57 nsew signal output
rlabel metal3 s 38621 8 39421 128 6 gpo[27]
port 58 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 gpo[28]
port 59 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 gpo[29]
port 60 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 gpo[2]
port 61 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 gpo[30]
port 62 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 gpo[31]
port 63 nsew signal output
rlabel metal3 s 38621 21088 39421 21208 6 gpo[32]
port 64 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 gpo[33]
port 65 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 gpo[3]
port 66 nsew signal output
rlabel metal2 s 34150 40765 34206 41565 6 gpo[4]
port 67 nsew signal output
rlabel metal2 s 5170 40765 5226 41565 6 gpo[5]
port 68 nsew signal output
rlabel metal2 s 9678 40765 9734 41565 6 gpo[6]
port 69 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 gpo[7]
port 70 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 gpo[8]
port 71 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 gpo[9]
port 72 nsew signal output
rlabel metal3 s 38621 19048 39421 19168 6 nrst
port 73 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 39421 41565
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5070438
string GDS_FILE /home/designer-25/CUP/openlane/Eighty_Twos/runs/23_08_08_18_39/results/signoff/Eighty_Twos.magic.gds
string GDS_START 1047140
<< end >>

