VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pushing_pixels
  CLASS BLOCK ;
  FOREIGN pushing_pixels ;
  ORIGIN 0.000 0.000 ;
  SIZE 1376.390 BY 1387.110 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1375.030 1383.110 1375.310 1387.110 ;
    END
  END clk
  PIN color[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END color[0]
  PIN color[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END color[10]
  PIN color[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END color[11]
  PIN color[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 367.170 1383.110 367.450 1387.110 ;
    END
  END color[12]
  PIN color[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 872.710 1383.110 872.990 1387.110 ;
    END
  END color[13]
  PIN color[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END color[14]
  PIN color[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1372.390 676.640 1376.390 677.240 ;
    END
  END color[15]
  PIN color[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END color[16]
  PIN color[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1372.390 853.440 1376.390 854.040 ;
    END
  END color[17]
  PIN color[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END color[18]
  PIN color[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END color[19]
  PIN color[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1383.110 1040.430 1387.110 ;
    END
  END color[1]
  PIN color[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1207.590 1383.110 1207.870 1387.110 ;
    END
  END color[20]
  PIN color[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END color[21]
  PIN color[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1372.390 142.840 1376.390 143.440 ;
    END
  END color[22]
  PIN color[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END color[23]
  PIN color[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.040 4.000 1241.640 ;
    END
  END color[2]
  PIN color[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END color[3]
  PIN color[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END color[4]
  PIN color[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END color[5]
  PIN color[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 199.730 1383.110 200.010 1387.110 ;
    END
  END color[6]
  PIN color[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1372.390 319.640 1376.390 320.240 ;
    END
  END color[7]
  PIN color[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END color[8]
  PIN color[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1372.390 1030.240 1376.390 1030.840 ;
    END
  END color[9]
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1372.390 1207.040 1376.390 1207.640 ;
    END
  END cs
  PIN is_mandelbrot
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 534.610 1383.110 534.890 1387.110 ;
    END
  END is_mandelbrot
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 702.050 1383.110 702.330 1387.110 ;
    END
  END nrst
  PIN spi_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END spi_clk
  PIN spi_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END spi_data
  PIN spi_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 1383.110 29.350 1387.110 ;
    END
  END spi_en
  PIN valid_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1372.390 496.440 1376.390 497.040 ;
    END
  END valid_out
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1373.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1373.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1373.840 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1370.800 1373.685 ;
      LAYER met1 ;
        RECT 0.070 10.640 1375.330 1373.840 ;
      LAYER met2 ;
        RECT 0.100 1382.830 28.790 1383.110 ;
        RECT 29.630 1382.830 199.450 1383.110 ;
        RECT 200.290 1382.830 366.890 1383.110 ;
        RECT 367.730 1382.830 534.330 1383.110 ;
        RECT 535.170 1382.830 701.770 1383.110 ;
        RECT 702.610 1382.830 872.430 1383.110 ;
        RECT 873.270 1382.830 1039.870 1383.110 ;
        RECT 1040.710 1382.830 1207.310 1383.110 ;
        RECT 1208.150 1382.830 1374.750 1383.110 ;
        RECT 0.100 4.280 1375.300 1382.830 ;
        RECT 0.650 3.670 167.250 4.280 ;
        RECT 168.090 3.670 334.690 4.280 ;
        RECT 335.530 3.670 502.130 4.280 ;
        RECT 502.970 3.670 672.790 4.280 ;
        RECT 673.630 3.670 840.230 4.280 ;
        RECT 841.070 3.670 1007.670 4.280 ;
        RECT 1008.510 3.670 1175.110 4.280 ;
        RECT 1175.950 3.670 1345.770 4.280 ;
        RECT 1346.610 3.670 1375.300 4.280 ;
      LAYER met3 ;
        RECT 4.000 1242.040 1372.390 1373.765 ;
        RECT 4.400 1240.640 1372.390 1242.040 ;
        RECT 4.000 1208.040 1372.390 1240.640 ;
        RECT 4.000 1206.640 1371.990 1208.040 ;
        RECT 4.000 1065.240 1372.390 1206.640 ;
        RECT 4.400 1063.840 1372.390 1065.240 ;
        RECT 4.000 1031.240 1372.390 1063.840 ;
        RECT 4.000 1029.840 1371.990 1031.240 ;
        RECT 4.000 888.440 1372.390 1029.840 ;
        RECT 4.400 887.040 1372.390 888.440 ;
        RECT 4.000 854.440 1372.390 887.040 ;
        RECT 4.000 853.040 1371.990 854.440 ;
        RECT 4.000 708.240 1372.390 853.040 ;
        RECT 4.400 706.840 1372.390 708.240 ;
        RECT 4.000 677.640 1372.390 706.840 ;
        RECT 4.000 676.240 1371.990 677.640 ;
        RECT 4.000 531.440 1372.390 676.240 ;
        RECT 4.400 530.040 1372.390 531.440 ;
        RECT 4.000 497.440 1372.390 530.040 ;
        RECT 4.000 496.040 1371.990 497.440 ;
        RECT 4.000 354.640 1372.390 496.040 ;
        RECT 4.400 353.240 1372.390 354.640 ;
        RECT 4.000 320.640 1372.390 353.240 ;
        RECT 4.000 319.240 1371.990 320.640 ;
        RECT 4.000 177.840 1372.390 319.240 ;
        RECT 4.400 176.440 1372.390 177.840 ;
        RECT 4.000 143.840 1372.390 176.440 ;
        RECT 4.000 142.440 1371.990 143.840 ;
        RECT 4.000 10.715 1372.390 142.440 ;
      LAYER met4 ;
        RECT 313.095 11.735 327.840 1366.625 ;
        RECT 330.240 11.735 404.640 1366.625 ;
        RECT 407.040 11.735 481.440 1366.625 ;
        RECT 483.840 11.735 558.240 1366.625 ;
        RECT 560.640 11.735 635.040 1366.625 ;
        RECT 637.440 11.735 711.840 1366.625 ;
        RECT 714.240 11.735 788.640 1366.625 ;
        RECT 791.040 11.735 865.440 1366.625 ;
        RECT 867.840 11.735 942.240 1366.625 ;
        RECT 944.640 11.735 1019.040 1366.625 ;
        RECT 1021.440 11.735 1029.185 1366.625 ;
  END
END pushing_pixels
END LIBRARY

