// This is the unpowered netlist.
module outel8227 (clk,
    cs,
    dataBusSelect,
    nrst,
    dataBusIn,
    dataBusOut,
    gpio);
 input clk;
 input cs;
 output dataBusSelect;
 input nrst;
 input [7:0] dataBusIn;
 output [7:0] dataBusOut;
 inout [25:0] gpio;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire \top8227.PSRCurrentValue[0] ;
 wire \top8227.PSRCurrentValue[1] ;
 wire \top8227.PSRCurrentValue[2] ;
 wire \top8227.PSRCurrentValue[3] ;
 wire \top8227.PSRCurrentValue[6] ;
 wire \top8227.PSRCurrentValue[7] ;
 wire \top8227.branchBackward ;
 wire \top8227.branchForward ;
 wire \top8227.demux.isAddressing ;
 wire \top8227.demux.nmi ;
 wire \top8227.demux.reset ;
 wire \top8227.demux.setInterruptFlag ;
 wire \top8227.demux.state_machine.currentAddress[0] ;
 wire \top8227.demux.state_machine.currentAddress[10] ;
 wire \top8227.demux.state_machine.currentAddress[11] ;
 wire \top8227.demux.state_machine.currentAddress[12] ;
 wire \top8227.demux.state_machine.currentAddress[1] ;
 wire \top8227.demux.state_machine.currentAddress[2] ;
 wire \top8227.demux.state_machine.currentAddress[3] ;
 wire \top8227.demux.state_machine.currentAddress[4] ;
 wire \top8227.demux.state_machine.currentAddress[5] ;
 wire \top8227.demux.state_machine.currentAddress[6] ;
 wire \top8227.demux.state_machine.currentAddress[7] ;
 wire \top8227.demux.state_machine.currentAddress[8] ;
 wire \top8227.demux.state_machine.currentAddress[9] ;
 wire \top8227.demux.state_machine.currentInstruction[0] ;
 wire \top8227.demux.state_machine.currentInstruction[1] ;
 wire \top8227.demux.state_machine.currentInstruction[2] ;
 wire \top8227.demux.state_machine.currentInstruction[3] ;
 wire \top8227.demux.state_machine.currentInstruction[4] ;
 wire \top8227.demux.state_machine.currentInstruction[5] ;
 wire \top8227.demux.state_machine.timeState[0] ;
 wire \top8227.demux.state_machine.timeState[1] ;
 wire \top8227.demux.state_machine.timeState[2] ;
 wire \top8227.demux.state_machine.timeState[3] ;
 wire \top8227.demux.state_machine.timeState[4] ;
 wire \top8227.demux.state_machine.timeState[5] ;
 wire \top8227.demux.state_machine.timeState[6] ;
 wire \top8227.freeCarry ;
 wire \top8227.instructionLoader.interruptInjector.interruptRequest ;
 wire \top8227.instructionLoader.interruptInjector.irqGenerated ;
 wire \top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ ;
 wire \top8227.instructionLoader.interruptInjector.irqSync.nextQ2 ;
 wire \top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ;
 wire \top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI ;
 wire \top8227.instructionLoader.interruptInjector.nmiSync.in ;
 wire \top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 ;
 wire \top8227.instructionLoader.interruptInjector.resetDetected ;
 wire \top8227.internalDataflow.accRegToDB[0] ;
 wire \top8227.internalDataflow.accRegToDB[1] ;
 wire \top8227.internalDataflow.accRegToDB[2] ;
 wire \top8227.internalDataflow.accRegToDB[3] ;
 wire \top8227.internalDataflow.accRegToDB[4] ;
 wire \top8227.internalDataflow.accRegToDB[5] ;
 wire \top8227.internalDataflow.accRegToDB[6] ;
 wire \top8227.internalDataflow.accRegToDB[7] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[16] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[17] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[18] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[19] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[20] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[21] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[22] ;
 wire \top8227.internalDataflow.addressHighBusModule.busInputs[23] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[16] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[17] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[18] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[19] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[20] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[21] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[22] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[23] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[24] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[25] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[26] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[27] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[28] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[29] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[30] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[31] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[32] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[33] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[34] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[35] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[36] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[37] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[38] ;
 wire \top8227.internalDataflow.addressLowBusModule.busInputs[39] ;
 wire \top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[0] ;
 wire \top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[1] ;
 wire \top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[2] ;
 wire \top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[3] ;
 wire \top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[6] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[32] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[33] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[34] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[35] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[36] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[37] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[38] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[39] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[40] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[41] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[42] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[43] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[44] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[45] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[46] ;
 wire \top8227.internalDataflow.stackBusModule.busInputs[47] ;
 wire \top8227.negEdgeDetector.q1 ;
 wire \top8227.pulse_slower.currentEnableState[0] ;
 wire \top8227.pulse_slower.currentEnableState[1] ;
 wire \top8227.pulse_slower.nextEnableState[0] ;
 wire \top8227.pulse_slower.nextEnableState[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\top8227.PSRCurrentValue[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\top8227.PSRCurrentValue[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net18));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__clkbuf_4 _1509_ (.A(\top8227.demux.state_machine.timeState[2] ),
    .X(_0814_));
 sky130_fd_sc_hd__buf_2 _1510_ (.A(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _1511_ (.A(\top8227.branchBackward ),
    .B(\top8227.branchForward ),
    .Y(_0816_));
 sky130_fd_sc_hd__and2_1 _1512_ (.A(_0815_),
    .B(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _1513_ (.A(\top8227.demux.state_machine.timeState[4] ),
    .X(_0818_));
 sky130_fd_sc_hd__clkbuf_4 _1514_ (.A(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__buf_2 _1515_ (.A(\top8227.demux.state_machine.currentInstruction[3] ),
    .X(_0820_));
 sky130_fd_sc_hd__buf_2 _1516_ (.A(\top8227.demux.state_machine.currentInstruction[2] ),
    .X(_0821_));
 sky130_fd_sc_hd__or4b_1 _1517_ (.A(\top8227.demux.state_machine.currentInstruction[1] ),
    .B(\top8227.demux.state_machine.currentInstruction[0] ),
    .C(_0820_),
    .D_N(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_4 _1518_ (.A(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__or2_1 _1519_ (.A(\top8227.demux.state_machine.currentInstruction[5] ),
    .B(\top8227.demux.state_machine.currentInstruction[4] ),
    .X(_0824_));
 sky130_fd_sc_hd__clkbuf_4 _1520_ (.A(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__buf_2 _1521_ (.A(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__inv_2 _1522_ (.A(\top8227.PSRCurrentValue[0] ),
    .Y(_0827_));
 sky130_fd_sc_hd__clkbuf_2 _1523_ (.A(\top8227.demux.state_machine.currentInstruction[1] ),
    .X(_0828_));
 sky130_fd_sc_hd__or4bb_1 _1524_ (.A(_0828_),
    .B(_0820_),
    .C_N(_0821_),
    .D_N(\top8227.demux.state_machine.currentInstruction[0] ),
    .X(_0829_));
 sky130_fd_sc_hd__clkbuf_4 _1525_ (.A(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__or3_1 _1526_ (.A(_0827_),
    .B(_0830_),
    .C(_0826_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_4 _1527_ (.A(\top8227.demux.state_machine.currentInstruction[5] ),
    .X(_0832_));
 sky130_fd_sc_hd__or4b_1 _1528_ (.A(\top8227.demux.state_machine.currentInstruction[1] ),
    .B(\top8227.demux.state_machine.currentInstruction[0] ),
    .C(\top8227.demux.state_machine.currentInstruction[2] ),
    .D_N(\top8227.demux.state_machine.currentInstruction[3] ),
    .X(_0833_));
 sky130_fd_sc_hd__buf_4 _1529_ (.A(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_4 _1530_ (.A(\top8227.demux.state_machine.currentInstruction[4] ),
    .X(_0835_));
 sky130_fd_sc_hd__or4b_1 _1531_ (.A(_0832_),
    .B(_0834_),
    .C(_0835_),
    .D_N(\top8227.PSRCurrentValue[7] ),
    .X(_0836_));
 sky130_fd_sc_hd__o311a_1 _1532_ (.A1(\top8227.PSRCurrentValue[0] ),
    .A2(_0823_),
    .A3(_0826_),
    .B1(_0831_),
    .C1(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__or4bb_1 _1533_ (.A(_0828_),
    .B(_0821_),
    .C_N(_0820_),
    .D_N(\top8227.demux.state_machine.currentInstruction[0] ),
    .X(_0838_));
 sky130_fd_sc_hd__clkbuf_4 _1534_ (.A(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__nor2_1 _1535_ (.A(_0826_),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__or4bb_1 _1536_ (.A(\top8227.demux.state_machine.currentInstruction[0] ),
    .B(\top8227.demux.state_machine.currentInstruction[3] ),
    .C_N(\top8227.demux.state_machine.currentInstruction[2] ),
    .D_N(_0828_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_4 _1537_ (.A(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__o21ai_1 _1538_ (.A1(_0826_),
    .A2(_0842_),
    .B1(\top8227.PSRCurrentValue[1] ),
    .Y(_0843_));
 sky130_fd_sc_hd__o21ai_2 _1539_ (.A1(\top8227.PSRCurrentValue[1] ),
    .A2(_0840_),
    .B1(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__or4bb_1 _1540_ (.A(\top8227.demux.state_machine.currentInstruction[0] ),
    .B(\top8227.demux.state_machine.currentInstruction[2] ),
    .C_N(\top8227.demux.state_machine.currentInstruction[3] ),
    .D_N(\top8227.demux.state_machine.currentInstruction[1] ),
    .X(_0845_));
 sky130_fd_sc_hd__buf_2 _1541_ (.A(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__or2_1 _1542_ (.A(_0826_),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__nor2_1 _1543_ (.A(_0832_),
    .B(_0835_),
    .Y(_0848_));
 sky130_fd_sc_hd__clkbuf_4 _1544_ (.A(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__buf_2 _1545_ (.A(_0828_),
    .X(_0850_));
 sky130_fd_sc_hd__clkbuf_4 _1546_ (.A(\top8227.demux.state_machine.currentInstruction[0] ),
    .X(_0851_));
 sky130_fd_sc_hd__buf_2 _1547_ (.A(_0821_),
    .X(_0852_));
 sky130_fd_sc_hd__clkbuf_2 _1548_ (.A(_0820_),
    .X(_0853_));
 sky130_fd_sc_hd__and4bb_2 _1549_ (.A_N(_0850_),
    .B_N(_0851_),
    .C(_0852_),
    .D(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _1550_ (.A(_0849_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__and4b_2 _1551_ (.A_N(_0850_),
    .B(_0851_),
    .C(_0852_),
    .D(_0853_),
    .X(_0856_));
 sky130_fd_sc_hd__nand3_1 _1552_ (.A(\top8227.PSRCurrentValue[6] ),
    .B(_0849_),
    .C(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__o221a_2 _1553_ (.A1(\top8227.PSRCurrentValue[7] ),
    .A2(_0847_),
    .B1(_0855_),
    .B2(\top8227.PSRCurrentValue[6] ),
    .C1(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__buf_2 _1554_ (.A(\top8227.demux.state_machine.timeState[6] ),
    .X(_0859_));
 sky130_fd_sc_hd__a41o_1 _1555_ (.A1(_0819_),
    .A2(_0837_),
    .A3(_0844_),
    .A4(_0858_),
    .B1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _1556_ (.A(_0823_),
    .B(_0825_),
    .Y(_0861_));
 sky130_fd_sc_hd__nor2_1 _1557_ (.A(_0830_),
    .B(_0825_),
    .Y(_0862_));
 sky130_fd_sc_hd__a21oi_1 _1558_ (.A1(_0839_),
    .A2(_0842_),
    .B1(_0825_),
    .Y(_0863_));
 sky130_fd_sc_hd__nand4b_4 _1559_ (.A_N(_0828_),
    .B(_0851_),
    .C(_0821_),
    .D(_0820_),
    .Y(_0864_));
 sky130_fd_sc_hd__or4bb_4 _1560_ (.A(_0828_),
    .B(\top8227.demux.state_machine.currentInstruction[0] ),
    .C_N(_0821_),
    .D_N(_0820_),
    .X(_0865_));
 sky130_fd_sc_hd__a41o_1 _1561_ (.A1(_0864_),
    .A2(_0834_),
    .A3(_0846_),
    .A4(_0865_),
    .B1(_0825_),
    .X(_0866_));
 sky130_fd_sc_hd__or4b_1 _1562_ (.A(_0861_),
    .B(_0862_),
    .C(_0863_),
    .D_N(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__clkbuf_4 _1563_ (.A(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__o21a_1 _1564_ (.A1(_0817_),
    .A2(_0860_),
    .B1(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__or4bb_1 _1565_ (.A(_0821_),
    .B(_0820_),
    .C_N(_0828_),
    .D_N(_0851_),
    .X(_0870_));
 sky130_fd_sc_hd__buf_4 _1566_ (.A(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__nor2_4 _1567_ (.A(_0825_),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__or2b_1 _1568_ (.A(_0835_),
    .B_N(_0832_),
    .X(_0873_));
 sky130_fd_sc_hd__buf_4 _1569_ (.A(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__or4b_1 _1570_ (.A(_0828_),
    .B(_0821_),
    .C(_0820_),
    .D_N(_0851_),
    .X(_0875_));
 sky130_fd_sc_hd__clkbuf_4 _1571_ (.A(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__nor2_2 _1572_ (.A(_0874_),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__or2b_1 _1573_ (.A(_0832_),
    .B_N(_0835_),
    .X(_0878_));
 sky130_fd_sc_hd__buf_4 _1574_ (.A(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__a21oi_1 _1575_ (.A1(_0830_),
    .A2(_0839_),
    .B1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__a21oi_2 _1576_ (.A1(_0839_),
    .A2(_0834_),
    .B1(_0874_),
    .Y(_0881_));
 sky130_fd_sc_hd__or4_2 _1577_ (.A(_0872_),
    .B(_0877_),
    .C(_0880_),
    .D(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__buf_4 _1578_ (.A(_0874_),
    .X(_0883_));
 sky130_fd_sc_hd__nor2_4 _1579_ (.A(_0883_),
    .B(_0842_),
    .Y(_0884_));
 sky130_fd_sc_hd__nand4b_4 _1580_ (.A_N(_0853_),
    .B(_0852_),
    .C(_0851_),
    .D(_0850_),
    .Y(_0885_));
 sky130_fd_sc_hd__nor2_2 _1581_ (.A(_0883_),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__or2_2 _1582_ (.A(_0884_),
    .B(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__o21a_1 _1583_ (.A1(_0882_),
    .A2(_0887_),
    .B1(_0859_),
    .X(_0888_));
 sky130_fd_sc_hd__nor2_2 _1584_ (.A(_0874_),
    .B(_0830_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_2 _1585_ (.A(_0874_),
    .B(_0823_),
    .Y(_0890_));
 sky130_fd_sc_hd__nor2_4 _1586_ (.A(_0874_),
    .B(_0871_),
    .Y(_0891_));
 sky130_fd_sc_hd__a22o_1 _1587_ (.A1(_0815_),
    .A2(_0890_),
    .B1(_0891_),
    .B2(_0819_),
    .X(_0892_));
 sky130_fd_sc_hd__and4b_1 _1588_ (.A_N(_0821_),
    .B(_0820_),
    .C(_0828_),
    .D(\top8227.demux.state_machine.currentInstruction[0] ),
    .X(_0893_));
 sky130_fd_sc_hd__clkbuf_4 _1589_ (.A(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__and2_1 _1590_ (.A(_0848_),
    .B(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__clkbuf_4 _1591_ (.A(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__and4b_1 _1592_ (.A_N(_0851_),
    .B(_0852_),
    .C(_0853_),
    .D(_0850_),
    .X(_0897_));
 sky130_fd_sc_hd__and2_2 _1593_ (.A(_0849_),
    .B(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__a22o_1 _1594_ (.A1(\top8227.demux.state_machine.timeState[3] ),
    .A2(_0896_),
    .B1(_0898_),
    .B2(_0819_),
    .X(_0899_));
 sky130_fd_sc_hd__a211o_1 _1595_ (.A1(_0815_),
    .A2(_0889_),
    .B1(_0892_),
    .C1(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__and2b_2 _1596_ (.A_N(_0832_),
    .B(_0835_),
    .X(_0901_));
 sky130_fd_sc_hd__and2_2 _1597_ (.A(_0894_),
    .B(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__and2b_2 _1598_ (.A_N(_0835_),
    .B(_0832_),
    .X(_0903_));
 sky130_fd_sc_hd__and2_2 _1599_ (.A(_0903_),
    .B(_0897_),
    .X(_0904_));
 sky130_fd_sc_hd__nor2_2 _1600_ (.A(_0883_),
    .B(_0864_),
    .Y(_0905_));
 sky130_fd_sc_hd__or3_1 _1601_ (.A(_0902_),
    .B(_0904_),
    .C(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__clkbuf_4 _1602_ (.A(\top8227.demux.state_machine.timeState[0] ),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_4 _1603_ (.A(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__and3_1 _1604_ (.A(_0908_),
    .B(_0901_),
    .C(_0854_),
    .X(_0909_));
 sky130_fd_sc_hd__a21o_1 _1605_ (.A1(_0819_),
    .A2(_0906_),
    .B1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__buf_4 _1606_ (.A(_0879_),
    .X(_0911_));
 sky130_fd_sc_hd__nor2_4 _1607_ (.A(_0911_),
    .B(_0864_),
    .Y(_0912_));
 sky130_fd_sc_hd__and2_1 _1608_ (.A(_0903_),
    .B(_0894_),
    .X(_0913_));
 sky130_fd_sc_hd__clkbuf_4 _1609_ (.A(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__nor2_2 _1610_ (.A(_0874_),
    .B(_0846_),
    .Y(_0915_));
 sky130_fd_sc_hd__clkbuf_4 _1611_ (.A(\top8227.demux.state_machine.timeState[5] ),
    .X(_0916_));
 sky130_fd_sc_hd__o31a_1 _1612_ (.A1(_0912_),
    .A2(_0914_),
    .A3(_0915_),
    .B1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__or4_2 _1613_ (.A(_0888_),
    .B(_0900_),
    .C(_0910_),
    .D(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__or4b_1 _1614_ (.A(\top8227.demux.state_machine.currentInstruction[0] ),
    .B(_0821_),
    .C(_0820_),
    .D_N(_0828_),
    .X(_0919_));
 sky130_fd_sc_hd__buf_4 _1615_ (.A(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__and4_2 _1616_ (.A(_0850_),
    .B(_0851_),
    .C(_0852_),
    .D(_0853_),
    .X(_0921_));
 sky130_fd_sc_hd__a2bb2o_1 _1617_ (.A1_N(_0874_),
    .A2_N(_0920_),
    .B1(_0921_),
    .B2(_0849_),
    .X(_0922_));
 sky130_fd_sc_hd__nor2_4 _1618_ (.A(_0879_),
    .B(_0920_),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_2 _1619_ (.A(_0911_),
    .B(_0876_),
    .Y(_0924_));
 sky130_fd_sc_hd__or4_4 _1620_ (.A(_0850_),
    .B(_0851_),
    .C(_0852_),
    .D(_0853_),
    .X(_0925_));
 sky130_fd_sc_hd__nor2_1 _1621_ (.A(_0911_),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__or4_1 _1622_ (.A(_0922_),
    .B(_0923_),
    .C(_0924_),
    .D(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nand2_4 _1623_ (.A(_0832_),
    .B(_0835_),
    .Y(_0928_));
 sky130_fd_sc_hd__a31o_1 _1624_ (.A1(_0871_),
    .A2(_0925_),
    .A3(_0920_),
    .B1(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__inv_2 _1625_ (.A(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__a21oi_1 _1626_ (.A1(_0864_),
    .A2(_0885_),
    .B1(_0928_),
    .Y(_0931_));
 sky130_fd_sc_hd__nor2_2 _1627_ (.A(_0928_),
    .B(_0842_),
    .Y(_0932_));
 sky130_fd_sc_hd__and4b_1 _1628_ (.A_N(_0852_),
    .B(_0853_),
    .C(_0832_),
    .D(_0835_),
    .X(_0933_));
 sky130_fd_sc_hd__nor2_2 _1629_ (.A(_0928_),
    .B(_0865_),
    .Y(_0934_));
 sky130_fd_sc_hd__or4_1 _1630_ (.A(_0931_),
    .B(_0932_),
    .C(_0933_),
    .D(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__or3b_2 _1631_ (.A(_0850_),
    .B(_0853_),
    .C_N(_0852_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_4 _1632_ (.A(_0928_),
    .X(_0937_));
 sky130_fd_sc_hd__nor2_1 _1633_ (.A(_0936_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__nand2_1 _1634_ (.A(_0903_),
    .B(_0921_),
    .Y(_0939_));
 sky130_fd_sc_hd__or4b_1 _1635_ (.A(_0930_),
    .B(_0935_),
    .C(_0938_),
    .D_N(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__a31oi_4 _1636_ (.A1(_0823_),
    .A2(_0871_),
    .A3(_0834_),
    .B1(_0879_),
    .Y(_0941_));
 sky130_fd_sc_hd__a21oi_1 _1637_ (.A1(_0876_),
    .A2(_0920_),
    .B1(_0826_),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_2 _1638_ (.A(_0883_),
    .B(_0925_),
    .Y(_0943_));
 sky130_fd_sc_hd__and2_2 _1639_ (.A(_0901_),
    .B(_0921_),
    .X(_0944_));
 sky130_fd_sc_hd__or3_1 _1640_ (.A(_0942_),
    .B(_0943_),
    .C(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__nor2_1 _1641_ (.A(_0911_),
    .B(_0842_),
    .Y(_0946_));
 sky130_fd_sc_hd__nor2_1 _1642_ (.A(_0879_),
    .B(_0846_),
    .Y(_0947_));
 sky130_fd_sc_hd__or2_1 _1643_ (.A(_0946_),
    .B(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__nor2_4 _1644_ (.A(_0879_),
    .B(_0885_),
    .Y(_0949_));
 sky130_fd_sc_hd__nor2_4 _1645_ (.A(_0825_),
    .B(_0885_),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_2 _1646_ (.A(_0883_),
    .B(_0865_),
    .Y(_0951_));
 sky130_fd_sc_hd__and2_2 _1647_ (.A(_0901_),
    .B(_0897_),
    .X(_0952_));
 sky130_fd_sc_hd__or4_1 _1648_ (.A(_0949_),
    .B(_0950_),
    .C(_0951_),
    .D(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__or4_1 _1649_ (.A(_0941_),
    .B(_0945_),
    .C(_0948_),
    .D(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__clkbuf_4 _1650_ (.A(_0819_),
    .X(_0955_));
 sky130_fd_sc_hd__o31a_1 _1651_ (.A1(_0927_),
    .A2(_0940_),
    .A3(_0954_),
    .B1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__inv_2 _1652_ (.A(\top8227.demux.state_machine.timeState[4] ),
    .Y(_0957_));
 sky130_fd_sc_hd__or3_1 _1653_ (.A(_0957_),
    .B(_0874_),
    .C(_0936_),
    .X(_0958_));
 sky130_fd_sc_hd__nand2_1 _1654_ (.A(_0849_),
    .B(_0894_),
    .Y(_0959_));
 sky130_fd_sc_hd__nor2_2 _1655_ (.A(\top8227.demux.state_machine.timeState[2] ),
    .B(\top8227.demux.state_machine.timeState[6] ),
    .Y(_0960_));
 sky130_fd_sc_hd__or3_1 _1656_ (.A(_0960_),
    .B(_0879_),
    .C(_0864_),
    .X(_0961_));
 sky130_fd_sc_hd__nor3_1 _1657_ (.A(\top8227.demux.state_machine.timeState[4] ),
    .B(_0814_),
    .C(\top8227.demux.state_machine.timeState[6] ),
    .Y(_0962_));
 sky130_fd_sc_hd__o211a_1 _1658_ (.A1(\top8227.demux.reset ),
    .A2(_0962_),
    .B1(_0894_),
    .C1(_0849_),
    .X(_0963_));
 sky130_fd_sc_hd__a31oi_1 _1659_ (.A1(_0958_),
    .A2(_0959_),
    .A3(_0961_),
    .B1(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__or2_2 _1660_ (.A(\top8227.demux.state_machine.timeState[4] ),
    .B(_0814_),
    .X(_0965_));
 sky130_fd_sc_hd__o41a_1 _1661_ (.A1(_0872_),
    .A2(_0877_),
    .A3(_0880_),
    .A4(_0881_),
    .B1(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__or2_1 _1662_ (.A(_0907_),
    .B(_0929_),
    .X(_0967_));
 sky130_fd_sc_hd__o31a_2 _1663_ (.A1(_0964_),
    .A2(_0930_),
    .A3(_0966_),
    .B1(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__or2_2 _1664_ (.A(\top8227.pulse_slower.currentEnableState[1] ),
    .B(\top8227.pulse_slower.currentEnableState[0] ),
    .X(_0969_));
 sky130_fd_sc_hd__inv_2 _1665_ (.A(_0969_),
    .Y(\top8227.pulse_slower.nextEnableState[0] ));
 sky130_fd_sc_hd__nor4_1 _1666_ (.A(\top8227.demux.state_machine.currentAddress[8] ),
    .B(\top8227.demux.state_machine.currentAddress[0] ),
    .C(\top8227.demux.state_machine.currentAddress[2] ),
    .D(\top8227.demux.state_machine.currentAddress[9] ),
    .Y(_0970_));
 sky130_fd_sc_hd__nand2_4 _1667_ (.A(\top8227.demux.isAddressing ),
    .B(net33),
    .Y(_0971_));
 sky130_fd_sc_hd__o211a_4 _1668_ (.A1(gpio[19]),
    .A2(_0968_),
    .B1(\top8227.pulse_slower.nextEnableState[0] ),
    .C1(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__o31ai_4 _1669_ (.A1(_0869_),
    .A2(_0918_),
    .A3(_0956_),
    .B1(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__clkinv_4 _1670_ (.A(net29),
    .Y(gpio[21]));
 sky130_fd_sc_hd__a21o_1 _1671_ (.A1(_0971_),
    .A2(_0968_),
    .B1(gpio[19]),
    .X(_0974_));
 sky130_fd_sc_hd__nand2_1 _1672_ (.A(\top8227.pulse_slower.nextEnableState[0] ),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__buf_4 _1673_ (.A(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__nor2_1 _1674_ (.A(\top8227.instructionLoader.interruptInjector.resetDetected ),
    .B(gpio[21]),
    .Y(_0977_));
 sky130_fd_sc_hd__nor2_2 _1675_ (.A(_0976_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__buf_4 _1676_ (.A(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__and2_1 _1677_ (.A(\top8227.demux.isAddressing ),
    .B(net33),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_4 _1678_ (.A(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__clkbuf_4 _1679_ (.A(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a21oi_2 _1680_ (.A1(_0971_),
    .A2(_0968_),
    .B1(gpio[19]),
    .Y(_0983_));
 sky130_fd_sc_hd__nor2_1 _1681_ (.A(_0969_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__clkbuf_4 _1682_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__buf_4 _1683_ (.A(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_4 _1684_ (.A(\top8227.demux.state_machine.currentAddress[1] ),
    .X(_0987_));
 sky130_fd_sc_hd__nor2_1 _1685_ (.A(_0987_),
    .B(\top8227.demux.state_machine.currentAddress[12] ),
    .Y(_0988_));
 sky130_fd_sc_hd__and2b_1 _1686_ (.A_N(\top8227.demux.state_machine.currentAddress[6] ),
    .B(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__nor2_1 _1687_ (.A(_0907_),
    .B(_0818_),
    .Y(_0990_));
 sky130_fd_sc_hd__and2b_1 _1688_ (.A_N(_0814_),
    .B(_0859_),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_2 _1689_ (.A(_0990_),
    .B(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__clkbuf_4 _1690_ (.A(_0907_),
    .X(_0993_));
 sky130_fd_sc_hd__o31ai_1 _1691_ (.A1(\top8227.demux.state_machine.currentAddress[7] ),
    .A2(\top8227.demux.state_machine.currentAddress[3] ),
    .A3(\top8227.demux.state_machine.currentAddress[11] ),
    .B1(_0818_),
    .Y(_0994_));
 sky130_fd_sc_hd__nor2_1 _1692_ (.A(\top8227.demux.state_machine.currentAddress[10] ),
    .B(\top8227.demux.state_machine.currentAddress[4] ),
    .Y(_0995_));
 sky130_fd_sc_hd__or3b_2 _1693_ (.A(_0907_),
    .B(_0818_),
    .C_N(_0814_),
    .X(_0996_));
 sky130_fd_sc_hd__nand2_1 _1694_ (.A(_0907_),
    .B(\top8227.demux.state_machine.currentAddress[5] ),
    .Y(_0997_));
 sky130_fd_sc_hd__o221a_1 _1695_ (.A1(_0993_),
    .A2(_0994_),
    .B1(_0995_),
    .B2(_0996_),
    .C1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__o21ai_1 _1696_ (.A1(_0989_),
    .A2(_0992_),
    .B1(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__and3_2 _1697_ (.A(_0982_),
    .B(_0986_),
    .C(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__clkbuf_4 _1698_ (.A(_0993_),
    .X(_1001_));
 sky130_fd_sc_hd__buf_2 _1699_ (.A(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__buf_2 _1700_ (.A(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_4 _1701_ (.A(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_4 _1702_ (.A(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__buf_4 _1703_ (.A(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(_1006_),
    .A1(\top8227.demux.state_machine.timeState[3] ),
    .S(_0986_),
    .X(_1007_));
 sky130_fd_sc_hd__or3_1 _1705_ (.A(_0979_),
    .B(_1000_),
    .C(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_1 _1706_ (.A(_1008_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _1707_ (.A(\top8227.demux.state_machine.timeState[1] ),
    .X(_1009_));
 sky130_fd_sc_hd__buf_4 _1708_ (.A(_0976_),
    .X(_1010_));
 sky130_fd_sc_hd__and3b_1 _1709_ (.A_N(_1000_),
    .B(_0977_),
    .C(_0986_),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_2 _1710_ (.A(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_4 _1711_ (.A(_0859_),
    .X(_1013_));
 sky130_fd_sc_hd__a22o_1 _1712_ (.A1(_1009_),
    .A2(_1010_),
    .B1(_1012_),
    .B2(_1013_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _1713_ (.A(_0815_),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_4 _1714_ (.A(_0955_),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_1 _1715_ (.A1(_1014_),
    .A2(_1010_),
    .B1(_1012_),
    .B2(_1015_),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _1716_ (.A1(net73),
    .A2(_1010_),
    .B1(_1012_),
    .B2(_0916_),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _1717_ (.A1(_1015_),
    .A2(_1010_),
    .B1(_1012_),
    .B2(_1006_),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_1 _1718_ (.A1(_0916_),
    .A2(_1010_),
    .B1(_1012_),
    .B2(_1009_),
    .X(_0018_));
 sky130_fd_sc_hd__a22o_1 _1719_ (.A1(_1013_),
    .A2(_1010_),
    .B1(_1012_),
    .B2(_1014_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _1720_ (.A(\top8227.demux.state_machine.currentAddress[7] ),
    .X(_1016_));
 sky130_fd_sc_hd__nor3_4 _1721_ (.A(\top8227.demux.nmi ),
    .B(\top8227.instructionLoader.interruptInjector.resetDetected ),
    .C(\top8227.instructionLoader.interruptInjector.irqGenerated ),
    .Y(_1017_));
 sky130_fd_sc_hd__clkbuf_4 _1722_ (.A(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__o21ai_1 _1723_ (.A1(net1),
    .A2(net2),
    .B1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__clkbuf_4 _1724_ (.A(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__buf_4 _1725_ (.A(net8),
    .X(_1021_));
 sky130_fd_sc_hd__nand2_1 _1726_ (.A(net7),
    .B(_1017_),
    .Y(_1022_));
 sky130_fd_sc_hd__nor2_1 _1727_ (.A(_1021_),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__and2_2 _1728_ (.A(net6),
    .B(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__buf_2 _1729_ (.A(net5),
    .X(_1025_));
 sky130_fd_sc_hd__nand3_1 _1730_ (.A(net4),
    .B(net3),
    .C(_1018_),
    .Y(_1026_));
 sky130_fd_sc_hd__or2_1 _1731_ (.A(_1025_),
    .B(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a21oi_1 _1732_ (.A1(_1020_),
    .A2(_1024_),
    .B1(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(_1016_),
    .A1(_1028_),
    .S(_0979_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_1 _1734_ (.A(_1029_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_2 _1735_ (.A(_0976_),
    .B(_0977_),
    .X(_1030_));
 sky130_fd_sc_hd__clkbuf_4 _1736_ (.A(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__buf_2 _1737_ (.A(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__clkbuf_4 _1738_ (.A(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__clkbuf_4 _1739_ (.A(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_4 _1740_ (.A(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__nor2_1 _1741_ (.A(_1025_),
    .B(_1026_),
    .Y(_1036_));
 sky130_fd_sc_hd__and2_1 _1742_ (.A(_0978_),
    .B(_1019_),
    .X(_1037_));
 sky130_fd_sc_hd__clkbuf_4 _1743_ (.A(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__and3_1 _1744_ (.A(_1023_),
    .B(_1036_),
    .C(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__buf_2 _1745_ (.A(net6),
    .X(_1040_));
 sky130_fd_sc_hd__a22o_1 _1746_ (.A1(\top8227.demux.state_machine.currentAddress[6] ),
    .A2(_1035_),
    .B1(_1039_),
    .B2(_1040_),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_2 _1747_ (.A(net2),
    .B(_1017_),
    .Y(_1041_));
 sky130_fd_sc_hd__nand2_1 _1748_ (.A(net4),
    .B(_1017_),
    .Y(_1042_));
 sky130_fd_sc_hd__nand2_1 _1749_ (.A(net3),
    .B(_1017_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _1750_ (.A(_1042_),
    .B(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__o21ai_1 _1751_ (.A1(_1041_),
    .A2(_1044_),
    .B1(_1026_),
    .Y(_1045_));
 sky130_fd_sc_hd__and3_1 _1752_ (.A(_1025_),
    .B(_0979_),
    .C(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__a21o_1 _1753_ (.A1(net60),
    .A2(_1035_),
    .B1(_1046_),
    .X(_0007_));
 sky130_fd_sc_hd__or2_2 _1754_ (.A(net4),
    .B(_1043_),
    .X(_1047_));
 sky130_fd_sc_hd__and4bb_1 _1755_ (.A_N(_0977_),
    .B_N(_1047_),
    .C(_1025_),
    .D(_0986_),
    .X(_1048_));
 sky130_fd_sc_hd__nand2_2 _1756_ (.A(_1021_),
    .B(_1017_),
    .Y(_1049_));
 sky130_fd_sc_hd__nor2_1 _1757_ (.A(net7),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__a32o_1 _1758_ (.A1(net2),
    .A2(_1048_),
    .A3(_1050_),
    .B1(_1035_),
    .B2(net58),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_2 _1759_ (.A(net5),
    .B(_1017_),
    .Y(_1051_));
 sky130_fd_sc_hd__nor2_2 _1760_ (.A(_1044_),
    .B(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__and3_2 _1761_ (.A(_0979_),
    .B(_1020_),
    .C(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__a21o_1 _1762_ (.A1(net54),
    .A2(_1035_),
    .B1(_1053_),
    .X(_0011_));
 sky130_fd_sc_hd__and4b_1 _1763_ (.A_N(net2),
    .B(_0978_),
    .C(_1018_),
    .D(net1),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_4 _1764_ (.A(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__or2_2 _1765_ (.A(net3),
    .B(_1042_),
    .X(_1056_));
 sky130_fd_sc_hd__nor2_2 _1766_ (.A(_1025_),
    .B(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__nor2_1 _1767_ (.A(_1041_),
    .B(_1044_),
    .Y(_1058_));
 sky130_fd_sc_hd__and3_1 _1768_ (.A(_0978_),
    .B(_1058_),
    .C(_1051_),
    .X(_1059_));
 sky130_fd_sc_hd__inv_2 _1769_ (.A(_1049_),
    .Y(_1060_));
 sky130_fd_sc_hd__and3_1 _1770_ (.A(_1042_),
    .B(_1043_),
    .C(_1051_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_4 _1771_ (.A(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__a32o_1 _1772_ (.A1(_1038_),
    .A2(_1060_),
    .A3(_1062_),
    .B1(_1034_),
    .B2(net91),
    .X(_1063_));
 sky130_fd_sc_hd__a211o_1 _1773_ (.A1(_1055_),
    .A2(_1057_),
    .B1(_1059_),
    .C1(_1063_),
    .X(_0005_));
 sky130_fd_sc_hd__nor2_1 _1774_ (.A(_1025_),
    .B(_1047_),
    .Y(_1064_));
 sky130_fd_sc_hd__nor2_1 _1775_ (.A(_1041_),
    .B(_1050_),
    .Y(_1065_));
 sky130_fd_sc_hd__nor2_1 _1776_ (.A(_1034_),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__a22o_1 _1777_ (.A1(\top8227.demux.state_machine.currentAddress[5] ),
    .A2(_1035_),
    .B1(_1064_),
    .B2(_1066_),
    .X(_0008_));
 sky130_fd_sc_hd__o21a_1 _1778_ (.A1(_1021_),
    .A2(_1047_),
    .B1(_1056_),
    .X(_1067_));
 sky130_fd_sc_hd__or4_1 _1779_ (.A(_1025_),
    .B(_1034_),
    .C(_1041_),
    .D(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__a21bo_1 _1780_ (.A1(net59),
    .A2(_1035_),
    .B1_N(_1068_),
    .X(_0000_));
 sky130_fd_sc_hd__a22o_1 _1781_ (.A1(_0987_),
    .A2(_1035_),
    .B1(_1052_),
    .B2(_1055_),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _1782_ (.A1(\top8227.demux.state_machine.currentAddress[12] ),
    .A2(_1035_),
    .B1(_1055_),
    .B2(_1062_),
    .X(_0003_));
 sky130_fd_sc_hd__nand2_1 _1783_ (.A(net2),
    .B(_1050_),
    .Y(_1069_));
 sky130_fd_sc_hd__a22o_1 _1784_ (.A1(net61),
    .A2(_1035_),
    .B1(_1048_),
    .B2(_1069_),
    .X(_0002_));
 sky130_fd_sc_hd__nor2_1 _1785_ (.A(net3),
    .B(_1042_),
    .Y(_1070_));
 sky130_fd_sc_hd__and2_1 _1786_ (.A(_1025_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_4 _1787_ (.A(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__a22o_1 _1788_ (.A1(net77),
    .A2(_1035_),
    .B1(_1055_),
    .B2(_1072_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_2 _1789_ (.A(_1070_),
    .B(_1062_),
    .X(_1073_));
 sky130_fd_sc_hd__nand2_1 _1790_ (.A(_1060_),
    .B(_1056_),
    .Y(_1074_));
 sky130_fd_sc_hd__a32o_1 _1791_ (.A1(_1020_),
    .A2(_1073_),
    .A3(_1074_),
    .B1(_1072_),
    .B2(net2),
    .X(_1075_));
 sky130_fd_sc_hd__a31o_1 _1792_ (.A1(_1060_),
    .A2(_1064_),
    .A3(_1065_),
    .B1(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(\top8227.demux.state_machine.currentAddress[9] ),
    .A1(_1076_),
    .S(_0979_),
    .X(_1077_));
 sky130_fd_sc_hd__clkbuf_1 _1794_ (.A(_1077_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_4 _1795_ (.A(_0971_),
    .X(_1078_));
 sky130_fd_sc_hd__and2_2 _1796_ (.A(_1078_),
    .B(_0968_),
    .X(_1079_));
 sky130_fd_sc_hd__inv_2 _1797_ (.A(_1079_),
    .Y(gpio[22]));
 sky130_fd_sc_hd__and4b_2 _1798_ (.A_N(_1040_),
    .B(_1021_),
    .C(net7),
    .D(_1018_),
    .X(_1080_));
 sky130_fd_sc_hd__a32o_1 _1799_ (.A1(_1037_),
    .A2(_1057_),
    .A3(_1080_),
    .B1(_1031_),
    .B2(_0902_),
    .X(_1081_));
 sky130_fd_sc_hd__and3_1 _1800_ (.A(_0978_),
    .B(_1019_),
    .C(_1024_),
    .X(_1082_));
 sky130_fd_sc_hd__a22o_1 _1801_ (.A1(_0914_),
    .A2(_1031_),
    .B1(_1062_),
    .B2(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__and2_1 _1802_ (.A(_0832_),
    .B(_0835_),
    .X(_1084_));
 sky130_fd_sc_hd__and2b_2 _1803_ (.A_N(_1040_),
    .B(_1023_),
    .X(_1085_));
 sky130_fd_sc_hd__nor2_2 _1804_ (.A(net29),
    .B(_1041_),
    .Y(_1086_));
 sky130_fd_sc_hd__and2_2 _1805_ (.A(_1057_),
    .B(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__a32o_1 _1806_ (.A1(_0894_),
    .A2(_1084_),
    .A3(_1031_),
    .B1(_1085_),
    .B2(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__or3_1 _1807_ (.A(_1081_),
    .B(_1083_),
    .C(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__nor2_2 _1808_ (.A(_0871_),
    .B(_0928_),
    .Y(_1090_));
 sky130_fd_sc_hd__clkbuf_4 _1809_ (.A(_1030_),
    .X(_1091_));
 sky130_fd_sc_hd__clkbuf_4 _1810_ (.A(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__or3_1 _1811_ (.A(_1040_),
    .B(net7),
    .C(_1049_),
    .X(_1093_));
 sky130_fd_sc_hd__a21oi_1 _1812_ (.A1(_1027_),
    .A2(_1047_),
    .B1(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__a22o_1 _1813_ (.A1(_1090_),
    .A2(_1092_),
    .B1(_1038_),
    .B2(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__buf_4 _1814_ (.A(_0896_),
    .X(_1096_));
 sky130_fd_sc_hd__nand2_2 _1815_ (.A(_1022_),
    .B(_1049_),
    .Y(_1097_));
 sky130_fd_sc_hd__a21oi_4 _1816_ (.A1(_1040_),
    .A2(_1018_),
    .B1(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__and3_1 _1817_ (.A(_0979_),
    .B(_1020_),
    .C(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__a22o_1 _1818_ (.A1(_1096_),
    .A2(_1032_),
    .B1(_1062_),
    .B2(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__a2bb2o_1 _1819_ (.A1_N(_0939_),
    .A2_N(_0978_),
    .B1(_1072_),
    .B2(_1082_),
    .X(_1101_));
 sky130_fd_sc_hd__nor4_2 _1820_ (.A(_0976_),
    .B(net29),
    .C(_1041_),
    .D(_1073_),
    .Y(_1102_));
 sky130_fd_sc_hd__and2_2 _1821_ (.A(_1040_),
    .B(_1050_),
    .X(_1103_));
 sky130_fd_sc_hd__a221o_1 _1822_ (.A1(_0944_),
    .A2(_1030_),
    .B1(_1102_),
    .B2(_1103_),
    .C1(_1059_),
    .X(_1104_));
 sky130_fd_sc_hd__a31o_1 _1823_ (.A1(_1037_),
    .A2(_1072_),
    .A3(_1080_),
    .B1(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__a311o_1 _1824_ (.A1(_0849_),
    .A2(_0921_),
    .A3(_1032_),
    .B1(_1101_),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__and4bb_2 _1825_ (.A_N(_1021_),
    .B_N(net7),
    .C(_1018_),
    .D(_1040_),
    .X(_1107_));
 sky130_fd_sc_hd__and3_2 _1826_ (.A(_0978_),
    .B(_1019_),
    .C(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__a22o_1 _1827_ (.A1(_0886_),
    .A2(_1032_),
    .B1(_1057_),
    .B2(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__nor2_1 _1828_ (.A(_0937_),
    .B(_0885_),
    .Y(_1110_));
 sky130_fd_sc_hd__and2b_2 _1829_ (.A_N(_1040_),
    .B(_1050_),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _1830_ (.A1(_1110_),
    .A2(_1032_),
    .B1(_1087_),
    .B2(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__and2_1 _1831_ (.A(_0978_),
    .B(_1057_),
    .X(_1113_));
 sky130_fd_sc_hd__a32o_1 _1832_ (.A1(_1020_),
    .A2(_1111_),
    .A3(_1113_),
    .B1(_1091_),
    .B2(_0949_),
    .X(_1114_));
 sky130_fd_sc_hd__inv_2 _1833_ (.A(_1097_),
    .Y(_1115_));
 sky130_fd_sc_hd__a32o_1 _1834_ (.A1(_1038_),
    .A2(_1064_),
    .A3(_1115_),
    .B1(_1091_),
    .B2(_0950_),
    .X(_1116_));
 sky130_fd_sc_hd__a211o_1 _1835_ (.A1(_1036_),
    .A2(_1108_),
    .B1(_1114_),
    .C1(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__or4_1 _1836_ (.A(_1106_),
    .B(_1109_),
    .C(_1112_),
    .D(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__or4_1 _1837_ (.A(_1089_),
    .B(_1095_),
    .C(_1100_),
    .D(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_1 _1838_ (.A(_0830_),
    .B(_0911_),
    .Y(_1120_));
 sky130_fd_sc_hd__nor2_1 _1839_ (.A(_0830_),
    .B(_0937_),
    .Y(_1121_));
 sky130_fd_sc_hd__a32o_1 _1840_ (.A1(_1020_),
    .A2(_1103_),
    .A3(_1113_),
    .B1(_1091_),
    .B2(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__a221o_1 _1841_ (.A1(_1120_),
    .A2(_1092_),
    .B1(_1080_),
    .B2(net26),
    .C1(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__a32o_1 _1842_ (.A1(_0849_),
    .A2(_0856_),
    .A3(_1032_),
    .B1(_1024_),
    .B2(_1053_),
    .X(_1124_));
 sky130_fd_sc_hd__a221o_1 _1843_ (.A1(_0862_),
    .A2(_1034_),
    .B1(_1053_),
    .B2(_1103_),
    .C1(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__a22o_1 _1844_ (.A1(_0905_),
    .A2(_1031_),
    .B1(_1072_),
    .B2(_1108_),
    .X(_1126_));
 sky130_fd_sc_hd__buf_4 _1845_ (.A(_0912_),
    .X(_1127_));
 sky130_fd_sc_hd__a22o_1 _1846_ (.A1(_1127_),
    .A2(_1031_),
    .B1(_1062_),
    .B2(_1108_),
    .X(_1128_));
 sky130_fd_sc_hd__or2_1 _1847_ (.A(_1126_),
    .B(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__and3_1 _1848_ (.A(_1025_),
    .B(_0978_),
    .C(_1070_),
    .X(_1130_));
 sky130_fd_sc_hd__nor2_1 _1849_ (.A(_0864_),
    .B(_0937_),
    .Y(_1131_));
 sky130_fd_sc_hd__a32o_1 _1850_ (.A1(_1020_),
    .A2(_1111_),
    .A3(_1130_),
    .B1(_1032_),
    .B2(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__a221o_1 _1851_ (.A1(_0889_),
    .A2(_1034_),
    .B1(_1057_),
    .B2(_1099_),
    .C1(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__or4_1 _1852_ (.A(_1123_),
    .B(_1125_),
    .C(_1129_),
    .D(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__nor2_1 _1853_ (.A(_0911_),
    .B(_0871_),
    .Y(_1135_));
 sky130_fd_sc_hd__nor2_1 _1854_ (.A(_1023_),
    .B(_1107_),
    .Y(_1136_));
 sky130_fd_sc_hd__a22o_1 _1855_ (.A1(_1064_),
    .A2(_1097_),
    .B1(_1136_),
    .B2(_1036_),
    .X(_1137_));
 sky130_fd_sc_hd__a21o_1 _1856_ (.A1(_1060_),
    .A2(_1062_),
    .B1(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__or2_1 _1857_ (.A(_1080_),
    .B(_1103_),
    .X(_1139_));
 sky130_fd_sc_hd__inv_2 _1858_ (.A(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__o311a_1 _1859_ (.A1(net7),
    .A2(_1049_),
    .A3(_1062_),
    .B1(_1138_),
    .C1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _1860_ (.A1(_1135_),
    .A2(_1092_),
    .B1(_1038_),
    .B2(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__a22o_1 _1861_ (.A1(_0891_),
    .A2(_1092_),
    .B1(_1055_),
    .B2(_1098_),
    .X(_1143_));
 sky130_fd_sc_hd__a22o_1 _1862_ (.A1(_0872_),
    .A2(_1033_),
    .B1(_1098_),
    .B2(net26),
    .X(_1144_));
 sky130_fd_sc_hd__or3_1 _1863_ (.A(_1142_),
    .B(_1143_),
    .C(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__nor2_2 _1864_ (.A(_0911_),
    .B(_0839_),
    .Y(_1146_));
 sky130_fd_sc_hd__nor4_1 _1865_ (.A(_1049_),
    .B(_1073_),
    .C(_1094_),
    .D(_1139_),
    .Y(_1147_));
 sky130_fd_sc_hd__nor2_1 _1866_ (.A(_0839_),
    .B(_0937_),
    .Y(_1148_));
 sky130_fd_sc_hd__a22o_1 _1867_ (.A1(_1087_),
    .A2(_1098_),
    .B1(_1148_),
    .B2(_1030_),
    .X(_1149_));
 sky130_fd_sc_hd__a221o_1 _1868_ (.A1(_1146_),
    .A2(_1031_),
    .B1(_1086_),
    .B2(_1147_),
    .C1(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__nor2_2 _1869_ (.A(_0874_),
    .B(_0839_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand2_1 _1870_ (.A(net2),
    .B(_1024_),
    .Y(_1152_));
 sky130_fd_sc_hd__or3_1 _1871_ (.A(_0976_),
    .B(_1073_),
    .C(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__o2bb2a_1 _1872_ (.A1_N(_1151_),
    .A2_N(_1030_),
    .B1(_1153_),
    .B2(_0977_),
    .X(_1154_));
 sky130_fd_sc_hd__inv_2 _1873_ (.A(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__a32o_1 _1874_ (.A1(_1037_),
    .A2(_1052_),
    .A3(_1080_),
    .B1(_1031_),
    .B2(_0840_),
    .X(_1156_));
 sky130_fd_sc_hd__or3_1 _1875_ (.A(_1150_),
    .B(_1155_),
    .C(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__nor2_1 _1876_ (.A(_0826_),
    .B(_0876_),
    .Y(_1158_));
 sky130_fd_sc_hd__a22o_1 _1877_ (.A1(_0877_),
    .A2(_1031_),
    .B1(_1085_),
    .B2(_1102_),
    .X(_1159_));
 sky130_fd_sc_hd__a221o_1 _1878_ (.A1(_1158_),
    .A2(_1034_),
    .B1(_1024_),
    .B2(_1055_),
    .C1(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__a32o_1 _1879_ (.A1(_1020_),
    .A2(_1103_),
    .A3(_1130_),
    .B1(_1033_),
    .B2(_0924_),
    .X(_1161_));
 sky130_fd_sc_hd__or4_1 _1880_ (.A(_1145_),
    .B(_1157_),
    .C(_1160_),
    .D(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__or3_1 _1881_ (.A(_1119_),
    .B(_1134_),
    .C(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__clkbuf_1 _1882_ (.A(_1163_),
    .X(_0020_));
 sky130_fd_sc_hd__and4_2 _1883_ (.A(_1040_),
    .B(_1021_),
    .C(net7),
    .D(_1018_),
    .X(_1164_));
 sky130_fd_sc_hd__a32o_1 _1884_ (.A1(_1020_),
    .A2(_1130_),
    .A3(_1164_),
    .B1(_1091_),
    .B2(_0904_),
    .X(_1165_));
 sky130_fd_sc_hd__a221o_1 _1885_ (.A1(_0898_),
    .A2(_1092_),
    .B1(_1072_),
    .B2(_1099_),
    .C1(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__a32o_1 _1886_ (.A1(_1072_),
    .A2(_1086_),
    .A3(_1093_),
    .B1(_1091_),
    .B2(_0932_),
    .X(_1167_));
 sky130_fd_sc_hd__a221o_1 _1887_ (.A1(_0884_),
    .A2(_1092_),
    .B1(_1057_),
    .B2(_1082_),
    .C1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__a22o_1 _1888_ (.A1(_0952_),
    .A2(_1091_),
    .B1(_1054_),
    .B2(_1103_),
    .X(_1169_));
 sky130_fd_sc_hd__a221o_1 _1889_ (.A1(_0946_),
    .A2(_1092_),
    .B1(_1080_),
    .B2(_1087_),
    .C1(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__or3_1 _1890_ (.A(_1166_),
    .B(_1168_),
    .C(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__nor2_1 _1891_ (.A(_0826_),
    .B(_0842_),
    .Y(_1172_));
 sky130_fd_sc_hd__a22o_1 _1892_ (.A1(_1172_),
    .A2(_1092_),
    .B1(_1053_),
    .B2(_1164_),
    .X(_1173_));
 sky130_fd_sc_hd__a2bb2o_1 _1893_ (.A1_N(_0847_),
    .A2_N(_0979_),
    .B1(_1053_),
    .B2(_1098_),
    .X(_1174_));
 sky130_fd_sc_hd__nor2_1 _1894_ (.A(_0937_),
    .B(_0920_),
    .Y(_1175_));
 sky130_fd_sc_hd__a221oi_1 _1895_ (.A1(_1040_),
    .A2(_1018_),
    .B1(_1027_),
    .B2(_1047_),
    .C1(_1069_),
    .Y(_1176_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(_1175_),
    .A1(_1176_),
    .S(_0978_),
    .X(_1177_));
 sky130_fd_sc_hd__a221o_1 _1897_ (.A1(_0923_),
    .A2(_1092_),
    .B1(_1054_),
    .B2(_1080_),
    .C1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__nor2_1 _1898_ (.A(_0826_),
    .B(_0920_),
    .Y(_1179_));
 sky130_fd_sc_hd__nor2_1 _1899_ (.A(_0883_),
    .B(_0920_),
    .Y(_1180_));
 sky130_fd_sc_hd__a22o_1 _1900_ (.A1(_1180_),
    .A2(_1091_),
    .B1(_1087_),
    .B2(_1164_),
    .X(_1181_));
 sky130_fd_sc_hd__a221o_1 _1901_ (.A1(_1179_),
    .A2(_1092_),
    .B1(_1055_),
    .B2(_1107_),
    .C1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__or4_1 _1902_ (.A(_1173_),
    .B(_1174_),
    .C(_1178_),
    .D(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_4 _1903_ (.A(_0915_),
    .X(_1184_));
 sky130_fd_sc_hd__a32o_1 _1904_ (.A1(_1038_),
    .A2(_1062_),
    .A3(_1085_),
    .B1(_1033_),
    .B2(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__nor2_1 _1905_ (.A(_0937_),
    .B(_0846_),
    .Y(_1186_));
 sky130_fd_sc_hd__a22o_1 _1906_ (.A1(_1087_),
    .A2(_1107_),
    .B1(_1186_),
    .B2(_1031_),
    .X(_1187_));
 sky130_fd_sc_hd__a32o_1 _1907_ (.A1(_1020_),
    .A2(_1113_),
    .A3(_1164_),
    .B1(_1032_),
    .B2(_0947_),
    .X(_1188_));
 sky130_fd_sc_hd__or2_1 _1908_ (.A(_1187_),
    .B(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__or2_1 _1909_ (.A(_1185_),
    .B(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__or4_1 _1910_ (.A(_1145_),
    .B(_1171_),
    .C(_1183_),
    .D(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__or2_1 _1911_ (.A(_1119_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_1 _1912_ (.A(_1192_),
    .X(_0021_));
 sky130_fd_sc_hd__a2bb2o_1 _1913_ (.A1_N(_0855_),
    .A2_N(_0979_),
    .B1(_1053_),
    .B2(_1085_),
    .X(_1193_));
 sky130_fd_sc_hd__a32o_1 _1914_ (.A1(_1038_),
    .A2(_1057_),
    .A3(_1085_),
    .B1(_1033_),
    .B2(_0890_),
    .X(_1194_));
 sky130_fd_sc_hd__nor2_2 _1915_ (.A(_0823_),
    .B(_0911_),
    .Y(_1195_));
 sky130_fd_sc_hd__and4_1 _1916_ (.A(_1038_),
    .B(_1051_),
    .C(_1056_),
    .D(_1080_),
    .X(_1196_));
 sky130_fd_sc_hd__nor2_1 _1917_ (.A(_0823_),
    .B(_0937_),
    .Y(_1197_));
 sky130_fd_sc_hd__a22o_1 _1918_ (.A1(_1197_),
    .A2(_1091_),
    .B1(_1087_),
    .B2(_1103_),
    .X(_1198_));
 sky130_fd_sc_hd__a211o_1 _1919_ (.A1(_1195_),
    .A2(_1033_),
    .B1(_1196_),
    .C1(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__or3_1 _1920_ (.A(_1193_),
    .B(_1194_),
    .C(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__a22o_1 _1921_ (.A1(_0951_),
    .A2(_1033_),
    .B1(_1055_),
    .B2(_1164_),
    .X(_1201_));
 sky130_fd_sc_hd__a22o_1 _1922_ (.A1(_0934_),
    .A2(_1032_),
    .B1(_1024_),
    .B2(_1087_),
    .X(_1202_));
 sky130_fd_sc_hd__a31o_1 _1923_ (.A1(_0901_),
    .A2(_0854_),
    .A3(_1033_),
    .B1(_1039_),
    .X(_1203_));
 sky130_fd_sc_hd__or3_1 _1924_ (.A(_1201_),
    .B(_1202_),
    .C(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__a221o_1 _1925_ (.A1(_0861_),
    .A2(_1034_),
    .B1(_1053_),
    .B2(_1111_),
    .C1(_1173_),
    .X(_1205_));
 sky130_fd_sc_hd__or4_1 _1926_ (.A(_1171_),
    .B(_1200_),
    .C(_1204_),
    .D(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__or3_1 _1927_ (.A(_1118_),
    .B(_1134_),
    .C(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _1928_ (.A(_1207_),
    .X(_0022_));
 sky130_fd_sc_hd__or4_1 _1929_ (.A(_1089_),
    .B(_1106_),
    .C(_1129_),
    .D(_1157_),
    .X(_1208_));
 sky130_fd_sc_hd__nor2_4 _1930_ (.A(_0911_),
    .B(_0834_),
    .Y(_1209_));
 sky130_fd_sc_hd__a22o_1 _1931_ (.A1(_1209_),
    .A2(_1033_),
    .B1(_1055_),
    .B2(_1085_),
    .X(_1210_));
 sky130_fd_sc_hd__a211o_1 _1932_ (.A1(_1052_),
    .A2(_1108_),
    .B1(_1169_),
    .C1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__nor2_2 _1933_ (.A(_0883_),
    .B(_0834_),
    .Y(_1212_));
 sky130_fd_sc_hd__a22o_1 _1934_ (.A1(_1212_),
    .A2(_1091_),
    .B1(net26),
    .B2(_1107_),
    .X(_1213_));
 sky130_fd_sc_hd__nor2_1 _1935_ (.A(_0834_),
    .B(_0937_),
    .Y(_1214_));
 sky130_fd_sc_hd__a32o_1 _1936_ (.A1(_1072_),
    .A2(_1086_),
    .A3(_1111_),
    .B1(_1214_),
    .B2(_1032_),
    .X(_1215_));
 sky130_fd_sc_hd__or3_1 _1937_ (.A(_0826_),
    .B(_0834_),
    .C(_0979_),
    .X(_1216_));
 sky130_fd_sc_hd__or4b_1 _1938_ (.A(_1100_),
    .B(_1213_),
    .C(_1215_),
    .D_N(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__or4_1 _1939_ (.A(_1124_),
    .B(_1132_),
    .C(_1174_),
    .D(_1193_),
    .X(_1218_));
 sky130_fd_sc_hd__or4_1 _1940_ (.A(_1208_),
    .B(_1211_),
    .C(_1217_),
    .D(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__or4_1 _1941_ (.A(_1166_),
    .B(_1190_),
    .C(_1204_),
    .D(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _1942_ (.A(_1220_),
    .X(_0023_));
 sky130_fd_sc_hd__or4_1 _1943_ (.A(_1114_),
    .B(_1142_),
    .C(_1161_),
    .D(_1167_),
    .X(_1221_));
 sky130_fd_sc_hd__or4_1 _1944_ (.A(_1081_),
    .B(_1128_),
    .C(_1132_),
    .D(_1150_),
    .X(_1222_));
 sky130_fd_sc_hd__or4_1 _1945_ (.A(_1095_),
    .B(_1104_),
    .C(_1123_),
    .D(_1210_),
    .X(_1223_));
 sky130_fd_sc_hd__or4_1 _1946_ (.A(_1170_),
    .B(_1178_),
    .C(_1189_),
    .D(_1203_),
    .X(_1224_));
 sky130_fd_sc_hd__or4_1 _1947_ (.A(_1221_),
    .B(_1222_),
    .C(_1223_),
    .D(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__nor2_1 _1948_ (.A(_0937_),
    .B(_0925_),
    .Y(_1226_));
 sky130_fd_sc_hd__a22o_1 _1949_ (.A1(_1226_),
    .A2(_1033_),
    .B1(_1055_),
    .B2(_1111_),
    .X(_1227_));
 sky130_fd_sc_hd__or4_1 _1950_ (.A(_1088_),
    .B(_1112_),
    .C(_1202_),
    .D(_1215_),
    .X(_1228_));
 sky130_fd_sc_hd__a32o_1 _1951_ (.A1(_1038_),
    .A2(_1072_),
    .A3(_1085_),
    .B1(_1034_),
    .B2(_0926_),
    .X(_1229_));
 sky130_fd_sc_hd__or4_1 _1952_ (.A(_1199_),
    .B(_1227_),
    .C(_1228_),
    .D(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__or2_1 _1953_ (.A(_1225_),
    .B(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _1954_ (.A(_1231_),
    .X(_0024_));
 sky130_fd_sc_hd__a211o_1 _1955_ (.A1(_0943_),
    .A2(_1034_),
    .B1(_1143_),
    .C1(_1149_),
    .X(_1232_));
 sky130_fd_sc_hd__o2111a_1 _1956_ (.A1(net4),
    .A2(_1093_),
    .B1(_1018_),
    .C1(_1025_),
    .D1(net3),
    .X(_1233_));
 sky130_fd_sc_hd__a31o_1 _1957_ (.A1(_1051_),
    .A2(_1056_),
    .A3(_1103_),
    .B1(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__a21o_1 _1958_ (.A1(_1038_),
    .A2(_1234_),
    .B1(_1213_),
    .X(_1235_));
 sky130_fd_sc_hd__or4_1 _1959_ (.A(_1155_),
    .B(_1159_),
    .C(_1177_),
    .D(_1187_),
    .X(_1236_));
 sky130_fd_sc_hd__or4_1 _1960_ (.A(_1181_),
    .B(_1198_),
    .C(_1235_),
    .D(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__or4_1 _1961_ (.A(_1083_),
    .B(_1095_),
    .C(_1232_),
    .D(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__or4_1 _1962_ (.A(_1101_),
    .B(_1122_),
    .C(_1201_),
    .D(_1227_),
    .X(_1239_));
 sky130_fd_sc_hd__or2_1 _1963_ (.A(_1133_),
    .B(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__or4_1 _1964_ (.A(_1109_),
    .B(_1126_),
    .C(_1165_),
    .D(_1168_),
    .X(_1241_));
 sky130_fd_sc_hd__or4_1 _1965_ (.A(_1185_),
    .B(_1194_),
    .C(_1228_),
    .D(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__or3_1 _1966_ (.A(_1238_),
    .B(_1240_),
    .C(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _1967_ (.A(_1243_),
    .X(_0025_));
 sky130_fd_sc_hd__and2b_1 _1968_ (.A_N(\top8227.pulse_slower.currentEnableState[1] ),
    .B(net64),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _1969_ (.A(_1244_),
    .X(\top8227.pulse_slower.nextEnableState[1] ));
 sky130_fd_sc_hd__inv_2 _1970_ (.A(gpio[17]),
    .Y(\top8227.instructionLoader.interruptInjector.interruptRequest ));
 sky130_fd_sc_hd__inv_2 _1971_ (.A(gpio[16]),
    .Y(\top8227.instructionLoader.interruptInjector.nmiSync.in ));
 sky130_fd_sc_hd__clkbuf_4 _1972_ (.A(_0972_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_4 _1973_ (.A(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__buf_4 _1974_ (.A(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__and3_2 _1975_ (.A(_1002_),
    .B(_0903_),
    .C(_0854_),
    .X(_1248_));
 sky130_fd_sc_hd__o211a_1 _1976_ (.A1(_0894_),
    .A2(_0854_),
    .B1(_1084_),
    .C1(_0908_),
    .X(_1249_));
 sky130_fd_sc_hd__a21oi_1 _1977_ (.A1(_0839_),
    .A2(_0846_),
    .B1(_0928_),
    .Y(_1250_));
 sky130_fd_sc_hd__and2_2 _1978_ (.A(_0908_),
    .B(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__or3_1 _1979_ (.A(_1248_),
    .B(_1249_),
    .C(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__o31a_1 _1980_ (.A1(_0877_),
    .A2(_1212_),
    .A3(_1151_),
    .B1(_1003_),
    .X(_1253_));
 sky130_fd_sc_hd__or2_1 _1981_ (.A(_1195_),
    .B(_1135_),
    .X(_1254_));
 sky130_fd_sc_hd__o21a_1 _1982_ (.A1(_1254_),
    .A2(_0923_),
    .B1(_1004_),
    .X(_1255_));
 sky130_fd_sc_hd__o21a_1 _1983_ (.A1(_0872_),
    .A2(_1158_),
    .B1(_1005_),
    .X(_1256_));
 sky130_fd_sc_hd__or4_1 _1984_ (.A(_1252_),
    .B(_1253_),
    .C(_1255_),
    .D(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__and2_1 _1985_ (.A(_0907_),
    .B(_1158_),
    .X(_1258_));
 sky130_fd_sc_hd__nor2_1 _1986_ (.A(_1248_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_2 _1987_ (.A(_1078_),
    .B(_0985_),
    .Y(_1260_));
 sky130_fd_sc_hd__or3b_4 _1988_ (.A(_1259_),
    .B(_1260_),
    .C_N(\top8227.PSRCurrentValue[3] ),
    .X(_1261_));
 sky130_fd_sc_hd__nor2_2 _1989_ (.A(_0907_),
    .B(_0957_),
    .Y(_1262_));
 sky130_fd_sc_hd__or2_2 _1990_ (.A(\top8227.demux.state_machine.currentAddress[10] ),
    .B(\top8227.demux.state_machine.currentAddress[4] ),
    .X(_1263_));
 sky130_fd_sc_hd__a21o_1 _1991_ (.A1(_1262_),
    .A2(_1263_),
    .B1(_1078_),
    .X(_1264_));
 sky130_fd_sc_hd__a21o_2 _1992_ (.A1(_0957_),
    .A2(_0815_),
    .B1(_0908_),
    .X(_1265_));
 sky130_fd_sc_hd__or2_1 _1993_ (.A(_0987_),
    .B(\top8227.demux.state_machine.currentAddress[6] ),
    .X(_1266_));
 sky130_fd_sc_hd__clkinv_4 _1994_ (.A(\top8227.demux.state_machine.timeState[0] ),
    .Y(_1267_));
 sky130_fd_sc_hd__and3_1 _1995_ (.A(_1267_),
    .B(\top8227.demux.state_machine.currentAddress[12] ),
    .C(_0965_),
    .X(_1268_));
 sky130_fd_sc_hd__a221o_1 _1996_ (.A1(_1004_),
    .A2(_1016_),
    .B1(_1265_),
    .B2(_1266_),
    .C1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__a31oi_4 _1997_ (.A1(_0837_),
    .A2(_0844_),
    .A3(_0858_),
    .B1(_0957_),
    .Y(_1270_));
 sky130_fd_sc_hd__and2_1 _1998_ (.A(\top8227.branchForward ),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__o21a_1 _1999_ (.A1(_1127_),
    .A2(_0887_),
    .B1(_1004_),
    .X(_1272_));
 sky130_fd_sc_hd__nand2_2 _2000_ (.A(_0960_),
    .B(_0990_),
    .Y(_1273_));
 sky130_fd_sc_hd__or2_2 _2001_ (.A(_0908_),
    .B(_0815_),
    .X(_1274_));
 sky130_fd_sc_hd__or2_2 _2002_ (.A(_0819_),
    .B(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__and2_1 _2003_ (.A(_0914_),
    .B(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__a211o_1 _2004_ (.A1(_1184_),
    .A2(_1273_),
    .B1(_1276_),
    .C1(_0982_),
    .X(_1277_));
 sky130_fd_sc_hd__and3_1 _2005_ (.A(\top8227.demux.state_machine.timeState[1] ),
    .B(_0849_),
    .C(_0894_),
    .X(_1278_));
 sky130_fd_sc_hd__and3_1 _2006_ (.A(_1003_),
    .B(_0894_),
    .C(_0901_),
    .X(_1279_));
 sky130_fd_sc_hd__or2_1 _2007_ (.A(_1278_),
    .B(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__a21oi_1 _2008_ (.A1(_0839_),
    .A2(_0846_),
    .B1(_0879_),
    .Y(_1281_));
 sky130_fd_sc_hd__and2_1 _2009_ (.A(_1003_),
    .B(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__or4_1 _2010_ (.A(_1272_),
    .B(_1277_),
    .C(_1280_),
    .D(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__o22a_1 _2011_ (.A1(_1264_),
    .A2(_1269_),
    .B1(_1271_),
    .B2(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__and2_1 _2012_ (.A(\top8227.branchBackward ),
    .B(_1270_),
    .X(_1285_));
 sky130_fd_sc_hd__o21a_1 _2013_ (.A1(_0923_),
    .A2(_0950_),
    .B1(_1003_),
    .X(_1286_));
 sky130_fd_sc_hd__o21a_1 _2014_ (.A1(_1209_),
    .A2(_0949_),
    .B1(_1002_),
    .X(_1287_));
 sky130_fd_sc_hd__and2_1 _2015_ (.A(_1096_),
    .B(_1275_),
    .X(_1288_));
 sky130_fd_sc_hd__o21a_1 _2016_ (.A1(_0955_),
    .A2(_1013_),
    .B1(_1127_),
    .X(_1289_));
 sky130_fd_sc_hd__or4_1 _2017_ (.A(_0981_),
    .B(_1287_),
    .C(_1288_),
    .D(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__a21oi_4 _2018_ (.A1(_0830_),
    .A2(_0842_),
    .B1(_0879_),
    .Y(_1291_));
 sky130_fd_sc_hd__o21a_1 _2019_ (.A1(_1254_),
    .A2(_1291_),
    .B1(_1003_),
    .X(_1292_));
 sky130_fd_sc_hd__or4_1 _2020_ (.A(_1253_),
    .B(_1286_),
    .C(_1290_),
    .D(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__nor2_2 _2021_ (.A(_0883_),
    .B(_0936_),
    .Y(_1294_));
 sky130_fd_sc_hd__a31oi_4 _2022_ (.A1(_0871_),
    .A2(_0876_),
    .A3(_0920_),
    .B1(_0825_),
    .Y(_1295_));
 sky130_fd_sc_hd__and2_2 _2023_ (.A(_1003_),
    .B(_0891_),
    .X(_1296_));
 sky130_fd_sc_hd__a221o_1 _2024_ (.A1(_0955_),
    .A2(_1294_),
    .B1(_1295_),
    .B2(_1003_),
    .C1(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__and2_2 _2025_ (.A(_1003_),
    .B(_0868_),
    .X(_1298_));
 sky130_fd_sc_hd__or3_1 _2026_ (.A(_1252_),
    .B(_1297_),
    .C(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__or3_1 _2027_ (.A(_1285_),
    .B(_1293_),
    .C(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__or2_2 _2028_ (.A(\top8227.demux.state_machine.currentAddress[3] ),
    .B(\top8227.demux.state_machine.currentAddress[11] ),
    .X(_1301_));
 sky130_fd_sc_hd__or4_1 _2029_ (.A(\top8227.demux.state_machine.currentAddress[12] ),
    .B(\top8227.demux.state_machine.currentAddress[10] ),
    .C(\top8227.demux.state_machine.currentAddress[4] ),
    .D(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__a221o_1 _2030_ (.A1(_0987_),
    .A2(_1262_),
    .B1(_1302_),
    .B2(_1004_),
    .C1(_1078_),
    .X(_1303_));
 sky130_fd_sc_hd__and4b_1 _2031_ (.A_N(_1284_),
    .B(_0985_),
    .C(_1300_),
    .D(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__buf_2 _2032_ (.A(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__o21a_1 _2033_ (.A1(_0912_),
    .A2(_1120_),
    .B1(_1001_),
    .X(_1306_));
 sky130_fd_sc_hd__nor2_1 _2034_ (.A(_1285_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__or4_1 _2035_ (.A(_0877_),
    .B(_0943_),
    .C(_0944_),
    .D(_0952_),
    .X(_1308_));
 sky130_fd_sc_hd__and2_1 _2036_ (.A(_0815_),
    .B(_0884_),
    .X(_1309_));
 sky130_fd_sc_hd__o21a_1 _2037_ (.A1(_0872_),
    .A2(_0881_),
    .B1(_1002_),
    .X(_1310_));
 sky130_fd_sc_hd__a211o_1 _2038_ (.A1(_1002_),
    .A2(_1308_),
    .B1(_1309_),
    .C1(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__o21ai_4 _2039_ (.A1(_1298_),
    .A2(_1311_),
    .B1(_0972_),
    .Y(_1312_));
 sky130_fd_sc_hd__a21oi_1 _2040_ (.A1(\top8227.demux.state_machine.currentAddress[12] ),
    .A2(_1262_),
    .B1(_0971_),
    .Y(_1313_));
 sky130_fd_sc_hd__o21ai_1 _2041_ (.A1(_0908_),
    .A2(_0994_),
    .B1(_0997_),
    .Y(_1314_));
 sky130_fd_sc_hd__o21ai_2 _2042_ (.A1(_1175_),
    .A2(_1090_),
    .B1(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__or2_1 _2043_ (.A(_0907_),
    .B(\top8227.demux.state_machine.timeState[4] ),
    .X(_1316_));
 sky130_fd_sc_hd__clkbuf_4 _2044_ (.A(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__o31a_1 _2045_ (.A1(_0941_),
    .A2(_0949_),
    .A3(_1291_),
    .B1(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__o41a_1 _2046_ (.A1(_1146_),
    .A2(_1151_),
    .A3(_0891_),
    .A4(_1318_),
    .B1(_0955_),
    .X(_1319_));
 sky130_fd_sc_hd__o21a_1 _2047_ (.A1(_0923_),
    .A2(_0950_),
    .B1(_0818_),
    .X(_1320_));
 sky130_fd_sc_hd__and4b_4 _2048_ (.A_N(_0852_),
    .B(_0853_),
    .C(_0903_),
    .D(_0850_),
    .X(_1321_));
 sky130_fd_sc_hd__and2_1 _2049_ (.A(_0993_),
    .B(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__o41a_1 _2050_ (.A1(_0902_),
    .A2(_0947_),
    .A3(_1320_),
    .A4(_1322_),
    .B1(_1317_),
    .X(_1323_));
 sky130_fd_sc_hd__and2_1 _2051_ (.A(_1001_),
    .B(_0887_),
    .X(_1324_));
 sky130_fd_sc_hd__a31oi_2 _2052_ (.A1(_0876_),
    .A2(_0834_),
    .A3(_0865_),
    .B1(_0883_),
    .Y(_1325_));
 sky130_fd_sc_hd__a21o_1 _2053_ (.A1(_0818_),
    .A2(_1325_),
    .B1(_0980_),
    .X(_1326_));
 sky130_fd_sc_hd__o21a_1 _2054_ (.A1(_0850_),
    .A2(_0851_),
    .B1(_0933_),
    .X(_1327_));
 sky130_fd_sc_hd__o31a_1 _2055_ (.A1(_0934_),
    .A2(_1295_),
    .A3(_1327_),
    .B1(_0818_),
    .X(_1328_));
 sky130_fd_sc_hd__or4_1 _2056_ (.A(_1323_),
    .B(_1324_),
    .C(_1326_),
    .D(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__nor2_1 _2057_ (.A(_1319_),
    .B(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__a211o_4 _2058_ (.A1(_1313_),
    .A2(_1315_),
    .B1(_1330_),
    .C1(_0976_),
    .X(_1331_));
 sky130_fd_sc_hd__and2b_1 _2059_ (.A_N(_1312_),
    .B(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_4 _2060_ (.A(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__or2_1 _2061_ (.A(_1285_),
    .B(_1306_),
    .X(_1334_));
 sky130_fd_sc_hd__or2_2 _2062_ (.A(\top8227.branchBackward ),
    .B(\top8227.branchForward ),
    .X(_1335_));
 sky130_fd_sc_hd__a31oi_2 _2063_ (.A1(_1014_),
    .A2(_0868_),
    .A3(_1335_),
    .B1(_0981_),
    .Y(_1336_));
 sky130_fd_sc_hd__inv_2 _2064_ (.A(\top8227.demux.state_machine.currentAddress[1] ),
    .Y(_1337_));
 sky130_fd_sc_hd__o22ai_2 _2065_ (.A1(_0995_),
    .A2(_0996_),
    .B1(_0992_),
    .B2(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__nor2_1 _2066_ (.A(_1078_),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__or3_1 _2067_ (.A(_0976_),
    .B(_1336_),
    .C(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__and4_1 _2068_ (.A(_0972_),
    .B(_1312_),
    .C(_1334_),
    .D(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_4 _2069_ (.A(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__a21oi_4 _2070_ (.A1(_1307_),
    .A2(_1333_),
    .B1(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__o41a_1 _2071_ (.A1(_0941_),
    .A2(_0949_),
    .A3(_1291_),
    .A4(_1281_),
    .B1(_0818_),
    .X(_1344_));
 sky130_fd_sc_hd__or2_1 _2072_ (.A(_1320_),
    .B(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__and2b_1 _2073_ (.A_N(_0853_),
    .B(_0852_),
    .X(_1346_));
 sky130_fd_sc_hd__and4_1 _2074_ (.A(_0850_),
    .B(\top8227.demux.state_machine.timeState[4] ),
    .C(_0903_),
    .D(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a221o_1 _2075_ (.A1(_0814_),
    .A2(_0889_),
    .B1(_0915_),
    .B2(\top8227.demux.state_machine.timeState[6] ),
    .C1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__o311a_1 _2076_ (.A1(\top8227.demux.state_machine.timeState[4] ),
    .A2(\top8227.demux.state_machine.timeState[6] ),
    .A3(\top8227.demux.state_machine.timeState[1] ),
    .B1(_0901_),
    .C1(_0856_),
    .X(_1349_));
 sky130_fd_sc_hd__a221o_1 _2077_ (.A1(_0814_),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\top8227.demux.state_machine.timeState[4] ),
    .C1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__o21a_1 _2078_ (.A1(_1151_),
    .A2(_0902_),
    .B1(\top8227.demux.state_machine.timeState[4] ),
    .X(_1351_));
 sky130_fd_sc_hd__a22oi_1 _2079_ (.A1(_0859_),
    .A2(_0896_),
    .B1(_0914_),
    .B2(_0814_),
    .Y(_1352_));
 sky130_fd_sc_hd__or4b_1 _2080_ (.A(_1348_),
    .B(_1350_),
    .C(_1351_),
    .D_N(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__a311o_1 _2081_ (.A1(_0814_),
    .A2(_0868_),
    .A3(_1335_),
    .B1(_1326_),
    .C1(_1328_),
    .X(_1354_));
 sky130_fd_sc_hd__inv_2 _2082_ (.A(_1313_),
    .Y(_1355_));
 sky130_fd_sc_hd__o32a_1 _2083_ (.A1(_1345_),
    .A2(_1353_),
    .A3(_1354_),
    .B1(_1338_),
    .B2(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__a21bo_1 _2084_ (.A1(_0908_),
    .A2(_0884_),
    .B1_N(_0958_),
    .X(_1357_));
 sky130_fd_sc_hd__o31a_1 _2085_ (.A1(_0886_),
    .A2(_0932_),
    .A3(_1321_),
    .B1(_0908_),
    .X(_1358_));
 sky130_fd_sc_hd__nor2_1 _2086_ (.A(_1357_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__inv_2 _2087_ (.A(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__a32o_2 _2088_ (.A1(\top8227.pulse_slower.nextEnableState[0] ),
    .A2(_0974_),
    .A3(_1356_),
    .B1(_1360_),
    .B2(_0972_),
    .X(_1361_));
 sky130_fd_sc_hd__o41a_1 _2089_ (.A1(_0902_),
    .A2(_1131_),
    .A3(_1195_),
    .A4(_0949_),
    .B1(_0993_),
    .X(_1362_));
 sky130_fd_sc_hd__o311a_1 _2090_ (.A1(_0908_),
    .A2(\top8227.demux.state_machine.currentAddress[1] ),
    .A3(_1090_),
    .B1(_1317_),
    .C1(_0980_),
    .X(_1363_));
 sky130_fd_sc_hd__or4_1 _2091_ (.A(_0907_),
    .B(\top8227.demux.state_machine.currentAddress[1] ),
    .C(_1016_),
    .D(\top8227.demux.state_machine.currentAddress[11] ),
    .X(_1364_));
 sky130_fd_sc_hd__a211o_1 _2092_ (.A1(\top8227.demux.state_machine.currentAddress[5] ),
    .A2(_1090_),
    .B1(\top8227.demux.state_machine.currentAddress[10] ),
    .C1(_1267_),
    .X(_1365_));
 sky130_fd_sc_hd__a211o_1 _2093_ (.A1(_1364_),
    .A2(_1365_),
    .B1(\top8227.demux.state_machine.currentAddress[3] ),
    .C1(_0971_),
    .X(_1366_));
 sky130_fd_sc_hd__o21ai_1 _2094_ (.A1(_1362_),
    .A2(_1363_),
    .B1(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__or3_2 _2095_ (.A(_0969_),
    .B(_0983_),
    .C(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__o41a_1 _2096_ (.A1(_1110_),
    .A2(_1135_),
    .A3(_0948_),
    .A4(_1214_),
    .B1(_0993_),
    .X(_1369_));
 sky130_fd_sc_hd__or4_1 _2097_ (.A(\top8227.demux.state_machine.currentAddress[11] ),
    .B(\top8227.demux.state_machine.currentAddress[12] ),
    .C(\top8227.demux.state_machine.currentAddress[4] ),
    .D(_0971_),
    .X(_1370_));
 sky130_fd_sc_hd__a22o_1 _2098_ (.A1(_1175_),
    .A2(_1314_),
    .B1(_1370_),
    .B2(_0993_),
    .X(_1371_));
 sky130_fd_sc_hd__o21ai_1 _2099_ (.A1(_0981_),
    .A2(_1369_),
    .B1(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__or3_2 _2100_ (.A(_0969_),
    .B(_0983_),
    .C(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__o31a_1 _2101_ (.A1(_0891_),
    .A2(_0923_),
    .A3(_0951_),
    .B1(_0993_),
    .X(_1374_));
 sky130_fd_sc_hd__o21a_1 _2102_ (.A1(_1209_),
    .A2(_0938_),
    .B1(_0993_),
    .X(_1375_));
 sky130_fd_sc_hd__o21a_1 _2103_ (.A1(_1179_),
    .A2(_0950_),
    .B1(_0908_),
    .X(_1376_));
 sky130_fd_sc_hd__or4_2 _2104_ (.A(_1249_),
    .B(_1251_),
    .C(_1258_),
    .D(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__o41ai_4 _2105_ (.A1(_1374_),
    .A2(_1360_),
    .A3(_1375_),
    .A4(_1377_),
    .B1(_0972_),
    .Y(_1378_));
 sky130_fd_sc_hd__and4bb_1 _2106_ (.A_N(_1361_),
    .B_N(_1368_),
    .C(_1373_),
    .D(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_4 _2107_ (.A(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__a21oi_2 _2108_ (.A1(_1373_),
    .A2(_1378_),
    .B1(_1361_),
    .Y(_1381_));
 sky130_fd_sc_hd__and3_1 _2109_ (.A(_1373_),
    .B(_1361_),
    .C(_1368_),
    .X(_1382_));
 sky130_fd_sc_hd__or3_1 _2110_ (.A(_1380_),
    .B(_1381_),
    .C(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__buf_4 _2111_ (.A(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__and4bb_1 _2112_ (.A_N(_1378_),
    .B_N(_1361_),
    .C(_1368_),
    .D(_1373_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_4 _2113_ (.A(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__nand2_1 _2114_ (.A(_1373_),
    .B(_1368_),
    .Y(_1387_));
 sky130_fd_sc_hd__and2_2 _2115_ (.A(_1387_),
    .B(_1381_),
    .X(_1388_));
 sky130_fd_sc_hd__and4b_1 _2116_ (.A_N(_1378_),
    .B(_1361_),
    .C(_1368_),
    .D(_1373_),
    .X(_1389_));
 sky130_fd_sc_hd__buf_2 _2117_ (.A(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__and4_4 _2118_ (.A(_1373_),
    .B(_1378_),
    .C(_1361_),
    .D(_1368_),
    .X(_1391_));
 sky130_fd_sc_hd__a22o_1 _2119_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[38] ),
    .A2(_1390_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[30] ),
    .X(_1392_));
 sky130_fd_sc_hd__a221o_1 _2120_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[38] ),
    .A2(_1380_),
    .B1(_1388_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[46] ),
    .C1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__a21oi_1 _2121_ (.A1(\top8227.internalDataflow.accRegToDB[6] ),
    .A2(_1386_),
    .B1(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__a2111oi_1 _2122_ (.A1(_0972_),
    .A2(_1288_),
    .B1(_1380_),
    .C1(_1381_),
    .D1(_1382_),
    .Y(_1395_));
 sky130_fd_sc_hd__a21oi_2 _2123_ (.A1(_1384_),
    .A2(_1394_),
    .B1(net20),
    .Y(_1396_));
 sky130_fd_sc_hd__nor2_1 _2124_ (.A(_0872_),
    .B(_0877_),
    .Y(_1397_));
 sky130_fd_sc_hd__a2111o_1 _2125_ (.A1(_0819_),
    .A2(_0927_),
    .B1(_0945_),
    .C1(_0891_),
    .D1(_0923_),
    .X(_1398_));
 sky130_fd_sc_hd__a2bb2o_1 _2126_ (.A1_N(_0960_),
    .A2_N(_1397_),
    .B1(_1317_),
    .B2(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__or2_2 _2127_ (.A(_0814_),
    .B(_0859_),
    .X(_1400_));
 sky130_fd_sc_hd__a311oi_1 _2128_ (.A1(_0846_),
    .A2(_0842_),
    .A3(_0885_),
    .B1(_0911_),
    .C1(_0957_),
    .Y(_1401_));
 sky130_fd_sc_hd__a221o_1 _2129_ (.A1(_1400_),
    .A2(_0880_),
    .B1(_0941_),
    .B2(_1316_),
    .C1(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__or2_1 _2130_ (.A(_0936_),
    .B(_0928_),
    .X(_1403_));
 sky130_fd_sc_hd__a311o_1 _2131_ (.A1(_0871_),
    .A2(_0925_),
    .A3(_0920_),
    .B1(_0928_),
    .C1(_1267_),
    .X(_1404_));
 sky130_fd_sc_hd__a32o_1 _2132_ (.A1(_0929_),
    .A2(_0939_),
    .A3(_1403_),
    .B1(_1404_),
    .B2(_0957_),
    .X(_1405_));
 sky130_fd_sc_hd__or2b_1 _2133_ (.A(_1402_),
    .B_N(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__o41a_1 _2134_ (.A1(_0931_),
    .A2(_0932_),
    .A3(_0933_),
    .A4(_0934_),
    .B1(_0818_),
    .X(_1407_));
 sky130_fd_sc_hd__a221o_1 _2135_ (.A1(_1294_),
    .A2(_0965_),
    .B1(_0884_),
    .B2(_1400_),
    .C1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__or2_1 _2136_ (.A(_1406_),
    .B(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__a22o_1 _2137_ (.A1(_1400_),
    .A2(_1151_),
    .B1(_0952_),
    .B2(_1316_),
    .X(_1410_));
 sky130_fd_sc_hd__a21oi_2 _2138_ (.A1(_0834_),
    .A2(_0885_),
    .B1(_0883_),
    .Y(_1411_));
 sky130_fd_sc_hd__and2_1 _2139_ (.A(_1400_),
    .B(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__a2111o_1 _2140_ (.A1(_0819_),
    .A2(_0906_),
    .B1(_1410_),
    .C1(_1412_),
    .D1(_0909_),
    .X(_1413_));
 sky130_fd_sc_hd__o21a_1 _2141_ (.A1(\top8227.demux.state_machine.timeState[1] ),
    .A2(\top8227.demux.state_machine.timeState[5] ),
    .B1(_0914_),
    .X(_1414_));
 sky130_fd_sc_hd__o21a_1 _2142_ (.A1(_0859_),
    .A2(\top8227.demux.state_machine.timeState[5] ),
    .B1(_0912_),
    .X(_1415_));
 sky130_fd_sc_hd__a221o_1 _2143_ (.A1(\top8227.demux.state_machine.timeState[5] ),
    .A2(_0915_),
    .B1(_0951_),
    .B2(_1317_),
    .C1(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__or4_1 _2144_ (.A(_0981_),
    .B(_0899_),
    .C(_1414_),
    .D(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__nor4_1 _2145_ (.A(_1399_),
    .B(_1409_),
    .C(_1413_),
    .D(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand2_1 _2146_ (.A(_0950_),
    .B(_1317_),
    .Y(_1419_));
 sky130_fd_sc_hd__or3_1 _2147_ (.A(_1001_),
    .B(_0955_),
    .C(_0859_),
    .X(_1420_));
 sky130_fd_sc_hd__o21ai_1 _2148_ (.A1(_0817_),
    .A2(_1420_),
    .B1(_0868_),
    .Y(_1421_));
 sky130_fd_sc_hd__a21oi_2 _2149_ (.A1(_1001_),
    .A2(_1263_),
    .B1(_0971_),
    .Y(_1422_));
 sky130_fd_sc_hd__a21bo_1 _2150_ (.A1(_1001_),
    .A2(_1016_),
    .B1_N(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__a21oi_1 _2151_ (.A1(\top8227.demux.state_machine.currentAddress[6] ),
    .A2(_1265_),
    .B1(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__a311o_1 _2152_ (.A1(net28),
    .A2(_1419_),
    .A3(_1421_),
    .B1(_1424_),
    .C1(_0975_),
    .X(_1425_));
 sky130_fd_sc_hd__o21a_1 _2153_ (.A1(_0912_),
    .A2(_0915_),
    .B1(\top8227.demux.state_machine.timeState[1] ),
    .X(_1426_));
 sky130_fd_sc_hd__a221o_1 _2154_ (.A1(_0916_),
    .A2(_0896_),
    .B1(_0914_),
    .B2(_1013_),
    .C1(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__o21a_1 _2155_ (.A1(_0819_),
    .A2(_0991_),
    .B1(\top8227.demux.state_machine.currentAddress[6] ),
    .X(_1428_));
 sky130_fd_sc_hd__and2_1 _2156_ (.A(_1267_),
    .B(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__a32o_1 _2157_ (.A1(\top8227.demux.state_machine.currentAddress[12] ),
    .A2(_0990_),
    .A3(_0991_),
    .B1(_1262_),
    .B2(_1016_),
    .X(_1430_));
 sky130_fd_sc_hd__or3_1 _2158_ (.A(_1078_),
    .B(_1429_),
    .C(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__o31a_1 _2159_ (.A1(_0981_),
    .A2(_1306_),
    .A3(_1427_),
    .B1(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__and3_1 _2160_ (.A(_0985_),
    .B(_1425_),
    .C(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__buf_2 _2161_ (.A(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__a21oi_4 _2162_ (.A1(_0985_),
    .A2(_1432_),
    .B1(_1425_),
    .Y(_1435_));
 sky130_fd_sc_hd__o21a_1 _2163_ (.A1(_1127_),
    .A2(_0887_),
    .B1(_0955_),
    .X(_1436_));
 sky130_fd_sc_hd__o21a_1 _2164_ (.A1(_1294_),
    .A2(_0896_),
    .B1(_1002_),
    .X(_1437_));
 sky130_fd_sc_hd__or3_1 _2165_ (.A(_1322_),
    .B(_1436_),
    .C(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__o211ai_2 _2166_ (.A1(_1013_),
    .A2(_1009_),
    .B1(_1096_),
    .C1(_1245_),
    .Y(_1439_));
 sky130_fd_sc_hd__nor4_1 _2167_ (.A(_1434_),
    .B(_1435_),
    .C(_1438_),
    .D(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__a221o_1 _2168_ (.A1(net7),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[22] ),
    .C1(net19),
    .X(_1441_));
 sky130_fd_sc_hd__a22o_1 _2169_ (.A1(_1343_),
    .A2(_1396_),
    .B1(_1441_),
    .B2(_1342_),
    .X(_1442_));
 sky130_fd_sc_hd__a22o_1 _2170_ (.A1(_1001_),
    .A2(_0889_),
    .B1(_0896_),
    .B2(_1014_),
    .X(_1443_));
 sky130_fd_sc_hd__a22o_1 _2171_ (.A1(_0819_),
    .A2(_0896_),
    .B1(_0912_),
    .B2(_0815_),
    .X(_1444_));
 sky130_fd_sc_hd__nor2_1 _2172_ (.A(_1443_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _2173_ (.A(\top8227.demux.state_machine.currentAddress[12] ),
    .B(_1265_),
    .Y(_1446_));
 sky130_fd_sc_hd__a21oi_1 _2174_ (.A1(_1263_),
    .A2(_1317_),
    .B1(_0971_),
    .Y(_1447_));
 sky130_fd_sc_hd__or2_1 _2175_ (.A(_1016_),
    .B(_1301_),
    .X(_1448_));
 sky130_fd_sc_hd__a22o_1 _2176_ (.A1(_0993_),
    .A2(_1448_),
    .B1(_1265_),
    .B2(\top8227.demux.state_machine.currentAddress[6] ),
    .X(_1449_));
 sky130_fd_sc_hd__a21oi_1 _2177_ (.A1(_0987_),
    .A2(_1275_),
    .B1(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__and3_1 _2178_ (.A(_1446_),
    .B(_1447_),
    .C(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__or4_1 _2179_ (.A(_1146_),
    .B(_0881_),
    .C(_0941_),
    .D(_1295_),
    .X(_1452_));
 sky130_fd_sc_hd__o31a_1 _2180_ (.A1(_0868_),
    .A2(_1308_),
    .A3(_1452_),
    .B1(_1001_),
    .X(_1453_));
 sky130_fd_sc_hd__a22o_1 _2181_ (.A1(_0815_),
    .A2(_0886_),
    .B1(_0950_),
    .B2(_0993_),
    .X(_1454_));
 sky130_fd_sc_hd__a211o_1 _2182_ (.A1(_0815_),
    .A2(_1321_),
    .B1(_1278_),
    .C1(_0981_),
    .X(_1455_));
 sky130_fd_sc_hd__a2111o_1 _2183_ (.A1(_0859_),
    .A2(_0915_),
    .B1(_1309_),
    .C1(_1454_),
    .D1(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__nor3_1 _2184_ (.A(_1453_),
    .B(_1374_),
    .C(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__o22a_2 _2185_ (.A1(_0981_),
    .A2(_1445_),
    .B1(_1451_),
    .B2(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__o21a_1 _2186_ (.A1(_0896_),
    .A2(_0912_),
    .B1(_1002_),
    .X(_1459_));
 sky130_fd_sc_hd__o31a_1 _2187_ (.A1(_1271_),
    .A2(_1443_),
    .A3(_1459_),
    .B1(_0972_),
    .X(_1460_));
 sky130_fd_sc_hd__o21a_1 _2188_ (.A1(_0890_),
    .A2(_1250_),
    .B1(_1001_),
    .X(_1461_));
 sky130_fd_sc_hd__nor2_1 _2189_ (.A(_1461_),
    .B(_1444_),
    .Y(_1462_));
 sky130_fd_sc_hd__o21ai_1 _2190_ (.A1(_0988_),
    .A2(_0992_),
    .B1(_0998_),
    .Y(_1463_));
 sky130_fd_sc_hd__a21oi_1 _2191_ (.A1(_1226_),
    .A2(_1463_),
    .B1(_1078_),
    .Y(_1464_));
 sky130_fd_sc_hd__a21oi_2 _2192_ (.A1(_1078_),
    .A2(_1462_),
    .B1(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__or3b_1 _2193_ (.A(_0969_),
    .B(_0983_),
    .C_N(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__or2_1 _2194_ (.A(_1460_),
    .B(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__nor2_2 _2195_ (.A(_1458_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__and2_2 _2196_ (.A(_1460_),
    .B(_1458_),
    .X(_1469_));
 sky130_fd_sc_hd__o21a_1 _2197_ (.A1(_0949_),
    .A2(_1291_),
    .B1(_1002_),
    .X(_1470_));
 sky130_fd_sc_hd__a211o_1 _2198_ (.A1(_0955_),
    .A2(_1294_),
    .B1(_1289_),
    .C1(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__o21a_1 _2199_ (.A1(_1285_),
    .A2(_1471_),
    .B1(_0972_),
    .X(_1472_));
 sky130_fd_sc_hd__or3_1 _2200_ (.A(_0975_),
    .B(_1465_),
    .C(_1458_),
    .X(_1473_));
 sky130_fd_sc_hd__and4b_1 _2201_ (.A_N(_1469_),
    .B(_1472_),
    .C(_1467_),
    .D(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__buf_2 _2202_ (.A(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__and4b_4 _2203_ (.A_N(_1458_),
    .B(_1460_),
    .C(_0984_),
    .D(_1466_),
    .X(_1476_));
 sky130_fd_sc_hd__nor4_1 _2204_ (.A(_0976_),
    .B(_1460_),
    .C(_1465_),
    .D(_1458_),
    .Y(_1477_));
 sky130_fd_sc_hd__and3_2 _2205_ (.A(_0985_),
    .B(_1465_),
    .C(_1458_),
    .X(_1478_));
 sky130_fd_sc_hd__a22o_1 _2206_ (.A1(net7),
    .A2(net25),
    .B1(_1478_),
    .B2(\top8227.internalDataflow.accRegToDB[6] ),
    .X(_1479_));
 sky130_fd_sc_hd__a221o_1 _2207_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[22] ),
    .A2(_1469_),
    .B1(_1476_),
    .B2(\top8227.PSRCurrentValue[6] ),
    .C1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__a211o_1 _2208_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[22] ),
    .A2(_1468_),
    .B1(_1475_),
    .C1(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_2 _2209_ (.A0(_1442_),
    .A1(_1481_),
    .S(_1333_),
    .X(_1482_));
 sky130_fd_sc_hd__nand2_1 _2210_ (.A(_1305_),
    .B(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__o21ai_4 _2211_ (.A1(_1248_),
    .A2(_1255_),
    .B1(_1245_),
    .Y(_1484_));
 sky130_fd_sc_hd__a2111oi_2 _2212_ (.A1(_1004_),
    .A2(_0884_),
    .B1(_1287_),
    .C1(_1297_),
    .D1(_1282_),
    .Y(_1485_));
 sky130_fd_sc_hd__or4_1 _2213_ (.A(_1184_),
    .B(_0950_),
    .C(_1291_),
    .D(_1411_),
    .X(_1486_));
 sky130_fd_sc_hd__a211o_1 _2214_ (.A1(_1013_),
    .A2(_1184_),
    .B1(_1289_),
    .C1(_0982_),
    .X(_1487_));
 sky130_fd_sc_hd__a2111o_1 _2215_ (.A1(_0914_),
    .A2(_1274_),
    .B1(_1280_),
    .C1(_1487_),
    .D1(_1251_),
    .X(_1488_));
 sky130_fd_sc_hd__a221oi_2 _2216_ (.A1(_1335_),
    .A2(_1270_),
    .B1(_1486_),
    .B2(_1004_),
    .C1(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__nand2_1 _2217_ (.A(\top8227.demux.state_machine.currentAddress[12] ),
    .B(_1275_),
    .Y(_1490_));
 sky130_fd_sc_hd__a31o_1 _2218_ (.A1(_1447_),
    .A2(_1450_),
    .A3(_1490_),
    .B1(_0976_),
    .X(_1491_));
 sky130_fd_sc_hd__a21o_2 _2219_ (.A1(_1485_),
    .A2(_1489_),
    .B1(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_4 _2220_ (.A(_1331_),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_4 _2221_ (.A0(_1396_),
    .A1(_1481_),
    .S(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _2222_ (.A0(_1484_),
    .A1(_1492_),
    .S(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__o21a_1 _2223_ (.A1(_1002_),
    .A2(_1009_),
    .B1(_1127_),
    .X(_1496_));
 sky130_fd_sc_hd__o21ai_1 _2224_ (.A1(_1437_),
    .A2(_1496_),
    .B1(_0972_),
    .Y(_1497_));
 sky130_fd_sc_hd__nand2_1 _2225_ (.A(_0957_),
    .B(_0960_),
    .Y(_1498_));
 sky130_fd_sc_hd__and3_1 _2226_ (.A(_1267_),
    .B(\top8227.demux.state_machine.currentAddress[12] ),
    .C(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__a32o_1 _2227_ (.A1(_1267_),
    .A2(_0987_),
    .A3(_0965_),
    .B1(_1448_),
    .B2(_1262_),
    .X(_1500_));
 sky130_fd_sc_hd__or4_1 _2228_ (.A(_1264_),
    .B(_1429_),
    .C(_1499_),
    .D(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__o21a_1 _2229_ (.A1(_0916_),
    .A2(_0965_),
    .B1(_0896_),
    .X(_1502_));
 sky130_fd_sc_hd__a221o_1 _2230_ (.A1(_1014_),
    .A2(_0912_),
    .B1(_1184_),
    .B2(_1009_),
    .C1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__a211o_1 _2231_ (.A1(_1498_),
    .A2(_1321_),
    .B1(_1347_),
    .C1(_0981_),
    .X(_1504_));
 sky130_fd_sc_hd__or3_1 _2232_ (.A(_1270_),
    .B(_1503_),
    .C(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__and3_1 _2233_ (.A(_0985_),
    .B(_1501_),
    .C(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__o21ai_1 _2234_ (.A1(_0860_),
    .A2(_1274_),
    .B1(_0868_),
    .Y(_1507_));
 sky130_fd_sc_hd__and2_1 _2235_ (.A(_1419_),
    .B(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__a211oi_2 _2236_ (.A1(net27),
    .A2(_1508_),
    .B1(_0975_),
    .C1(_1424_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor3_1 _2237_ (.A(_1497_),
    .B(_1506_),
    .C(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__o21a_1 _2238_ (.A1(\top8227.demux.state_machine.currentAddress[5] ),
    .A2(_0987_),
    .B1(_1001_),
    .X(_0120_));
 sky130_fd_sc_hd__and4_1 _2239_ (.A(gpio[19]),
    .B(_0981_),
    .C(\top8227.pulse_slower.nextEnableState[0] ),
    .D(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__a31o_1 _2240_ (.A1(_0984_),
    .A2(_1501_),
    .A3(_1505_),
    .B1(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__and2_1 _2241_ (.A(_1497_),
    .B(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__and3b_1 _2242_ (.A_N(_0122_),
    .B(_1497_),
    .C(_0118_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_4 _2243_ (.A(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__nor3_4 _2244_ (.A(_0119_),
    .B(_0123_),
    .C(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__and2_1 _2245_ (.A(_1439_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__nor2_1 _2246_ (.A(_1506_),
    .B(_0118_),
    .Y(_0128_));
 sky130_fd_sc_hd__and2b_1 _2247_ (.A_N(_0128_),
    .B(_0123_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_4 _2248_ (.A(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _2249_ (.A(_0128_),
    .B(_0123_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_4 _2250_ (.A(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__a221o_1 _2251_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[38] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[22] ),
    .C1(_0126_),
    .X(_0133_));
 sky130_fd_sc_hd__a221oi_2 _2252_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[30] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(net7),
    .C1(_0133_),
    .Y(_0134_));
 sky130_fd_sc_hd__or2_2 _2253_ (.A(_0127_),
    .B(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__a221o_1 _2254_ (.A1(_1004_),
    .A2(_1127_),
    .B1(_1184_),
    .B2(_1014_),
    .C1(_1288_),
    .X(_0136_));
 sky130_fd_sc_hd__a211o_1 _2255_ (.A1(_0955_),
    .A2(_1321_),
    .B1(_0136_),
    .C1(_1298_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_1 _2256_ (.A(_1245_),
    .B(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_4 _2257_ (.A(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2258_ (.A0(_1495_),
    .A1(_0135_),
    .S(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__or2_2 _2259_ (.A(_1483_),
    .B(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_1 _2260_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[37] ),
    .A2(_1390_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[29] ),
    .X(_0142_));
 sky130_fd_sc_hd__a221o_1 _2261_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[37] ),
    .A2(_1380_),
    .B1(_1388_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[45] ),
    .C1(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__a21oi_1 _2262_ (.A1(\top8227.internalDataflow.accRegToDB[5] ),
    .A2(_1386_),
    .B1(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__a21oi_2 _2263_ (.A1(_1384_),
    .A2(_0144_),
    .B1(net20),
    .Y(_0145_));
 sky130_fd_sc_hd__a221o_1 _2264_ (.A1(net6),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[21] ),
    .C1(net19),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _2265_ (.A1(_1343_),
    .A2(_0145_),
    .B1(_0146_),
    .B2(_1342_),
    .X(_0147_));
 sky130_fd_sc_hd__a221o_1 _2266_ (.A1(\top8227.internalDataflow.accRegToDB[5] ),
    .A2(_1478_),
    .B1(_1469_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[21] ),
    .C1(_1476_),
    .X(_0148_));
 sky130_fd_sc_hd__a21o_1 _2267_ (.A1(net6),
    .A2(net25),
    .B1(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__a211o_1 _2268_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[21] ),
    .A2(_1468_),
    .B1(_1475_),
    .C1(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_2 _2269_ (.A0(_0147_),
    .A1(_0150_),
    .S(_1333_),
    .X(_0151_));
 sky130_fd_sc_hd__nand2_1 _2270_ (.A(_1305_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__mux2_2 _2271_ (.A0(_0145_),
    .A1(_0150_),
    .S(_1493_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2272_ (.A0(_1484_),
    .A1(_1492_),
    .S(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__and2b_1 _2273_ (.A_N(_0139_),
    .B(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__a221o_1 _2274_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[37] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[21] ),
    .C1(_0126_),
    .X(_0156_));
 sky130_fd_sc_hd__a221oi_2 _2275_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[29] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(net6),
    .C1(_0156_),
    .Y(_0157_));
 sky130_fd_sc_hd__or2_1 _2276_ (.A(_0127_),
    .B(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__buf_2 _2277_ (.A(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _2278_ (.A(_0139_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__or3_4 _2279_ (.A(_0152_),
    .B(_0155_),
    .C(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_1 _2280_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[36] ),
    .A2(_1380_),
    .B1(_1388_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[44] ),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _2281_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[36] ),
    .A2(_1390_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[28] ),
    .X(_0163_));
 sky130_fd_sc_hd__a21bo_1 _2282_ (.A1(\top8227.internalDataflow.accRegToDB[4] ),
    .A2(_1386_),
    .B1_N(_1384_),
    .X(_0164_));
 sky130_fd_sc_hd__a21o_1 _2283_ (.A1(_1245_),
    .A2(_1288_),
    .B1(_1384_),
    .X(_0165_));
 sky130_fd_sc_hd__o31a_1 _2284_ (.A1(_0162_),
    .A2(_0163_),
    .A3(_0164_),
    .B1(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__a221o_1 _2285_ (.A1(net5),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[20] ),
    .C1(net19),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _2286_ (.A1(_1343_),
    .A2(_0166_),
    .B1(_0167_),
    .B2(_1342_),
    .X(_0168_));
 sky130_fd_sc_hd__nor3_1 _2287_ (.A(\top8227.demux.reset ),
    .B(\top8227.demux.nmi ),
    .C(\top8227.demux.setInterruptFlag ),
    .Y(_0169_));
 sky130_fd_sc_hd__a32o_1 _2288_ (.A1(_1014_),
    .A2(_1096_),
    .A3(_0169_),
    .B1(_1294_),
    .B2(_1003_),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _2289_ (.A1(net5),
    .A2(_1477_),
    .B1(_1476_),
    .B2(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__a221o_1 _2290_ (.A1(\top8227.internalDataflow.accRegToDB[4] ),
    .A2(_1478_),
    .B1(_1469_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[20] ),
    .C1(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__a211o_1 _2291_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[20] ),
    .A2(_1468_),
    .B1(_1475_),
    .C1(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_2 _2292_ (.A0(_0168_),
    .A1(_0173_),
    .S(_1333_),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _2293_ (.A(_1305_),
    .B(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__mux2_2 _2294_ (.A0(_0166_),
    .A1(_0173_),
    .S(_1493_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(_1484_),
    .A1(_1492_),
    .S(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a221o_1 _2296_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[36] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[20] ),
    .C1(_0126_),
    .X(_0178_));
 sky130_fd_sc_hd__a221oi_4 _2297_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[28] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(net5),
    .C1(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__or2_4 _2298_ (.A(_0127_),
    .B(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2299_ (.A0(_0177_),
    .A1(_0180_),
    .S(_0139_),
    .X(_0181_));
 sky130_fd_sc_hd__or2_2 _2300_ (.A(_0175_),
    .B(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_1 _2301_ (.A1(\top8227.internalDataflow.accRegToDB[3] ),
    .A2(_1478_),
    .B1(_1476_),
    .B2(\top8227.PSRCurrentValue[3] ),
    .X(_0183_));
 sky130_fd_sc_hd__a221o_1 _2302_ (.A1(net4),
    .A2(net25),
    .B1(_1469_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[19] ),
    .C1(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__a211oi_1 _2303_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[19] ),
    .A2(_1468_),
    .B1(_1475_),
    .C1(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_1 _2304_ (.A(_1331_),
    .B(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__a22o_1 _2305_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[35] ),
    .A2(_1390_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[27] ),
    .X(_0187_));
 sky130_fd_sc_hd__a221o_1 _2306_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[35] ),
    .A2(_1380_),
    .B1(_1388_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[43] ),
    .C1(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__a21bo_1 _2307_ (.A1(\top8227.internalDataflow.accRegToDB[3] ),
    .A2(_1386_),
    .B1_N(_1384_),
    .X(_0189_));
 sky130_fd_sc_hd__o21a_1 _2308_ (.A1(_0188_),
    .A2(_0189_),
    .B1(_0165_),
    .X(_0190_));
 sky130_fd_sc_hd__a221o_1 _2309_ (.A1(net4),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[19] ),
    .C1(net19),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _2310_ (.A1(_1343_),
    .A2(_0190_),
    .B1(_0191_),
    .B2(_1342_),
    .X(_0192_));
 sky130_fd_sc_hd__o22a_2 _2311_ (.A1(_1312_),
    .A2(_0186_),
    .B1(_0192_),
    .B2(_1333_),
    .X(_0193_));
 sky130_fd_sc_hd__and2_1 _2312_ (.A(_1305_),
    .B(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__inv_2 _2313_ (.A(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__o21a_2 _2314_ (.A1(_1493_),
    .A2(_0190_),
    .B1(_0186_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2315_ (.A0(_1484_),
    .A1(_1492_),
    .S(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__a221o_1 _2316_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[35] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[19] ),
    .C1(_0126_),
    .X(_0198_));
 sky130_fd_sc_hd__a221o_1 _2317_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[27] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(net4),
    .C1(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__or2b_1 _2318_ (.A(_0127_),
    .B_N(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__buf_2 _2319_ (.A(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(_0197_),
    .A1(_0201_),
    .S(_0139_),
    .X(_0202_));
 sky130_fd_sc_hd__xnor2_1 _2321_ (.A(_0195_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _2322_ (.A(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__a22o_1 _2323_ (.A1(\top8227.internalDataflow.accRegToDB[2] ),
    .A2(_1478_),
    .B1(_1476_),
    .B2(\top8227.PSRCurrentValue[2] ),
    .X(_0205_));
 sky130_fd_sc_hd__a221o_1 _2324_ (.A1(net3),
    .A2(net25),
    .B1(_1469_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[18] ),
    .C1(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__a211oi_1 _2325_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[18] ),
    .A2(_1468_),
    .B1(_1475_),
    .C1(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _2326_ (.A(_1331_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__a22o_1 _2327_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[34] ),
    .A2(_1390_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[26] ),
    .X(_0209_));
 sky130_fd_sc_hd__a221o_1 _2328_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[34] ),
    .A2(_1380_),
    .B1(_1388_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[42] ),
    .C1(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__a21oi_1 _2329_ (.A1(\top8227.internalDataflow.accRegToDB[2] ),
    .A2(_1386_),
    .B1(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_2 _2330_ (.A1(_1384_),
    .A2(_0211_),
    .B1(net20),
    .Y(_0212_));
 sky130_fd_sc_hd__a221o_1 _2331_ (.A1(net3),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[18] ),
    .C1(net19),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _2332_ (.A1(_1343_),
    .A2(_0212_),
    .B1(_0213_),
    .B2(_1342_),
    .X(_0214_));
 sky130_fd_sc_hd__o22a_2 _2333_ (.A1(_1312_),
    .A2(_0208_),
    .B1(_0214_),
    .B2(_1333_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_2 _2334_ (.A(_1305_),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__o21a_2 _2335_ (.A1(_1331_),
    .A2(_0212_),
    .B1(_0208_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2336_ (.A0(_1484_),
    .A1(_1492_),
    .S(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__o2111ai_2 _2337_ (.A1(_1013_),
    .A2(_1009_),
    .B1(_1096_),
    .C1(_1245_),
    .D1(_0126_),
    .Y(_0219_));
 sky130_fd_sc_hd__a22o_1 _2338_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[34] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[18] ),
    .X(_0220_));
 sky130_fd_sc_hd__a221o_1 _2339_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[26] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(net3),
    .C1(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__o21ba_2 _2340_ (.A1(\top8227.demux.nmi ),
    .A2(_0219_),
    .B1_N(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_2 _2341_ (.A0(_0218_),
    .A1(_0222_),
    .S(_0139_),
    .X(_0223_));
 sky130_fd_sc_hd__xnor2_4 _2342_ (.A(_0216_),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _2343_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[32] ),
    .B(_1390_),
    .Y(_0225_));
 sky130_fd_sc_hd__a22o_1 _2344_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[32] ),
    .A2(_1380_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[24] ),
    .X(_0226_));
 sky130_fd_sc_hd__a221oi_4 _2345_ (.A1(\top8227.internalDataflow.accRegToDB[0] ),
    .A2(_1386_),
    .B1(_1388_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[40] ),
    .C1(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__a21o_1 _2346_ (.A1(_1307_),
    .A2(_1333_),
    .B1(_1342_),
    .X(_0228_));
 sky130_fd_sc_hd__a311oi_1 _2347_ (.A1(_1384_),
    .A2(_0225_),
    .A3(_0227_),
    .B1(_0228_),
    .C1(net21),
    .Y(_0229_));
 sky130_fd_sc_hd__nand2_1 _2348_ (.A(_1245_),
    .B(_1438_),
    .Y(_0230_));
 sky130_fd_sc_hd__a211oi_1 _2349_ (.A1(_0230_),
    .A2(_1439_),
    .B1(_1434_),
    .C1(_1435_),
    .Y(_0231_));
 sky130_fd_sc_hd__a22o_1 _2350_ (.A1(net1),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[16] ),
    .X(_0232_));
 sky130_fd_sc_hd__o21a_1 _2351_ (.A1(_0231_),
    .A2(_0232_),
    .B1(_1342_),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _2352_ (.A1(net1),
    .A2(net25),
    .B1(_1478_),
    .B2(\top8227.internalDataflow.accRegToDB[0] ),
    .X(_0234_));
 sky130_fd_sc_hd__a221o_1 _2353_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[16] ),
    .A2(_1469_),
    .B1(_1476_),
    .B2(\top8227.PSRCurrentValue[0] ),
    .C1(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__a21oi_1 _2354_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[16] ),
    .A2(_1468_),
    .B1(_1475_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand3b_2 _2355_ (.A_N(_0235_),
    .B(_0236_),
    .C(_1331_),
    .Y(_0237_));
 sky130_fd_sc_hd__o32a_2 _2356_ (.A1(_1333_),
    .A2(_0229_),
    .A3(_0233_),
    .B1(_0237_),
    .B2(_1312_),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_1 _2357_ (.A(_1305_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__and4b_1 _2358_ (.A_N(_1013_),
    .B(_1245_),
    .C(_1278_),
    .D(_0126_),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _2359_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[32] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[16] ),
    .X(_0241_));
 sky130_fd_sc_hd__a221o_1 _2360_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[24] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(net1),
    .C1(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_2 _2361_ (.A(_0240_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__or2b_1 _2362_ (.A(_0243_),
    .B_N(_0139_),
    .X(_0244_));
 sky130_fd_sc_hd__a31oi_4 _2363_ (.A1(_1384_),
    .A2(_0225_),
    .A3(_0227_),
    .B1(net21),
    .Y(_0245_));
 sky130_fd_sc_hd__o21ai_1 _2364_ (.A1(_1493_),
    .A2(_0245_),
    .B1(_0237_),
    .Y(_0246_));
 sky130_fd_sc_hd__o211a_1 _2365_ (.A1(_1493_),
    .A2(_0245_),
    .B1(_1492_),
    .C1(_0237_),
    .X(_0247_));
 sky130_fd_sc_hd__a211o_1 _2366_ (.A1(_1484_),
    .A2(_0246_),
    .B1(_0247_),
    .C1(_0139_),
    .X(_0248_));
 sky130_fd_sc_hd__nand3_1 _2367_ (.A(_0239_),
    .B(_0244_),
    .C(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__or2_1 _2368_ (.A(_1248_),
    .B(_1258_),
    .X(_0250_));
 sky130_fd_sc_hd__o31a_1 _2369_ (.A1(_0881_),
    .A2(_0934_),
    .A3(_1186_),
    .B1(_1004_),
    .X(_0251_));
 sky130_fd_sc_hd__o21a_1 _2370_ (.A1(_0250_),
    .A2(_0251_),
    .B1(\top8227.PSRCurrentValue[0] ),
    .X(_0252_));
 sky130_fd_sc_hd__a221o_1 _2371_ (.A1(_0914_),
    .A2(_1317_),
    .B1(_1275_),
    .B2(_1184_),
    .C1(_1279_),
    .X(_0253_));
 sky130_fd_sc_hd__or3_1 _2372_ (.A(_0982_),
    .B(_1255_),
    .C(_1282_),
    .X(_0254_));
 sky130_fd_sc_hd__or4_1 _2373_ (.A(_1324_),
    .B(_0252_),
    .C(_0253_),
    .D(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__a2bb2o_1 _2374_ (.A1_N(_1337_),
    .A2_N(_0996_),
    .B1(_1263_),
    .B2(_1262_),
    .X(_0256_));
 sky130_fd_sc_hd__a221o_1 _2375_ (.A1(_1004_),
    .A2(_0987_),
    .B1(\top8227.freeCarry ),
    .B2(_0256_),
    .C1(_1355_),
    .X(_0257_));
 sky130_fd_sc_hd__o211a_1 _2376_ (.A1(_1271_),
    .A2(_0255_),
    .B1(_0257_),
    .C1(_0985_),
    .X(_0258_));
 sky130_fd_sc_hd__a21oi_1 _2377_ (.A1(_0244_),
    .A2(_0248_),
    .B1(_0239_),
    .Y(_0259_));
 sky130_fd_sc_hd__a21o_2 _2378_ (.A1(_0249_),
    .A2(_0258_),
    .B1(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_1 _2379_ (.A1(\top8227.internalDataflow.accRegToDB[1] ),
    .A2(_1478_),
    .B1(_1476_),
    .B2(\top8227.PSRCurrentValue[1] ),
    .X(_0261_));
 sky130_fd_sc_hd__a221o_1 _2380_ (.A1(net2),
    .A2(net94),
    .B1(_1469_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[17] ),
    .C1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__a211oi_2 _2381_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[17] ),
    .A2(_1468_),
    .B1(_1475_),
    .C1(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _2382_ (.A(_1493_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__a32oi_4 _2383_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[41] ),
    .A2(_1387_),
    .A3(_1381_),
    .B1(_1380_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[33] ),
    .Y(_0265_));
 sky130_fd_sc_hd__a22oi_2 _2384_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[33] ),
    .A2(_1390_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[25] ),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _2385_ (.A(\top8227.internalDataflow.accRegToDB[1] ),
    .B(_1386_),
    .Y(_0267_));
 sky130_fd_sc_hd__a41oi_4 _2386_ (.A1(_1384_),
    .A2(_0265_),
    .A3(_0266_),
    .A4(_0267_),
    .B1(net93),
    .Y(_0268_));
 sky130_fd_sc_hd__a221o_1 _2387_ (.A1(net2),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[17] ),
    .C1(_1440_),
    .X(_0269_));
 sky130_fd_sc_hd__a22o_1 _2388_ (.A1(_1343_),
    .A2(_0268_),
    .B1(_0269_),
    .B2(_1342_),
    .X(_0270_));
 sky130_fd_sc_hd__o22a_2 _2389_ (.A1(_1312_),
    .A2(_0264_),
    .B1(_0270_),
    .B2(_1333_),
    .X(_0271_));
 sky130_fd_sc_hd__and2_2 _2390_ (.A(_1305_),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _2391_ (.A(_1331_),
    .B(_0268_),
    .Y(_0273_));
 sky130_fd_sc_hd__a21oi_2 _2392_ (.A1(_1331_),
    .A2(_0263_),
    .B1(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(_1484_),
    .A1(_1492_),
    .S(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__and2b_1 _2394_ (.A_N(\top8227.demux.nmi ),
    .B(\top8227.demux.reset ),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _2395_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[33] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[17] ),
    .X(_0277_));
 sky130_fd_sc_hd__a221o_1 _2396_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[25] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(net2),
    .C1(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__o21ba_2 _2397_ (.A1(_0219_),
    .A2(_0276_),
    .B1_N(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_2 _2398_ (.A0(_0275_),
    .A1(_0279_),
    .S(_0139_),
    .X(_0280_));
 sky130_fd_sc_hd__xnor2_4 _2399_ (.A(_0272_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand2_1 _2400_ (.A(_1305_),
    .B(_0271_),
    .Y(_0282_));
 sky130_fd_sc_hd__nor2_1 _2401_ (.A(_0282_),
    .B(_0280_),
    .Y(_0283_));
 sky130_fd_sc_hd__a21oi_4 _2402_ (.A1(_0260_),
    .A2(_0281_),
    .B1(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__or2_1 _2403_ (.A(_0216_),
    .B(_0223_),
    .X(_0285_));
 sky130_fd_sc_hd__o21ai_4 _2404_ (.A1(_0224_),
    .A2(_0284_),
    .B1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor2_1 _2405_ (.A(_0195_),
    .B(_0202_),
    .Y(_0287_));
 sky130_fd_sc_hd__a21oi_2 _2406_ (.A1(_0204_),
    .A2(_0286_),
    .B1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__xor2_4 _2407_ (.A(_0224_),
    .B(_0284_),
    .X(_0289_));
 sky130_fd_sc_hd__xnor2_2 _2408_ (.A(_0260_),
    .B(_0281_),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_2 _2409_ (.A(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__o22ai_2 _2410_ (.A1(_0204_),
    .A2(_0286_),
    .B1(_0289_),
    .B2(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__and2_1 _2411_ (.A(_0175_),
    .B(_0181_),
    .X(_0293_));
 sky130_fd_sc_hd__inv_2 _2412_ (.A(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _2413_ (.A(_0182_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__a21o_1 _2414_ (.A1(_0288_),
    .A2(_0292_),
    .B1(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__inv_2 _2415_ (.A(_0161_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21a_1 _2416_ (.A1(_0155_),
    .A2(_0160_),
    .B1(_0152_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_2 _2417_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__a21o_1 _2418_ (.A1(_0182_),
    .A2(_0296_),
    .B1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__and2_1 _2419_ (.A(_1483_),
    .B(_0140_),
    .X(_0301_));
 sky130_fd_sc_hd__inv_2 _2420_ (.A(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _2421_ (.A(_0141_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__a21o_1 _2422_ (.A1(_0161_),
    .A2(_0300_),
    .B1(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__a22o_1 _2423_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[39] ),
    .A2(_1390_),
    .B1(_1391_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[31] ),
    .X(_0305_));
 sky130_fd_sc_hd__a221o_1 _2424_ (.A1(\top8227.internalDataflow.stackBusModule.busInputs[39] ),
    .A2(_1380_),
    .B1(_1388_),
    .B2(\top8227.internalDataflow.stackBusModule.busInputs[47] ),
    .C1(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__a21oi_1 _2425_ (.A1(\top8227.internalDataflow.accRegToDB[7] ),
    .A2(_1386_),
    .B1(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__a21oi_1 _2426_ (.A1(_1384_),
    .A2(_0307_),
    .B1(net20),
    .Y(_0308_));
 sky130_fd_sc_hd__a221o_1 _2427_ (.A1(_1021_),
    .A2(_1434_),
    .B1(_1435_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[23] ),
    .C1(net19),
    .X(_0309_));
 sky130_fd_sc_hd__a22o_1 _2428_ (.A1(_1343_),
    .A2(_0308_),
    .B1(_0309_),
    .B2(_1342_),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _2429_ (.A1(\top8227.internalDataflow.accRegToDB[7] ),
    .A2(_1478_),
    .B1(_1476_),
    .B2(\top8227.PSRCurrentValue[7] ),
    .X(_0311_));
 sky130_fd_sc_hd__a221o_1 _2430_ (.A1(net8),
    .A2(net25),
    .B1(_1469_),
    .B2(\top8227.internalDataflow.addressHighBusModule.busInputs[23] ),
    .C1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a211o_1 _2431_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ),
    .A2(_1468_),
    .B1(_1475_),
    .C1(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_2 _2432_ (.A0(_0310_),
    .A1(_0313_),
    .S(_1333_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _2433_ (.A(_1305_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__mux2_2 _2434_ (.A0(_0308_),
    .A1(_0313_),
    .S(_1493_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(_1484_),
    .A1(_1492_),
    .S(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__a221o_1 _2436_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[39] ),
    .A2(net24),
    .B1(_0125_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ),
    .C1(_0126_),
    .X(_0318_));
 sky130_fd_sc_hd__a221o_1 _2437_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[31] ),
    .A2(_0130_),
    .B1(_0132_),
    .B2(_1021_),
    .C1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__nand2b_4 _2438_ (.A_N(_0127_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(_0317_),
    .A1(_0320_),
    .S(_0139_),
    .X(_0321_));
 sky130_fd_sc_hd__and2_1 _2440_ (.A(_0315_),
    .B(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_2 _2441_ (.A(_0315_),
    .B(_0321_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor2_1 _2442_ (.A(_0322_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_1 _2443_ (.A1(_0141_),
    .A2(_0304_),
    .B1(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__and3_1 _2444_ (.A(_0141_),
    .B(_0304_),
    .C(_0324_),
    .X(_0326_));
 sky130_fd_sc_hd__nand3_1 _2445_ (.A(_0303_),
    .B(_0161_),
    .C(_0300_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand3_1 _2446_ (.A(_0299_),
    .B(_0182_),
    .C(_0296_),
    .Y(_0328_));
 sky130_fd_sc_hd__nand2_2 _2447_ (.A(_0300_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a21bo_1 _2448_ (.A1(_0304_),
    .A2(_0327_),
    .B1_N(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__o21a_1 _2449_ (.A1(_0325_),
    .A2(_0326_),
    .B1(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__inv_2 _2450_ (.A(_0322_),
    .Y(_0332_));
 sky130_fd_sc_hd__nand2_1 _2451_ (.A(_0141_),
    .B(_0304_),
    .Y(_0333_));
 sky130_fd_sc_hd__a21o_1 _2452_ (.A1(_0332_),
    .A2(_0333_),
    .B1(_0323_),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _2453_ (.A(_0295_),
    .B(_0288_),
    .X(_0335_));
 sky130_fd_sc_hd__a21o_1 _2454_ (.A1(_0182_),
    .A2(_0335_),
    .B1(_0299_),
    .X(_0336_));
 sky130_fd_sc_hd__a21o_1 _2455_ (.A1(_0161_),
    .A2(_0336_),
    .B1(_0303_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _2456_ (.A(_0141_),
    .B(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_1 _2457_ (.A(_0322_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__and3_1 _2458_ (.A(\top8227.PSRCurrentValue[3] ),
    .B(_1246_),
    .C(_0250_),
    .X(_0340_));
 sky130_fd_sc_hd__buf_2 _2459_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_1 _2460_ (.A(_1270_),
    .B(_1298_),
    .Y(_0342_));
 sky130_fd_sc_hd__a2111oi_1 _2461_ (.A1(_1005_),
    .A2(_1411_),
    .B1(_1276_),
    .C1(_1292_),
    .D1(_1248_),
    .Y(_0343_));
 sky130_fd_sc_hd__a22o_1 _2462_ (.A1(_1184_),
    .A2(_1273_),
    .B1(_1420_),
    .B2(_1127_),
    .X(_0344_));
 sky130_fd_sc_hd__o31a_1 _2463_ (.A1(_1005_),
    .A2(_1009_),
    .A3(_0965_),
    .B1(_1096_),
    .X(_0345_));
 sky130_fd_sc_hd__or3_1 _2464_ (.A(_1279_),
    .B(_0344_),
    .C(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__a211o_1 _2465_ (.A1(_1005_),
    .A2(_0923_),
    .B1(_1282_),
    .C1(_0982_),
    .X(_0347_));
 sky130_fd_sc_hd__or3_1 _2466_ (.A(_1357_),
    .B(_0346_),
    .C(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__a2111oi_1 _2467_ (.A1(_1005_),
    .A2(_0949_),
    .B1(_1251_),
    .C1(_1256_),
    .D1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__a31o_2 _2468_ (.A1(_0342_),
    .A2(net30),
    .A3(net23),
    .B1(_1491_),
    .X(_0350_));
 sky130_fd_sc_hd__inv_2 _2469_ (.A(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__o31a_1 _2470_ (.A1(_0339_),
    .A2(_0341_),
    .A3(_0323_),
    .B1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__o21a_1 _2471_ (.A1(_0877_),
    .A2(_1151_),
    .B1(_1005_),
    .X(_0353_));
 sky130_fd_sc_hd__o21a_1 _2472_ (.A1(_1249_),
    .A2(_0353_),
    .B1(_1245_),
    .X(_0354_));
 sky130_fd_sc_hd__inv_2 _2473_ (.A(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nor2_1 _2474_ (.A(_0239_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__o32a_2 _2475_ (.A1(_1261_),
    .A2(_0331_),
    .A3(_0334_),
    .B1(_0352_),
    .B2(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__o21a_1 _2476_ (.A1(_1493_),
    .A2(_0245_),
    .B1(_0237_),
    .X(_0358_));
 sky130_fd_sc_hd__o21a_1 _2477_ (.A1(_0886_),
    .A2(_1184_),
    .B1(_1014_),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _2478_ (.A(_1246_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_2 _2479_ (.A(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__a211oi_1 _2480_ (.A1(_1246_),
    .A2(_1257_),
    .B1(_0361_),
    .C1(_0827_),
    .Y(_0362_));
 sky130_fd_sc_hd__a41o_1 _2481_ (.A1(_0916_),
    .A2(\top8227.demux.setInterruptFlag ),
    .A3(_1078_),
    .A4(_1096_),
    .B1(_0832_),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_4 _2482_ (.A(_1267_),
    .B(_1260_),
    .Y(_0364_));
 sky130_fd_sc_hd__o21a_1 _2483_ (.A1(_0898_),
    .A2(_0905_),
    .B1(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _2484_ (.A0(_0362_),
    .A1(_0363_),
    .S(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__a21o_1 _2485_ (.A1(_0358_),
    .A2(_0361_),
    .B1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__a31o_1 _2486_ (.A1(_1247_),
    .A2(_1257_),
    .A3(_0357_),
    .B1(_0367_),
    .X(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[0] ));
 sky130_fd_sc_hd__nand2_1 _2487_ (.A(_1247_),
    .B(_0359_),
    .Y(_0368_));
 sky130_fd_sc_hd__o21a_1 _2488_ (.A1(_1295_),
    .A2(_1325_),
    .B1(_1015_),
    .X(_0369_));
 sky130_fd_sc_hd__o31a_1 _2489_ (.A1(_0943_),
    .A2(_0944_),
    .A3(_0952_),
    .B1(_1005_),
    .X(_0370_));
 sky130_fd_sc_hd__o31a_1 _2490_ (.A1(_0891_),
    .A2(_0934_),
    .A3(_1327_),
    .B1(_1015_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _2491_ (.A(_1309_),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__or4_2 _2492_ (.A(_0369_),
    .B(_1351_),
    .C(_0370_),
    .D(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__o21ai_1 _2493_ (.A1(_1345_),
    .A2(_0373_),
    .B1(_1246_),
    .Y(_0374_));
 sky130_fd_sc_hd__or4_1 _2494_ (.A(_0176_),
    .B(_0196_),
    .C(_0217_),
    .D(_0358_),
    .X(_0375_));
 sky130_fd_sc_hd__or4_1 _2495_ (.A(_0316_),
    .B(_1494_),
    .C(_0153_),
    .D(_0374_),
    .X(_0376_));
 sky130_fd_sc_hd__nor2_1 _2496_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__mux2_1 _2497_ (.A0(_0377_),
    .A1(_0361_),
    .S(_0274_),
    .X(_0378_));
 sky130_fd_sc_hd__a31o_1 _2498_ (.A1(\top8227.PSRCurrentValue[1] ),
    .A2(_0368_),
    .A3(_0374_),
    .B1(_0378_),
    .X(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[1] ));
 sky130_fd_sc_hd__a32o_1 _2499_ (.A1(_0916_),
    .A2(\top8227.demux.setInterruptFlag ),
    .A3(_1096_),
    .B1(_0926_),
    .B2(_1006_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _2500_ (.A(_1247_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__and3_1 _2501_ (.A(_1247_),
    .B(_0363_),
    .C(_0379_),
    .X(_0381_));
 sky130_fd_sc_hd__a31o_1 _2502_ (.A1(\top8227.PSRCurrentValue[2] ),
    .A2(_0368_),
    .A3(_0380_),
    .B1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__a21o_1 _2503_ (.A1(_0217_),
    .A2(_0361_),
    .B1(_0382_),
    .X(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[2] ));
 sky130_fd_sc_hd__a21o_1 _2504_ (.A1(_0849_),
    .A2(_0921_),
    .B1(_0904_),
    .X(_0383_));
 sky130_fd_sc_hd__a21oi_1 _2505_ (.A1(_0364_),
    .A2(_0383_),
    .B1(_0361_),
    .Y(_0384_));
 sky130_fd_sc_hd__a32o_1 _2506_ (.A1(_0364_),
    .A2(_0363_),
    .A3(_0383_),
    .B1(_0384_),
    .B2(\top8227.PSRCurrentValue[3] ),
    .X(_0385_));
 sky130_fd_sc_hd__a21o_1 _2507_ (.A1(_0196_),
    .A2(_0361_),
    .B1(_0385_),
    .X(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[3] ));
 sky130_fd_sc_hd__nand2_1 _2508_ (.A(_1246_),
    .B(_0250_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _2509_ (.A1(_1006_),
    .A2(_0950_),
    .B1(_0359_),
    .Y(_0387_));
 sky130_fd_sc_hd__o2bb2a_1 _2510_ (.A1_N(_0924_),
    .A2_N(_0364_),
    .B1(_0387_),
    .B2(_1260_),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_2 _2511_ (.A(gpio[20]),
    .B(_1010_),
    .Y(_0389_));
 sky130_fd_sc_hd__a32o_1 _2512_ (.A1(\top8227.PSRCurrentValue[6] ),
    .A2(_0386_),
    .A3(_0388_),
    .B1(_0389_),
    .B2(\top8227.negEdgeDetector.q1 ),
    .X(_0390_));
 sky130_fd_sc_hd__and3b_1 _2513_ (.A_N(_0387_),
    .B(_1494_),
    .C(_1247_),
    .X(_0391_));
 sky130_fd_sc_hd__inv_2 _2514_ (.A(_0323_),
    .Y(_0392_));
 sky130_fd_sc_hd__a2111o_1 _2515_ (.A1(_0338_),
    .A2(_0392_),
    .B1(_0339_),
    .C1(\top8227.PSRCurrentValue[3] ),
    .D1(_0386_),
    .X(_0393_));
 sky130_fd_sc_hd__or3b_1 _2516_ (.A(_0390_),
    .B(_0391_),
    .C_N(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(_0394_),
    .X(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[6] ));
 sky130_fd_sc_hd__and2_2 _2518_ (.A(clknet_4_6_0_clk),
    .B(\top8227.pulse_slower.nextEnableState[0] ),
    .X(_0395_));
 sky130_fd_sc_hd__buf_1 _2519_ (.A(_0395_),
    .X(gpio[24]));
 sky130_fd_sc_hd__nand2_2 _2520_ (.A(gpio[18]),
    .B(_1079_),
    .Y(net18));
 sky130_fd_sc_hd__nand2_1 _2521_ (.A(_0868_),
    .B(_0364_),
    .Y(_0396_));
 sky130_fd_sc_hd__and4b_1 _2522_ (.A_N(_1021_),
    .B(_0868_),
    .C(_0364_),
    .D(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _2523_ (.A1(net56),
    .A2(_0396_),
    .B1(_0397_),
    .B2(_0357_),
    .X(_0026_));
 sky130_fd_sc_hd__a21bo_1 _2524_ (.A1(_0987_),
    .A2(_1262_),
    .B1_N(_1422_),
    .X(_0398_));
 sky130_fd_sc_hd__o211a_1 _2525_ (.A1(_0982_),
    .A2(_1298_),
    .B1(_0398_),
    .C1(_0986_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\top8227.freeCarry ),
    .A1(_0357_),
    .S(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(_0400_),
    .X(_0027_));
 sky130_fd_sc_hd__inv_2 _2528_ (.A(net55),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(_0401_),
    .B(_0986_),
    .Y(_0028_));
 sky130_fd_sc_hd__or3_1 _2530_ (.A(\top8227.PSRCurrentValue[2] ),
    .B(\top8227.demux.setInterruptFlag ),
    .C(_1010_),
    .X(_0402_));
 sky130_fd_sc_hd__or2_1 _2531_ (.A(\top8227.demux.nmi ),
    .B(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _2532_ (.A1(\top8227.demux.nmi ),
    .A2(_0381_),
    .B1(_0403_),
    .B2(net53),
    .X(_0029_));
 sky130_fd_sc_hd__o21ba_1 _2533_ (.A1(net82),
    .A2(_0986_),
    .B1_N(_0389_),
    .X(_0030_));
 sky130_fd_sc_hd__nor2_1 _2534_ (.A(_1010_),
    .B(_1018_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2b_1 _2535_ (.A_N(_0380_),
    .B(_0363_),
    .Y(_0405_));
 sky130_fd_sc_hd__o21a_1 _2536_ (.A1(net67),
    .A2(_0404_),
    .B1(_0405_),
    .X(_0031_));
 sky130_fd_sc_hd__or3b_1 _2537_ (.A(\top8227.demux.nmi ),
    .B(\top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ),
    .C_N(\top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI ),
    .X(_0406_));
 sky130_fd_sc_hd__a21bo_1 _2538_ (.A1(\top8227.demux.nmi ),
    .A2(_0405_),
    .B1_N(_0406_),
    .X(_0032_));
 sky130_fd_sc_hd__or4b_1 _2539_ (.A(\top8227.PSRCurrentValue[2] ),
    .B(\top8227.demux.setInterruptFlag ),
    .C(\top8227.instructionLoader.interruptInjector.irqGenerated ),
    .D_N(\top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ ),
    .X(_0407_));
 sky130_fd_sc_hd__a21bo_1 _2540_ (.A1(net62),
    .A2(_0405_),
    .B1_N(_0407_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _2541_ (.A(_1315_),
    .B(_1464_),
    .Y(_0408_));
 sky130_fd_sc_hd__a211o_1 _2542_ (.A1(_1127_),
    .A2(_1274_),
    .B1(_1288_),
    .C1(_0982_),
    .X(_0409_));
 sky130_fd_sc_hd__a221o_1 _2543_ (.A1(_1006_),
    .A2(_1294_),
    .B1(_0882_),
    .B2(_1015_),
    .C1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__and3_1 _2544_ (.A(_0985_),
    .B(_0408_),
    .C(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__buf_4 _2545_ (.A(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(net10),
    .A1(_0358_),
    .S(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(_0413_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(net85),
    .A1(_0274_),
    .S(_0412_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_0414_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(net79),
    .A1(_0217_),
    .S(_0412_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _2551_ (.A(_0415_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(net13),
    .A1(_0196_),
    .S(_0412_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _2553_ (.A(_0416_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(net14),
    .A1(_0176_),
    .S(_0412_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _2555_ (.A(_0417_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2556_ (.A0(net86),
    .A1(_0153_),
    .S(_0412_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _2557_ (.A(_0418_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(net16),
    .A1(_1494_),
    .S(_0412_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _2559_ (.A(_0419_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(net84),
    .A1(_0316_),
    .S(_0412_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _2561_ (.A(_0420_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_1 _2562_ (.A(_0955_),
    .B(_0901_),
    .C(_0854_),
    .X(_0421_));
 sky130_fd_sc_hd__o221ai_1 _2563_ (.A1(_1016_),
    .A2(\top8227.demux.state_machine.currentAddress[6] ),
    .B1(_1428_),
    .B2(_0421_),
    .C1(_1267_),
    .Y(_0422_));
 sky130_fd_sc_hd__nor3_1 _2564_ (.A(_0909_),
    .B(_1270_),
    .C(_1427_),
    .Y(_0423_));
 sky130_fd_sc_hd__a221o_1 _2565_ (.A1(_0982_),
    .A2(_0422_),
    .B1(_0423_),
    .B2(_1336_),
    .C1(_0976_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_4 _2566_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__a2bb2oi_4 _2567_ (.A1_N(\top8227.demux.nmi ),
    .A2_N(\top8227.instructionLoader.interruptInjector.irqGenerated ),
    .B1(net29),
    .B2(_0401_),
    .Y(_0426_));
 sky130_fd_sc_hd__a31o_1 _2568_ (.A1(_0903_),
    .A2(_1346_),
    .A3(_0364_),
    .B1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _2569_ (.A(_0837_),
    .B(_0844_),
    .C(_0858_),
    .X(_0428_));
 sky130_fd_sc_hd__and2_1 _2570_ (.A(_0868_),
    .B(_1273_),
    .X(_0429_));
 sky130_fd_sc_hd__o41a_1 _2571_ (.A1(_1013_),
    .A2(_0816_),
    .A3(_0428_),
    .A4(_1274_),
    .B1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__or3_1 _2572_ (.A(_0859_),
    .B(\top8227.demux.state_machine.timeState[1] ),
    .C(\top8227.demux.state_machine.timeState[5] ),
    .X(_0431_));
 sky130_fd_sc_hd__or2_1 _2573_ (.A(\top8227.demux.state_machine.timeState[5] ),
    .B(\top8227.demux.state_machine.timeState[3] ),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _2574_ (.A1(_0818_),
    .A2(_0898_),
    .B1(_0951_),
    .B2(_1316_),
    .X(_0433_));
 sky130_fd_sc_hd__a221o_1 _2575_ (.A1(_0914_),
    .A2(_0431_),
    .B1(_0432_),
    .B2(_0896_),
    .C1(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o22a_1 _2576_ (.A1(\top8227.demux.state_machine.timeState[1] ),
    .A2(_0916_),
    .B1(_0912_),
    .B2(_0915_),
    .X(_0435_));
 sky130_fd_sc_hd__nand2_1 _2577_ (.A(_0971_),
    .B(_1419_),
    .Y(_0436_));
 sky130_fd_sc_hd__or4_1 _2578_ (.A(_1413_),
    .B(_0434_),
    .C(_0435_),
    .D(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__or4_1 _2579_ (.A(_1399_),
    .B(_1409_),
    .C(_0430_),
    .D(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__o21ai_1 _2580_ (.A1(_1002_),
    .A2(_0421_),
    .B1(_1016_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _2581_ (.A(\top8227.demux.state_machine.currentAddress[6] ),
    .B(_1273_),
    .Y(_0440_));
 sky130_fd_sc_hd__nand3_1 _2582_ (.A(_1422_),
    .B(_0439_),
    .C(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand3_1 _2583_ (.A(_0985_),
    .B(_0438_),
    .C(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__nor2b_2 _2584_ (.A(_0427_),
    .B_N(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__and2_2 _2585_ (.A(_0425_),
    .B(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_4 _2586_ (.A(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__or2_1 _2587_ (.A(_0231_),
    .B(_0232_),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_2 _2588_ (.A1(_1245_),
    .A2(_1334_),
    .B1(_1340_),
    .X(_0447_));
 sky130_fd_sc_hd__nor2b_2 _2589_ (.A(_0447_),
    .B_N(_1312_),
    .Y(_0448_));
 sky130_fd_sc_hd__and2b_1 _2590_ (.A_N(_0235_),
    .B(_0236_),
    .X(_0449_));
 sky130_fd_sc_hd__or3b_1 _2591_ (.A(_1312_),
    .B(_0447_),
    .C_N(_1493_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_2 _2592_ (.A(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_1 _2593_ (.A(_0449_),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__a221o_2 _2594_ (.A1(_0446_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0245_),
    .C1(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__or2_1 _2595_ (.A(_0442_),
    .B(_0426_),
    .X(_0454_));
 sky130_fd_sc_hd__buf_2 _2596_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__buf_2 _2597_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__buf_2 _2598_ (.A(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_4 _2599_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_4 _2600_ (.A(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__or2_1 _2601_ (.A(_0279_),
    .B(_0243_),
    .X(_0460_));
 sky130_fd_sc_hd__or2_1 _2602_ (.A(_0222_),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__nor3_1 _2603_ (.A(_0179_),
    .B(_0201_),
    .C(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__or2b_1 _2604_ (.A(_0159_),
    .B_N(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__or2_1 _2605_ (.A(_0134_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_1 _2606_ (.A(_0320_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _2607_ (.A(_0222_),
    .Y(_0466_));
 sky130_fd_sc_hd__nand2_1 _2608_ (.A(_0279_),
    .B(_0243_),
    .Y(_0467_));
 sky130_fd_sc_hd__nor2_1 _2609_ (.A(_0466_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__and2_1 _2610_ (.A(_0201_),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__and3_1 _2611_ (.A(_0180_),
    .B(_0427_),
    .C(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__and3_1 _2612_ (.A(_0135_),
    .B(_0159_),
    .C(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__inv_2 _2613_ (.A(_0455_),
    .Y(_0472_));
 sky130_fd_sc_hd__a21o_1 _2614_ (.A1(_0320_),
    .A2(_0471_),
    .B1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__o21ai_1 _2615_ (.A1(_0459_),
    .A2(_0465_),
    .B1(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__xnor2_1 _2616_ (.A(_0453_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__inv_2 _2617_ (.A(_0424_),
    .Y(_0476_));
 sky130_fd_sc_hd__clkbuf_4 _2618_ (.A(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__and2_1 _2619_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[16] ),
    .B(_0456_),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_1 _2620_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[16] ),
    .B(_0456_),
    .Y(_0479_));
 sky130_fd_sc_hd__nor2_1 _2621_ (.A(_0478_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__or2_1 _2622_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ),
    .B(_0456_),
    .X(_0481_));
 sky130_fd_sc_hd__and2_1 _2623_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[22] ),
    .B(_0456_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_1 _2624_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[22] ),
    .B(_0456_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_1 _2625_ (.A(_0482_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _2626_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[20] ),
    .Y(_0485_));
 sky130_fd_sc_hd__nor2_1 _2627_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[21] ),
    .B(_0456_),
    .Y(_0486_));
 sky130_fd_sc_hd__xnor2_1 _2628_ (.A(_0485_),
    .B(_0455_),
    .Y(_0487_));
 sky130_fd_sc_hd__or2_1 _2629_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[19] ),
    .B(_0455_),
    .X(_0488_));
 sky130_fd_sc_hd__xor2_1 _2630_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[18] ),
    .B(_0455_),
    .X(_0489_));
 sky130_fd_sc_hd__or3_1 _2631_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[17] ),
    .B(_0442_),
    .C(_0426_),
    .X(_0490_));
 sky130_fd_sc_hd__o21a_1 _2632_ (.A1(_0442_),
    .A2(_0426_),
    .B1(\top8227.internalDataflow.addressLowBusModule.busInputs[17] ),
    .X(_0491_));
 sky130_fd_sc_hd__a21o_1 _2633_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[16] ),
    .A2(_0490_),
    .B1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__and2_1 _2634_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[18] ),
    .B(_0455_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _2635_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[19] ),
    .B(_0455_),
    .X(_0494_));
 sky130_fd_sc_hd__a311o_1 _2636_ (.A1(_0488_),
    .A2(_0489_),
    .A3(_0492_),
    .B1(_0493_),
    .C1(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nand2_1 _2637_ (.A(_0487_),
    .B(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _2638_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[21] ),
    .B(_0456_),
    .Y(_0497_));
 sky130_fd_sc_hd__o221ai_4 _2639_ (.A1(_0485_),
    .A2(_0472_),
    .B1(_0486_),
    .B2(_0496_),
    .C1(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__and2_1 _2640_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ),
    .B(_0456_),
    .X(_0499_));
 sky130_fd_sc_hd__a311o_1 _2641_ (.A1(_0481_),
    .A2(_0484_),
    .A3(_0498_),
    .B1(_0482_),
    .C1(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__or2_1 _2642_ (.A(_0480_),
    .B(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__nand2_1 _2643_ (.A(_0480_),
    .B(_0500_),
    .Y(_0502_));
 sky130_fd_sc_hd__nor2_4 _2644_ (.A(_0476_),
    .B(_0443_),
    .Y(_0503_));
 sky130_fd_sc_hd__and3_1 _2645_ (.A(_0501_),
    .B(_0502_),
    .C(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__a221o_1 _2646_ (.A1(net75),
    .A2(_0445_),
    .B1(_0475_),
    .B2(_0477_),
    .C1(_0504_),
    .X(_0042_));
 sky130_fd_sc_hd__nor2_1 _2647_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[17] ),
    .B(_0459_),
    .Y(_0505_));
 sky130_fd_sc_hd__and2_1 _2648_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[17] ),
    .B(_0457_),
    .X(_0506_));
 sky130_fd_sc_hd__nor2_1 _2649_ (.A(_0505_),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__a21oi_1 _2650_ (.A1(_0480_),
    .A2(_0500_),
    .B1(_0478_),
    .Y(_0508_));
 sky130_fd_sc_hd__xnor2_1 _2651_ (.A(_0507_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nor2_1 _2652_ (.A(_0263_),
    .B(_0451_),
    .Y(_0510_));
 sky130_fd_sc_hd__a221o_2 _2653_ (.A1(_0269_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0268_),
    .C1(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__and2_1 _2654_ (.A(_0453_),
    .B(_0465_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_1 _2655_ (.A(_0459_),
    .B(_0453_),
    .Y(_0513_));
 sky130_fd_sc_hd__o211a_1 _2656_ (.A1(_0459_),
    .A2(_0512_),
    .B1(_0513_),
    .C1(_0473_),
    .X(_0514_));
 sky130_fd_sc_hd__xnor2_1 _2657_ (.A(_0511_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__nor2_1 _2658_ (.A(_0425_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__a221o_1 _2659_ (.A1(net90),
    .A2(_0445_),
    .B1(_0509_),
    .B2(_0503_),
    .C1(_0516_),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_1 _2660_ (.A(_0207_),
    .B(_0451_),
    .Y(_0517_));
 sky130_fd_sc_hd__a221o_2 _2661_ (.A1(_0213_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0212_),
    .C1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__a31o_1 _2662_ (.A1(_0453_),
    .A2(_0465_),
    .A3(_0511_),
    .B1(_0458_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _2663_ (.A(_0453_),
    .B(_0511_),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_1 _2664_ (.A(_0459_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__and3_1 _2665_ (.A(_0473_),
    .B(_0519_),
    .C(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__xor2_1 _2666_ (.A(_0518_),
    .B(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__xor2_1 _2667_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[18] ),
    .B(_0457_),
    .X(_0524_));
 sky130_fd_sc_hd__or2_1 _2668_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[17] ),
    .B(_0456_),
    .X(_0525_));
 sky130_fd_sc_hd__a311o_1 _2669_ (.A1(_0480_),
    .A2(_0500_),
    .A3(_0525_),
    .B1(_0506_),
    .C1(_0478_),
    .X(_0526_));
 sky130_fd_sc_hd__and2_1 _2670_ (.A(_0524_),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__or2_1 _2671_ (.A(_0524_),
    .B(_0526_),
    .X(_0528_));
 sky130_fd_sc_hd__and3b_1 _2672_ (.A_N(_0527_),
    .B(_0503_),
    .C(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__a221o_1 _2673_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[18] ),
    .A2(_0445_),
    .B1(_0523_),
    .B2(_0477_),
    .C1(_0529_),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_1 _2674_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[19] ),
    .B(_0458_),
    .Y(_0530_));
 sky130_fd_sc_hd__and2_1 _2675_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[19] ),
    .B(_0457_),
    .X(_0531_));
 sky130_fd_sc_hd__a21o_1 _2676_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[18] ),
    .A2(_0457_),
    .B1(_0527_),
    .X(_0532_));
 sky130_fd_sc_hd__o21bai_1 _2677_ (.A1(_0530_),
    .A2(_0531_),
    .B1_N(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__or3b_1 _2678_ (.A(_0530_),
    .B(_0531_),
    .C_N(_0532_),
    .X(_0534_));
 sky130_fd_sc_hd__nor2_1 _2679_ (.A(_0185_),
    .B(_0451_),
    .Y(_0535_));
 sky130_fd_sc_hd__a221o_2 _2680_ (.A1(_0191_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0190_),
    .C1(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _2681_ (.A(_0201_),
    .B(_0468_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _2682_ (.A(_0135_),
    .B(_0159_),
    .Y(_0538_));
 sky130_fd_sc_hd__or2_1 _2683_ (.A(_0472_),
    .B(_0443_),
    .X(_0539_));
 sky130_fd_sc_hd__or4bb_1 _2684_ (.A(_0538_),
    .B(_0539_),
    .C_N(_0320_),
    .D_N(_0180_),
    .X(_0540_));
 sky130_fd_sc_hd__or4_1 _2685_ (.A(_0537_),
    .B(_0518_),
    .C(_0520_),
    .D(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__nand4_1 _2686_ (.A(_0472_),
    .B(_0511_),
    .C(_0512_),
    .D(_0518_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _2687_ (.A(_0541_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__xnor2_1 _2688_ (.A(_0536_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_1 _2689_ (.A(_0425_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a31o_1 _2690_ (.A1(_0425_),
    .A2(_0533_),
    .A3(_0534_),
    .B1(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _2691_ (.A0(_0546_),
    .A1(\top8227.internalDataflow.addressHighBusModule.busInputs[19] ),
    .S(_0444_),
    .X(_0547_));
 sky130_fd_sc_hd__clkbuf_1 _2692_ (.A(_0547_),
    .X(_0045_));
 sky130_fd_sc_hd__xor2_1 _2693_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[20] ),
    .B(_0457_),
    .X(_0548_));
 sky130_fd_sc_hd__o21a_1 _2694_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[19] ),
    .A2(_0457_),
    .B1(_0532_),
    .X(_0549_));
 sky130_fd_sc_hd__or3_1 _2695_ (.A(_0531_),
    .B(_0548_),
    .C(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__o21ai_1 _2696_ (.A1(_0531_),
    .A2(_0549_),
    .B1(_0548_),
    .Y(_0551_));
 sky130_fd_sc_hd__and2b_1 _2697_ (.A_N(_0451_),
    .B(_0173_),
    .X(_0552_));
 sky130_fd_sc_hd__a221o_2 _2698_ (.A1(_0167_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0166_),
    .C1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(_0541_),
    .A1(_0542_),
    .S(_0536_),
    .X(_0554_));
 sky130_fd_sc_hd__xnor2_1 _2700_ (.A(_0553_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__a22o_1 _2701_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[20] ),
    .A2(_0445_),
    .B1(_0555_),
    .B2(_0477_),
    .X(_0556_));
 sky130_fd_sc_hd__a31o_1 _2702_ (.A1(_0503_),
    .A2(_0550_),
    .A3(_0551_),
    .B1(_0556_),
    .X(_0046_));
 sky130_fd_sc_hd__or2_1 _2703_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[21] ),
    .B(_0457_),
    .X(_0557_));
 sky130_fd_sc_hd__nand2_1 _2704_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[21] ),
    .B(_0457_),
    .Y(_0558_));
 sky130_fd_sc_hd__o21a_1 _2705_ (.A1(_0531_),
    .A2(_0549_),
    .B1(_0548_),
    .X(_0559_));
 sky130_fd_sc_hd__a21o_1 _2706_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[20] ),
    .A2(_0457_),
    .B1(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _2707_ (.A1(_0557_),
    .A2(_0558_),
    .B1(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a31o_1 _2708_ (.A1(_0557_),
    .A2(_0558_),
    .A3(_0560_),
    .B1(_0476_),
    .X(_0562_));
 sky130_fd_sc_hd__xnor2_1 _2709_ (.A(_0458_),
    .B(_0553_),
    .Y(_0563_));
 sky130_fd_sc_hd__nor2_1 _2710_ (.A(_0554_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__and2b_1 _2711_ (.A_N(_0451_),
    .B(_0150_),
    .X(_0565_));
 sky130_fd_sc_hd__a221o_1 _2712_ (.A1(_0146_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0145_),
    .C1(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__or2_1 _2713_ (.A(_0564_),
    .B(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__a21oi_1 _2714_ (.A1(_0564_),
    .A2(_0566_),
    .B1(_0425_),
    .Y(_0568_));
 sky130_fd_sc_hd__a2bb2o_1 _2715_ (.A1_N(_0561_),
    .A2_N(_0562_),
    .B1(_0567_),
    .B2(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(_0569_),
    .A1(\top8227.internalDataflow.addressHighBusModule.busInputs[21] ),
    .S(_0444_),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_1 _2717_ (.A(_0570_),
    .X(_0047_));
 sky130_fd_sc_hd__xnor2_1 _2718_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[22] ),
    .B(_0458_),
    .Y(_0571_));
 sky130_fd_sc_hd__a21bo_1 _2719_ (.A1(_0557_),
    .A2(_0560_),
    .B1_N(_0558_),
    .X(_0572_));
 sky130_fd_sc_hd__xnor2_1 _2720_ (.A(_0571_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__and2_1 _2721_ (.A(_0458_),
    .B(_0566_),
    .X(_0574_));
 sky130_fd_sc_hd__nor2_1 _2722_ (.A(_0458_),
    .B(_0566_),
    .Y(_0575_));
 sky130_fd_sc_hd__or4_1 _2723_ (.A(_0554_),
    .B(_0563_),
    .C(_0574_),
    .D(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__and2b_1 _2724_ (.A_N(_0451_),
    .B(_1481_),
    .X(_0577_));
 sky130_fd_sc_hd__a221o_2 _2725_ (.A1(_1441_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_1396_),
    .C1(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__xor2_1 _2726_ (.A(_0576_),
    .B(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__nor2_1 _2727_ (.A(_0425_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__a221o_1 _2728_ (.A1(net76),
    .A2(_0445_),
    .B1(_0573_),
    .B2(_0503_),
    .C1(_0580_),
    .X(_0048_));
 sky130_fd_sc_hd__or2b_1 _2729_ (.A(_0571_),
    .B_N(_0572_),
    .X(_0581_));
 sky130_fd_sc_hd__a21bo_1 _2730_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[22] ),
    .A2(_0459_),
    .B1_N(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__xor2_1 _2731_ (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[23] ),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__xnor2_1 _2732_ (.A(_0472_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__xnor2_1 _2733_ (.A(_0459_),
    .B(_0578_),
    .Y(_0585_));
 sky130_fd_sc_hd__and2b_1 _2734_ (.A_N(_0451_),
    .B(_0313_),
    .X(_0586_));
 sky130_fd_sc_hd__a221o_1 _2735_ (.A1(_0309_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0308_),
    .C1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__o21ai_1 _2736_ (.A1(_0576_),
    .A2(_0585_),
    .B1(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__or3_1 _2737_ (.A(_0576_),
    .B(_0587_),
    .C(_0585_),
    .X(_0589_));
 sky130_fd_sc_hd__a21oi_1 _2738_ (.A1(_0588_),
    .A2(_0589_),
    .B1(_0425_),
    .Y(_0590_));
 sky130_fd_sc_hd__a221o_1 _2739_ (.A1(\top8227.internalDataflow.addressHighBusModule.busInputs[23] ),
    .A2(_0445_),
    .B1(_0584_),
    .B2(_0503_),
    .C1(_0590_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _2740_ (.A1(_1014_),
    .A2(_0890_),
    .B1(_1214_),
    .B2(_1006_),
    .X(_0591_));
 sky130_fd_sc_hd__or4b_2 _2741_ (.A(_1348_),
    .B(_1496_),
    .C(_0591_),
    .D_N(_1352_),
    .X(_0592_));
 sky130_fd_sc_hd__nand2_4 _2742_ (.A(_1247_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__mux2_1 _2743_ (.A0(_0238_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[32] ),
    .S(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_1 _2744_ (.A(_0594_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(_0271_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[33] ),
    .S(_0593_),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_1 _2746_ (.A(_0595_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(_0215_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[34] ),
    .S(_0593_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_1 _2748_ (.A(_0596_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2749_ (.A0(_0193_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[35] ),
    .S(_0593_),
    .X(_0597_));
 sky130_fd_sc_hd__clkbuf_1 _2750_ (.A(_0597_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(_0174_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[36] ),
    .S(_0593_),
    .X(_0598_));
 sky130_fd_sc_hd__clkbuf_1 _2752_ (.A(_0598_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(_0151_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[37] ),
    .S(_0593_),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_1 _2754_ (.A(_0599_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(_1482_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[38] ),
    .S(_0593_),
    .X(_0600_));
 sky130_fd_sc_hd__clkbuf_1 _2756_ (.A(_0600_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(_0314_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[39] ),
    .S(_0593_),
    .X(_0601_));
 sky130_fd_sc_hd__clkbuf_1 _2758_ (.A(_0601_),
    .X(_0057_));
 sky130_fd_sc_hd__or3_1 _2759_ (.A(_0932_),
    .B(_0944_),
    .C(_1197_),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _2760_ (.A1(_1015_),
    .A2(_0948_),
    .B1(_0602_),
    .B2(_1006_),
    .X(_0603_));
 sky130_fd_sc_hd__and2_1 _2761_ (.A(_1246_),
    .B(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_4 _2762_ (.A(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(\top8227.internalDataflow.stackBusModule.busInputs[40] ),
    .A1(_0238_),
    .S(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_0606_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2765_ (.A0(\top8227.internalDataflow.stackBusModule.busInputs[41] ),
    .A1(_0271_),
    .S(_0605_),
    .X(_0607_));
 sky130_fd_sc_hd__clkbuf_1 _2766_ (.A(_0607_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2767_ (.A0(net68),
    .A1(_0215_),
    .S(_0605_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_1 _2768_ (.A(_0608_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(net72),
    .A1(_0193_),
    .S(_0605_),
    .X(_0609_));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(_0609_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2771_ (.A0(net65),
    .A1(_0174_),
    .S(_0605_),
    .X(_0610_));
 sky130_fd_sc_hd__clkbuf_1 _2772_ (.A(_0610_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(net71),
    .A1(_0151_),
    .S(_0605_),
    .X(_0611_));
 sky130_fd_sc_hd__clkbuf_1 _2774_ (.A(_0611_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(net66),
    .A1(_1482_),
    .S(_0605_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_1 _2776_ (.A(_0612_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(net81),
    .A1(_0314_),
    .S(_0605_),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_1 _2778_ (.A(_0613_),
    .X(_0065_));
 sky130_fd_sc_hd__a22o_1 _2779_ (.A1(\top8227.instructionLoader.interruptInjector.resetDetected ),
    .A2(_0986_),
    .B1(_0402_),
    .B2(\top8227.demux.reset ),
    .X(_0066_));
 sky130_fd_sc_hd__a221o_1 _2780_ (.A1(_1006_),
    .A2(\top8227.demux.state_machine.currentAddress[5] ),
    .B1(_1301_),
    .B2(_1262_),
    .C1(_1499_),
    .X(_0614_));
 sky130_fd_sc_hd__a21o_1 _2781_ (.A1(_1016_),
    .A2(_1317_),
    .B1(_1266_),
    .X(_0615_));
 sky130_fd_sc_hd__a221o_1 _2782_ (.A1(_1263_),
    .A2(_1265_),
    .B1(_1273_),
    .B2(_0615_),
    .C1(_1078_),
    .X(_0616_));
 sky130_fd_sc_hd__inv_2 _2783_ (.A(_1508_),
    .Y(_0617_));
 sky130_fd_sc_hd__and2b_1 _2784_ (.A_N(_0835_),
    .B(_0894_),
    .X(_0618_));
 sky130_fd_sc_hd__o32a_1 _2785_ (.A1(_1005_),
    .A2(_1009_),
    .A3(_0916_),
    .B1(_1184_),
    .B2(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _2786_ (.A(_1015_),
    .B(_0431_),
    .X(_0620_));
 sky130_fd_sc_hd__a221o_1 _2787_ (.A1(\top8227.demux.state_machine.timeState[3] ),
    .A2(_1096_),
    .B1(_1127_),
    .B2(_0620_),
    .C1(_0982_),
    .X(_0621_));
 sky130_fd_sc_hd__a211o_1 _2788_ (.A1(_1013_),
    .A2(_0618_),
    .B1(_0619_),
    .C1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__o21a_1 _2789_ (.A1(_1212_),
    .A2(_0887_),
    .B1(_1400_),
    .X(_0623_));
 sky130_fd_sc_hd__a2111o_1 _2790_ (.A1(_1294_),
    .A2(_1275_),
    .B1(_1347_),
    .C1(_0433_),
    .D1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or3_1 _2791_ (.A(_1406_),
    .B(_1399_),
    .C(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__or3_1 _2792_ (.A(_0910_),
    .B(_1410_),
    .C(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__or4_1 _2793_ (.A(_1407_),
    .B(_0617_),
    .C(_0622_),
    .D(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__o211a_4 _2794_ (.A1(_0614_),
    .A2(_0616_),
    .B1(_0986_),
    .C1(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _2795_ (.A0(gpio[8]),
    .A1(_0453_),
    .S(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_1 _2796_ (.A(_0629_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(gpio[9]),
    .A1(_0511_),
    .S(_0628_),
    .X(_0630_));
 sky130_fd_sc_hd__clkbuf_1 _2798_ (.A(_0630_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2799_ (.A0(gpio[10]),
    .A1(_0518_),
    .S(_0628_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _2800_ (.A(_0631_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2801_ (.A0(gpio[11]),
    .A1(_0536_),
    .S(_0628_),
    .X(_0632_));
 sky130_fd_sc_hd__clkbuf_1 _2802_ (.A(_0632_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(gpio[12]),
    .A1(_0553_),
    .S(_0628_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _2804_ (.A(_0633_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(gpio[13]),
    .A1(_0566_),
    .S(_0628_),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_1 _2806_ (.A(_0634_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2807_ (.A0(gpio[14]),
    .A1(_0578_),
    .S(_0628_),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_1 _2808_ (.A(_0635_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(gpio[15]),
    .A1(_0587_),
    .S(_0628_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_1 _2810_ (.A(_0636_),
    .X(_0074_));
 sky130_fd_sc_hd__inv_2 _2811_ (.A(_0243_),
    .Y(_0637_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(\top8227.internalDataflow.addressLowBusModule.busInputs[16] ),
    .A1(_0637_),
    .S(_0477_),
    .X(_0638_));
 sky130_fd_sc_hd__xnor2_1 _2813_ (.A(_0443_),
    .B(_0638_),
    .Y(_0075_));
 sky130_fd_sc_hd__o21ai_1 _2814_ (.A1(_0243_),
    .A2(_0472_),
    .B1(_0539_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _2815_ (.A(_0467_),
    .B(_0460_),
    .Y(_0640_));
 sky130_fd_sc_hd__xnor2_1 _2816_ (.A(_0639_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__and2b_1 _2817_ (.A_N(_0491_),
    .B(_0490_),
    .X(_0642_));
 sky130_fd_sc_hd__nand2_1 _2818_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[16] ),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__or2_1 _2819_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[16] ),
    .B(_0642_),
    .X(_0644_));
 sky130_fd_sc_hd__a32o_1 _2820_ (.A1(_0643_),
    .A2(_0503_),
    .A3(_0644_),
    .B1(_0445_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[17] ),
    .X(_0645_));
 sky130_fd_sc_hd__a21o_1 _2821_ (.A1(_0477_),
    .A2(_0641_),
    .B1(_0645_),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _2822_ (.A(_0489_),
    .B(_0492_),
    .X(_0646_));
 sky130_fd_sc_hd__nor2_1 _2823_ (.A(_0489_),
    .B(_0492_),
    .Y(_0647_));
 sky130_fd_sc_hd__or4_1 _2824_ (.A(_0646_),
    .B(_0477_),
    .C(_0443_),
    .D(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__a22o_1 _2825_ (.A1(_0459_),
    .A2(_0467_),
    .B1(_0460_),
    .B2(_0539_),
    .X(_0649_));
 sky130_fd_sc_hd__xnor2_1 _2826_ (.A(_0222_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__o2bb2a_1 _2827_ (.A1_N(\top8227.internalDataflow.addressLowBusModule.busInputs[18] ),
    .A2_N(_0445_),
    .B1(_0650_),
    .B2(_0425_),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _2828_ (.A(_0648_),
    .B(_0651_),
    .Y(_0077_));
 sky130_fd_sc_hd__and2b_1 _2829_ (.A_N(_0494_),
    .B(_0488_),
    .X(_0652_));
 sky130_fd_sc_hd__o21ai_1 _2830_ (.A1(_0493_),
    .A2(_0646_),
    .B1(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__o31a_1 _2831_ (.A1(_0493_),
    .A2(_0646_),
    .A3(_0652_),
    .B1(_0425_),
    .X(_0654_));
 sky130_fd_sc_hd__o32a_1 _2832_ (.A1(_0466_),
    .A2(_0467_),
    .A3(_0539_),
    .B1(_0461_),
    .B2(_0458_),
    .X(_0655_));
 sky130_fd_sc_hd__xor2_1 _2833_ (.A(_0201_),
    .B(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__a22o_1 _2834_ (.A1(_0653_),
    .A2(_0654_),
    .B1(_0656_),
    .B2(_0477_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(_0657_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[19] ),
    .S(_0444_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_1 _2836_ (.A(_0658_),
    .X(_0078_));
 sky130_fd_sc_hd__o21a_1 _2837_ (.A1(_0201_),
    .A2(_0461_),
    .B1(_0180_),
    .X(_0659_));
 sky130_fd_sc_hd__or2_1 _2838_ (.A(_0458_),
    .B(_0462_),
    .X(_0660_));
 sky130_fd_sc_hd__a21oi_1 _2839_ (.A1(_0427_),
    .A2(_0469_),
    .B1(_0180_),
    .Y(_0661_));
 sky130_fd_sc_hd__o21a_1 _2840_ (.A1(_0470_),
    .A2(_0661_),
    .B1(_0459_),
    .X(_0662_));
 sky130_fd_sc_hd__o21bai_1 _2841_ (.A1(_0659_),
    .A2(_0660_),
    .B1_N(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__and2_1 _2842_ (.A(_0496_),
    .B(_0503_),
    .X(_0664_));
 sky130_fd_sc_hd__o21a_1 _2843_ (.A1(_0487_),
    .A2(_0495_),
    .B1(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__a221o_1 _2844_ (.A1(net88),
    .A2(_0445_),
    .B1(_0663_),
    .B2(_0477_),
    .C1(_0665_),
    .X(_0079_));
 sky130_fd_sc_hd__o21a_1 _2845_ (.A1(_0472_),
    .A2(_0470_),
    .B1(_0660_),
    .X(_0666_));
 sky130_fd_sc_hd__xnor2_1 _2846_ (.A(_0159_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__o21ai_1 _2847_ (.A1(_0485_),
    .A2(_0472_),
    .B1(_0496_),
    .Y(_0668_));
 sky130_fd_sc_hd__or2_1 _2848_ (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[21] ),
    .B(_0458_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2_1 _2849_ (.A(_0497_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__xnor2_1 _2850_ (.A(_0668_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(_0667_),
    .A1(_0671_),
    .S(_0425_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(_0672_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[21] ),
    .S(_0444_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _2853_ (.A(_0673_),
    .X(_0080_));
 sky130_fd_sc_hd__nand2_1 _2854_ (.A(_0472_),
    .B(_0464_),
    .Y(_0674_));
 sky130_fd_sc_hd__a21o_1 _2855_ (.A1(_0135_),
    .A2(_0463_),
    .B1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__a21oi_1 _2856_ (.A1(_0157_),
    .A2(_0470_),
    .B1(_0135_),
    .Y(_0676_));
 sky130_fd_sc_hd__o21ai_1 _2857_ (.A1(_0471_),
    .A2(_0676_),
    .B1(_0459_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _2858_ (.A(_0675_),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__and2_1 _2859_ (.A(_0484_),
    .B(_0498_),
    .X(_0679_));
 sky130_fd_sc_hd__or2_1 _2860_ (.A(_0484_),
    .B(_0498_),
    .X(_0680_));
 sky130_fd_sc_hd__and3b_1 _2861_ (.A_N(_0679_),
    .B(_0503_),
    .C(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__a221o_1 _2862_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[22] ),
    .A2(_0445_),
    .B1(_0678_),
    .B2(_0477_),
    .C1(_0681_),
    .X(_0081_));
 sky130_fd_sc_hd__nor2_1 _2863_ (.A(_0482_),
    .B(_0679_),
    .Y(_0682_));
 sky130_fd_sc_hd__and2b_1 _2864_ (.A_N(_0499_),
    .B(_0481_),
    .X(_0683_));
 sky130_fd_sc_hd__xnor2_1 _2865_ (.A(_0682_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__o21a_1 _2866_ (.A1(_0472_),
    .A2(_0471_),
    .B1(_0674_),
    .X(_0685_));
 sky130_fd_sc_hd__xnor2_1 _2867_ (.A(_0320_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(_0684_),
    .A1(_0686_),
    .S(_0477_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _2869_ (.A0(_0687_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ),
    .S(_0444_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_1 _2870_ (.A(_0688_),
    .X(_0082_));
 sky130_fd_sc_hd__o31a_1 _2871_ (.A1(_1209_),
    .A2(_0942_),
    .A3(_0951_),
    .B1(_1015_),
    .X(_0689_));
 sky130_fd_sc_hd__o21a_1 _2872_ (.A1(_0931_),
    .A2(_0952_),
    .B1(_1006_),
    .X(_0690_));
 sky130_fd_sc_hd__o31ai_4 _2873_ (.A1(_0372_),
    .A2(_0689_),
    .A3(_0690_),
    .B1(_1247_),
    .Y(_0691_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(_0238_),
    .A1(\top8227.internalDataflow.accRegToDB[0] ),
    .S(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_0692_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(_0271_),
    .A1(\top8227.internalDataflow.accRegToDB[1] ),
    .S(_0691_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_0693_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(_0215_),
    .A1(\top8227.internalDataflow.accRegToDB[2] ),
    .S(net22),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _2879_ (.A(_0694_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2880_ (.A0(_0193_),
    .A1(\top8227.internalDataflow.accRegToDB[3] ),
    .S(_0691_),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_1 _2881_ (.A(_0695_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(_0174_),
    .A1(\top8227.internalDataflow.accRegToDB[4] ),
    .S(net22),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_1 _2883_ (.A(_0696_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(_0151_),
    .A1(\top8227.internalDataflow.accRegToDB[5] ),
    .S(net22),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_1 _2885_ (.A(_0697_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(_1482_),
    .A1(\top8227.internalDataflow.accRegToDB[6] ),
    .S(net22),
    .X(_0698_));
 sky130_fd_sc_hd__clkbuf_1 _2887_ (.A(_0698_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2888_ (.A0(_0314_),
    .A1(\top8227.internalDataflow.accRegToDB[7] ),
    .S(net22),
    .X(_0699_));
 sky130_fd_sc_hd__clkbuf_1 _2889_ (.A(_0699_),
    .X(_0090_));
 sky130_fd_sc_hd__o21a_1 _2890_ (.A1(_1014_),
    .A2(_0620_),
    .B1(_1321_),
    .X(_0700_));
 sky130_fd_sc_hd__o31a_1 _2891_ (.A1(_1009_),
    .A2(_1273_),
    .A3(_0432_),
    .B1(_1096_),
    .X(_0701_));
 sky130_fd_sc_hd__o41a_1 _2892_ (.A1(_1005_),
    .A2(_1009_),
    .A3(_0916_),
    .A4(_1400_),
    .B1(_1127_),
    .X(_0702_));
 sky130_fd_sc_hd__or4_1 _2893_ (.A(_0436_),
    .B(_0700_),
    .C(_0701_),
    .D(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__inv_2 _2894_ (.A(_1447_),
    .Y(_0704_));
 sky130_fd_sc_hd__a22o_1 _2895_ (.A1(_1016_),
    .A2(_1317_),
    .B1(_1275_),
    .B2(_0987_),
    .X(_0705_));
 sky130_fd_sc_hd__or4b_1 _2896_ (.A(_0704_),
    .B(_0614_),
    .C(_0705_),
    .D_N(_0440_),
    .X(_0706_));
 sky130_fd_sc_hd__o41a_1 _2897_ (.A1(_1407_),
    .A2(_0429_),
    .A3(_0626_),
    .A4(_0703_),
    .B1(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_4 _2898_ (.A(_0986_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__a21o_1 _2899_ (.A1(gpio[0]),
    .A2(_0708_),
    .B1(_0637_),
    .X(_0091_));
 sky130_fd_sc_hd__a21bo_1 _2900_ (.A1(gpio[1]),
    .A2(_0708_),
    .B1_N(_0279_),
    .X(_0092_));
 sky130_fd_sc_hd__a21o_1 _2901_ (.A1(gpio[2]),
    .A2(_0708_),
    .B1(_0466_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _2902_ (.A(gpio[3]),
    .B(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _2903_ (.A(_0201_),
    .B(_0709_),
    .Y(_0094_));
 sky130_fd_sc_hd__nand2_1 _2904_ (.A(gpio[4]),
    .B(_0708_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _2905_ (.A(_0180_),
    .B(_0710_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_1 _2906_ (.A(gpio[5]),
    .B(_0708_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _2907_ (.A(_0159_),
    .B(_0711_),
    .Y(_0096_));
 sky130_fd_sc_hd__nand2_1 _2908_ (.A(gpio[6]),
    .B(_0708_),
    .Y(_0712_));
 sky130_fd_sc_hd__nand2_1 _2909_ (.A(_0135_),
    .B(_0712_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _2910_ (.A(gpio[7]),
    .B(_0708_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _2911_ (.A(_0320_),
    .B(_0713_),
    .Y(_0098_));
 sky130_fd_sc_hd__nor2_1 _2912_ (.A(_1249_),
    .B(_1251_),
    .Y(_0714_));
 sky130_fd_sc_hd__or4bb_1 _2913_ (.A(_0982_),
    .B(_1286_),
    .C_N(net31),
    .D_N(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__nor3_1 _2914_ (.A(_0353_),
    .B(_0346_),
    .C(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a31o_4 _2915_ (.A1(_0342_),
    .A2(net32),
    .A3(_0716_),
    .B1(_1491_),
    .X(_0717_));
 sky130_fd_sc_hd__or2b_1 _2916_ (.A(_0259_),
    .B_N(_0249_),
    .X(_0718_));
 sky130_fd_sc_hd__xor2_1 _2917_ (.A(_0718_),
    .B(_0258_),
    .X(_0719_));
 sky130_fd_sc_hd__nand2_1 _2918_ (.A(_0351_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__and2_1 _2919_ (.A(_1246_),
    .B(_1376_),
    .X(_0721_));
 sky130_fd_sc_hd__nand2_4 _2920_ (.A(_1209_),
    .B(_0364_),
    .Y(_0722_));
 sky130_fd_sc_hd__nor2_1 _2921_ (.A(_0718_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__a32o_1 _2922_ (.A1(_1247_),
    .A2(_1296_),
    .A3(_0249_),
    .B1(_0272_),
    .B2(_0354_),
    .X(_0724_));
 sky130_fd_sc_hd__a2111o_1 _2923_ (.A1(_0259_),
    .A2(_0721_),
    .B1(_0723_),
    .C1(_0724_),
    .D1(_0351_),
    .X(_0725_));
 sky130_fd_sc_hd__a22o_1 _2924_ (.A1(net74),
    .A2(_0717_),
    .B1(_0720_),
    .B2(_0725_),
    .X(_0099_));
 sky130_fd_sc_hd__a211o_1 _2925_ (.A1(_0204_),
    .A2(_0286_),
    .B1(_0292_),
    .C1(_0287_),
    .X(_0726_));
 sky130_fd_sc_hd__or3_1 _2926_ (.A(_1261_),
    .B(_0290_),
    .C(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__o21ai_1 _2927_ (.A1(_1261_),
    .A2(_0726_),
    .B1(_0290_),
    .Y(_0728_));
 sky130_fd_sc_hd__and2_1 _2928_ (.A(_0282_),
    .B(_0280_),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_2 _2929_ (.A(_1246_),
    .B(_1296_),
    .Y(_0730_));
 sky130_fd_sc_hd__nand2_4 _2930_ (.A(_1246_),
    .B(_1376_),
    .Y(_0731_));
 sky130_fd_sc_hd__o32a_1 _2931_ (.A1(_0283_),
    .A2(_0729_),
    .A3(_0722_),
    .B1(_0216_),
    .B2(_0355_),
    .X(_0732_));
 sky130_fd_sc_hd__o211a_1 _2932_ (.A1(_0729_),
    .A2(_0730_),
    .B1(_0731_),
    .C1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__nor2_1 _2933_ (.A(_0283_),
    .B(_0731_),
    .Y(_0734_));
 sky130_fd_sc_hd__a2bb2o_1 _2934_ (.A1_N(_0733_),
    .A2_N(_0734_),
    .B1(\top8227.internalDataflow.addressLowBusModule.busInputs[25] ),
    .B2(_0717_),
    .X(_0735_));
 sky130_fd_sc_hd__a31o_1 _2935_ (.A1(_0351_),
    .A2(_0727_),
    .A3(_0728_),
    .B1(_0735_),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _2936_ (.A(_0216_),
    .B(_0223_),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_1 _2937_ (.A(_0354_),
    .B(_0194_),
    .Y(_0737_));
 sky130_fd_sc_hd__o221a_1 _2938_ (.A1(_0736_),
    .A2(_0730_),
    .B1(_0722_),
    .B2(_0224_),
    .C1(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__o211a_1 _2939_ (.A1(_0285_),
    .A2(_0731_),
    .B1(_0738_),
    .C1(_0350_),
    .X(_0739_));
 sky130_fd_sc_hd__o21ba_1 _2940_ (.A1(_0350_),
    .A2(_0289_),
    .B1_N(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__nor2_2 _2941_ (.A(_1484_),
    .B(_1259_),
    .Y(_0741_));
 sky130_fd_sc_hd__nor2_1 _2942_ (.A(_0290_),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__and2_1 _2943_ (.A(_0290_),
    .B(_0741_),
    .X(_0743_));
 sky130_fd_sc_hd__or3_1 _2944_ (.A(_0726_),
    .B(_0742_),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__xnor2_1 _2945_ (.A(_0289_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__mux2_1 _2946_ (.A0(_0740_),
    .A1(_0745_),
    .S(_0341_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(_0746_),
    .A1(\top8227.internalDataflow.addressLowBusModule.busInputs[26] ),
    .S(_0717_),
    .X(_0747_));
 sky130_fd_sc_hd__clkbuf_1 _2948_ (.A(_0747_),
    .X(_0101_));
 sky130_fd_sc_hd__and3_1 _2949_ (.A(_0289_),
    .B(_0291_),
    .C(_0741_),
    .X(_0748_));
 sky130_fd_sc_hd__or3_1 _2950_ (.A(_0289_),
    .B(_0291_),
    .C(_0741_),
    .X(_0749_));
 sky130_fd_sc_hd__or4b_1 _2951_ (.A(_1261_),
    .B(_0726_),
    .C(_0748_),
    .D_N(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__a21oi_1 _2952_ (.A1(_0204_),
    .A2(_0286_),
    .B1(_0350_),
    .Y(_0751_));
 sky130_fd_sc_hd__o21a_1 _2953_ (.A1(_0204_),
    .A2(_0286_),
    .B1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__and2_1 _2954_ (.A(_0195_),
    .B(_0202_),
    .X(_0753_));
 sky130_fd_sc_hd__o221a_1 _2955_ (.A1(_0355_),
    .A2(_0175_),
    .B1(_0753_),
    .B2(_0730_),
    .C1(_0731_),
    .X(_0754_));
 sky130_fd_sc_hd__o21ai_1 _2956_ (.A1(_0203_),
    .A2(_0722_),
    .B1(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__o211a_1 _2957_ (.A1(_0287_),
    .A2(_0731_),
    .B1(_0755_),
    .C1(_0350_),
    .X(_0756_));
 sky130_fd_sc_hd__a221o_1 _2958_ (.A1(\top8227.internalDataflow.addressLowBusModule.busInputs[27] ),
    .A2(_0717_),
    .B1(_0750_),
    .B2(_0752_),
    .C1(_0756_),
    .X(_0102_));
 sky130_fd_sc_hd__nand2_1 _2959_ (.A(_0351_),
    .B(_0335_),
    .Y(_0757_));
 sky130_fd_sc_hd__a21o_1 _2960_ (.A1(_0295_),
    .A2(_0288_),
    .B1(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__or2_1 _2961_ (.A(_0295_),
    .B(_0722_),
    .X(_0759_));
 sky130_fd_sc_hd__o221a_1 _2962_ (.A1(_0355_),
    .A2(_0152_),
    .B1(_0293_),
    .B2(_0730_),
    .C1(_0731_),
    .X(_0760_));
 sky130_fd_sc_hd__a22o_1 _2963_ (.A1(_0182_),
    .A2(_0721_),
    .B1(_0759_),
    .B2(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__a21oi_1 _2964_ (.A1(_0758_),
    .A2(_0761_),
    .B1(_0341_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand3_1 _2965_ (.A(_0295_),
    .B(_0288_),
    .C(_0292_),
    .Y(_0763_));
 sky130_fd_sc_hd__a32o_1 _2966_ (.A1(_0341_),
    .A2(_0296_),
    .A3(_0763_),
    .B1(_0717_),
    .B2(\top8227.internalDataflow.addressLowBusModule.busInputs[28] ),
    .X(_0764_));
 sky130_fd_sc_hd__or2_1 _2967_ (.A(_0762_),
    .B(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_0765_),
    .X(_0103_));
 sky130_fd_sc_hd__nand3_1 _2969_ (.A(_0299_),
    .B(_0182_),
    .C(_0335_),
    .Y(_0766_));
 sky130_fd_sc_hd__o221a_1 _2970_ (.A1(_0355_),
    .A2(_1483_),
    .B1(_0298_),
    .B2(_0730_),
    .C1(_0731_),
    .X(_0767_));
 sky130_fd_sc_hd__o21a_1 _2971_ (.A1(_0299_),
    .A2(_0722_),
    .B1(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__a21oi_1 _2972_ (.A1(_0161_),
    .A2(_0721_),
    .B1(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__a311o_1 _2973_ (.A1(_0351_),
    .A2(_0336_),
    .A3(_0766_),
    .B1(_0769_),
    .C1(_0341_),
    .X(_0770_));
 sky130_fd_sc_hd__a21oi_2 _2974_ (.A1(_0332_),
    .A2(_0333_),
    .B1(_0323_),
    .Y(_0771_));
 sky130_fd_sc_hd__a21oi_1 _2975_ (.A1(_0331_),
    .A2(_0771_),
    .B1(_0329_),
    .Y(_0772_));
 sky130_fd_sc_hd__and3_1 _2976_ (.A(_0329_),
    .B(_0331_),
    .C(_0771_),
    .X(_0773_));
 sky130_fd_sc_hd__or3_1 _2977_ (.A(_1261_),
    .B(_0772_),
    .C(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _2978_ (.A1(net69),
    .A2(_0717_),
    .B1(_0770_),
    .B2(_0774_),
    .X(_0104_));
 sky130_fd_sc_hd__or2_1 _2979_ (.A(_0303_),
    .B(_0722_),
    .X(_0775_));
 sky130_fd_sc_hd__o221a_1 _2980_ (.A1(_0355_),
    .A2(_0315_),
    .B1(_0301_),
    .B2(_0730_),
    .C1(_0731_),
    .X(_0776_));
 sky130_fd_sc_hd__a22o_1 _2981_ (.A1(_0141_),
    .A2(_0721_),
    .B1(_0775_),
    .B2(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _2982_ (.A(_0351_),
    .B(_0337_),
    .Y(_0778_));
 sky130_fd_sc_hd__a31o_1 _2983_ (.A1(_0303_),
    .A2(_0161_),
    .A3(_0336_),
    .B1(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__a21oi_1 _2984_ (.A1(_0777_),
    .A2(_0779_),
    .B1(_0341_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand2_1 _2985_ (.A(_0304_),
    .B(_0327_),
    .Y(_0781_));
 sky130_fd_sc_hd__xnor2_1 _2986_ (.A(_0781_),
    .B(_0329_),
    .Y(_0782_));
 sky130_fd_sc_hd__xnor2_1 _2987_ (.A(_0741_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__nor2_1 _2988_ (.A(_0325_),
    .B(_0326_),
    .Y(_0784_));
 sky130_fd_sc_hd__o31a_1 _2989_ (.A1(_0329_),
    .A2(_0784_),
    .A3(_0334_),
    .B1(_0781_),
    .X(_0785_));
 sky130_fd_sc_hd__a311oi_1 _2990_ (.A1(_0331_),
    .A2(_0771_),
    .A3(_0783_),
    .B1(_0785_),
    .C1(_1261_),
    .Y(_0786_));
 sky130_fd_sc_hd__a211o_1 _2991_ (.A1(net63),
    .A2(_0717_),
    .B1(_0780_),
    .C1(_0786_),
    .X(_0105_));
 sky130_fd_sc_hd__or3b_1 _2992_ (.A(_0781_),
    .B(_0329_),
    .C_N(_0741_),
    .X(_0787_));
 sky130_fd_sc_hd__a31o_1 _2993_ (.A1(_0330_),
    .A2(_0771_),
    .A3(_0787_),
    .B1(_0784_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _2994_ (.A(_0341_),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _2995_ (.A(_0324_),
    .Y(_0790_));
 sky130_fd_sc_hd__a21oi_1 _2996_ (.A1(_0338_),
    .A2(_0790_),
    .B1(_0350_),
    .Y(_0791_));
 sky130_fd_sc_hd__o21a_1 _2997_ (.A1(_0338_),
    .A2(_0790_),
    .B1(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__a2bb2o_1 _2998_ (.A1_N(_0322_),
    .A2_N(_0730_),
    .B1(_0258_),
    .B2(_0354_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(_0324_),
    .A1(_0793_),
    .S(_0722_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _3000_ (.A0(_0323_),
    .A1(_0794_),
    .S(_0731_),
    .X(_0795_));
 sky130_fd_sc_hd__or3_1 _3001_ (.A(_0341_),
    .B(_0792_),
    .C(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__a22o_1 _3002_ (.A1(net78),
    .A2(_0717_),
    .B1(_0789_),
    .B2(_0796_),
    .X(_0106_));
 sky130_fd_sc_hd__o21a_1 _3003_ (.A1(_0943_),
    .A2(_1121_),
    .B1(_1006_),
    .X(_0797_));
 sky130_fd_sc_hd__o21a_1 _3004_ (.A1(_0902_),
    .A2(_0949_),
    .B1(_1015_),
    .X(_0798_));
 sky130_fd_sc_hd__o21a_4 _3005_ (.A1(_0797_),
    .A2(_0798_),
    .B1(_1247_),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _3006_ (.A0(net80),
    .A1(_0238_),
    .S(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_1 _3007_ (.A(_0800_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _3008_ (.A0(\top8227.internalDataflow.stackBusModule.busInputs[33] ),
    .A1(_0271_),
    .S(_0799_),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_1 _3009_ (.A(_0801_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(net83),
    .A1(_0215_),
    .S(_0799_),
    .X(_0802_));
 sky130_fd_sc_hd__clkbuf_1 _3011_ (.A(_0802_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _3012_ (.A0(net70),
    .A1(_0193_),
    .S(_0799_),
    .X(_0803_));
 sky130_fd_sc_hd__clkbuf_1 _3013_ (.A(_0803_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _3014_ (.A0(net87),
    .A1(_0174_),
    .S(_0799_),
    .X(_0804_));
 sky130_fd_sc_hd__clkbuf_1 _3015_ (.A(_0804_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(net92),
    .A1(_0151_),
    .S(_0799_),
    .X(_0805_));
 sky130_fd_sc_hd__clkbuf_1 _3017_ (.A(_0805_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(\top8227.internalDataflow.stackBusModule.busInputs[38] ),
    .A1(_1482_),
    .S(_0799_),
    .X(_0806_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_0806_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(net89),
    .A1(_0314_),
    .S(_0799_),
    .X(_0807_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_0807_),
    .X(_0114_));
 sky130_fd_sc_hd__or3b_1 _3022_ (.A(_0396_),
    .B(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ),
    .C_N(_1021_),
    .X(_0808_));
 sky130_fd_sc_hd__a2bb2o_1 _3023_ (.A1_N(_0357_),
    .A2_N(_0808_),
    .B1(_0396_),
    .B2(net57),
    .X(_0115_));
 sky130_fd_sc_hd__or4_1 _3024_ (.A(\top8227.demux.state_machine.currentAddress[8] ),
    .B(\top8227.demux.state_machine.currentAddress[0] ),
    .C(\top8227.demux.state_machine.currentAddress[2] ),
    .D(\top8227.demux.state_machine.currentAddress[9] ),
    .X(_0809_));
 sky130_fd_sc_hd__o21ai_1 _3025_ (.A1(_0809_),
    .A2(_0999_),
    .B1(\top8227.demux.isAddressing ),
    .Y(_0810_));
 sky130_fd_sc_hd__o22a_1 _3026_ (.A1(\top8227.demux.isAddressing ),
    .A2(_0979_),
    .B1(_0810_),
    .B2(_1010_),
    .X(_0116_));
 sky130_fd_sc_hd__a21bo_1 _3027_ (.A1(_1015_),
    .A2(_0923_),
    .B1_N(_0387_),
    .X(_0811_));
 sky130_fd_sc_hd__o31a_1 _3028_ (.A1(_1344_),
    .A2(_0373_),
    .A3(_0811_),
    .B1(_1247_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _3029_ (.A0(\top8227.PSRCurrentValue[7] ),
    .A1(_0316_),
    .S(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_1 _3030_ (.A(_0813_),
    .X(_0117_));
 sky130_fd_sc_hd__dfstp_1 _3031_ (.CLK(clknet_4_10_0_clk),
    .D(_0000_),
    .SET_B(net47),
    .Q(\top8227.demux.state_machine.currentAddress[0] ));
 sky130_fd_sc_hd__dfrtp_2 _3032_ (.CLK(clknet_4_12_0_clk),
    .D(_0004_),
    .RESET_B(net45),
    .Q(\top8227.demux.state_machine.currentAddress[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3033_ (.CLK(clknet_4_10_0_clk),
    .D(_0005_),
    .RESET_B(net47),
    .Q(\top8227.demux.state_machine.currentAddress[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3034_ (.CLK(clknet_4_11_0_clk),
    .D(_0006_),
    .RESET_B(net45),
    .Q(\top8227.demux.state_machine.currentAddress[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3035_ (.CLK(clknet_4_10_0_clk),
    .D(_0007_),
    .RESET_B(net45),
    .Q(\top8227.demux.state_machine.currentAddress[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3036_ (.CLK(clknet_4_10_0_clk),
    .D(_0008_),
    .RESET_B(net46),
    .Q(\top8227.demux.state_machine.currentAddress[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3037_ (.CLK(clknet_4_14_0_clk),
    .D(_0009_),
    .RESET_B(net46),
    .Q(\top8227.demux.state_machine.currentAddress[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3038_ (.CLK(clknet_4_11_0_clk),
    .D(_0010_),
    .RESET_B(net45),
    .Q(\top8227.demux.state_machine.currentAddress[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3039_ (.CLK(clknet_4_10_0_clk),
    .D(_0011_),
    .RESET_B(net47),
    .Q(\top8227.demux.state_machine.currentAddress[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3040_ (.CLK(clknet_4_10_0_clk),
    .D(_0012_),
    .RESET_B(net47),
    .Q(\top8227.demux.state_machine.currentAddress[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3041_ (.CLK(clknet_4_10_0_clk),
    .D(_0001_),
    .RESET_B(net46),
    .Q(\top8227.demux.state_machine.currentAddress[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3042_ (.CLK(clknet_4_12_0_clk),
    .D(_0002_),
    .RESET_B(net46),
    .Q(\top8227.demux.state_machine.currentAddress[11] ));
 sky130_fd_sc_hd__dfrtp_4 _3043_ (.CLK(clknet_4_11_0_clk),
    .D(_0003_),
    .RESET_B(net45),
    .Q(\top8227.demux.state_machine.currentAddress[12] ));
 sky130_fd_sc_hd__dfstp_1 _3044_ (.CLK(clknet_4_15_0_clk),
    .D(_0013_),
    .SET_B(net48),
    .Q(\top8227.demux.state_machine.timeState[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3045_ (.CLK(clknet_4_13_0_clk),
    .D(_0014_),
    .RESET_B(net48),
    .Q(\top8227.demux.state_machine.timeState[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3046_ (.CLK(clknet_4_13_0_clk),
    .D(_0015_),
    .RESET_B(net48),
    .Q(\top8227.demux.state_machine.timeState[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3047_ (.CLK(clknet_4_13_0_clk),
    .D(_0016_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.timeState[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3048_ (.CLK(clknet_4_13_0_clk),
    .D(_0017_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.timeState[4] ));
 sky130_fd_sc_hd__dfrtp_2 _3049_ (.CLK(clknet_4_13_0_clk),
    .D(_0018_),
    .RESET_B(net48),
    .Q(\top8227.demux.state_machine.timeState[5] ));
 sky130_fd_sc_hd__dfrtp_2 _3050_ (.CLK(clknet_4_13_0_clk),
    .D(_0019_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.timeState[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3051_ (.CLK(clknet_4_6_0_clk),
    .D(_0026_),
    .RESET_B(net43),
    .Q(\top8227.branchForward ));
 sky130_fd_sc_hd__dfrtp_4 _3052_ (.CLK(clknet_4_15_0_clk),
    .D(_0020_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.currentInstruction[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3053_ (.CLK(clknet_4_15_0_clk),
    .D(_0021_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.currentInstruction[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3054_ (.CLK(clknet_4_14_0_clk),
    .D(_0022_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.currentInstruction[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3055_ (.CLK(clknet_4_15_0_clk),
    .D(_0023_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.currentInstruction[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3056_ (.CLK(clknet_4_14_0_clk),
    .D(_0024_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.currentInstruction[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3057_ (.CLK(clknet_4_14_0_clk),
    .D(_0025_),
    .RESET_B(net49),
    .Q(\top8227.demux.state_machine.currentInstruction[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3058_ (.CLK(clknet_4_12_0_clk),
    .D(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[0] ),
    .RESET_B(net39),
    .Q(\top8227.PSRCurrentValue[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3059_ (.CLK(clknet_4_12_0_clk),
    .D(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[1] ),
    .RESET_B(net39),
    .Q(\top8227.PSRCurrentValue[1] ));
 sky130_fd_sc_hd__dfrtp_2 _3060_ (.CLK(clknet_4_9_0_clk),
    .D(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[2] ),
    .RESET_B(net38),
    .Q(\top8227.PSRCurrentValue[2] ));
 sky130_fd_sc_hd__dfrtp_2 _3061_ (.CLK(clknet_4_9_0_clk),
    .D(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[3] ),
    .RESET_B(net39),
    .Q(\top8227.PSRCurrentValue[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3062_ (.CLK(clknet_4_9_0_clk),
    .D(\top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt[6] ),
    .RESET_B(net38),
    .Q(\top8227.PSRCurrentValue[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3063_ (.CLK(clknet_4_9_0_clk),
    .D(_0027_),
    .RESET_B(net45),
    .Q(\top8227.freeCarry ));
 sky130_fd_sc_hd__dfstp_1 _3064_ (.CLK(clknet_4_8_0_clk),
    .D(_0028_),
    .SET_B(net45),
    .Q(\top8227.instructionLoader.interruptInjector.resetDetected ));
 sky130_fd_sc_hd__dfrtp_1 _3065_ (.CLK(clknet_4_8_0_clk),
    .D(_0029_),
    .RESET_B(net38),
    .Q(\top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ));
 sky130_fd_sc_hd__dfrtp_1 _3066_ (.CLK(clknet_4_6_0_clk),
    .D(_0030_),
    .RESET_B(net48),
    .Q(\top8227.negEdgeDetector.q1 ));
 sky130_fd_sc_hd__dfrtp_2 _3067_ (.CLK(clknet_4_11_0_clk),
    .D(_0031_),
    .RESET_B(net38),
    .Q(\top8227.demux.setInterruptFlag ));
 sky130_fd_sc_hd__dfrtp_4 _3068_ (.CLK(clknet_4_8_0_clk),
    .D(_0032_),
    .RESET_B(net38),
    .Q(\top8227.demux.nmi ));
 sky130_fd_sc_hd__dfrtp_4 _3069_ (.CLK(clknet_4_8_0_clk),
    .D(_0033_),
    .RESET_B(net39),
    .Q(\top8227.instructionLoader.interruptInjector.irqGenerated ));
 sky130_fd_sc_hd__dfrtp_1 _3070_ (.CLK(clknet_4_15_0_clk),
    .D(\top8227.instructionLoader.interruptInjector.interruptRequest ),
    .RESET_B(net50),
    .Q(\top8227.instructionLoader.interruptInjector.irqSync.nextQ2 ));
 sky130_fd_sc_hd__dfrtp_2 _3071_ (.CLK(clknet_4_15_0_clk),
    .D(net51),
    .RESET_B(net50),
    .Q(\top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ ));
 sky130_fd_sc_hd__dfrtp_1 _3072_ (.CLK(clknet_4_2_0_clk),
    .D(\top8227.instructionLoader.interruptInjector.nmiSync.in ),
    .RESET_B(net37),
    .Q(\top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 ));
 sky130_fd_sc_hd__dfrtp_1 _3073_ (.CLK(clknet_4_8_0_clk),
    .D(net52),
    .RESET_B(net38),
    .Q(\top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI ));
 sky130_fd_sc_hd__dfrtp_1 _3074_ (.CLK(clknet_4_7_0_clk),
    .D(_0034_),
    .RESET_B(net48),
    .Q(net10));
 sky130_fd_sc_hd__dfrtp_1 _3075_ (.CLK(clknet_4_8_0_clk),
    .D(_0035_),
    .RESET_B(net38),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_1 _3076_ (.CLK(clknet_4_2_0_clk),
    .D(_0036_),
    .RESET_B(net34),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _3077_ (.CLK(clknet_4_6_0_clk),
    .D(_0037_),
    .RESET_B(net42),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _3078_ (.CLK(clknet_4_8_0_clk),
    .D(_0038_),
    .RESET_B(net38),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _3079_ (.CLK(clknet_4_2_0_clk),
    .D(_0039_),
    .RESET_B(net37),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _3080_ (.CLK(clknet_4_7_0_clk),
    .D(_0040_),
    .RESET_B(net48),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_1 _3081_ (.CLK(clknet_4_5_0_clk),
    .D(_0041_),
    .RESET_B(net41),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_2 _3082_ (.CLK(clknet_4_5_0_clk),
    .D(_0042_),
    .RESET_B(net41),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[16] ));
 sky130_fd_sc_hd__dfrtp_4 _3083_ (.CLK(clknet_4_5_0_clk),
    .D(_0043_),
    .RESET_B(net42),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[17] ));
 sky130_fd_sc_hd__dfrtp_4 _3084_ (.CLK(clknet_4_5_0_clk),
    .D(_0044_),
    .RESET_B(net41),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[18] ));
 sky130_fd_sc_hd__dfrtp_4 _3085_ (.CLK(clknet_4_5_0_clk),
    .D(_0045_),
    .RESET_B(net41),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[19] ));
 sky130_fd_sc_hd__dfrtp_2 _3086_ (.CLK(clknet_4_4_0_clk),
    .D(_0046_),
    .RESET_B(net41),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[20] ));
 sky130_fd_sc_hd__dfrtp_2 _3087_ (.CLK(clknet_4_4_0_clk),
    .D(_0047_),
    .RESET_B(net41),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[21] ));
 sky130_fd_sc_hd__dfrtp_2 _3088_ (.CLK(clknet_4_4_0_clk),
    .D(_0048_),
    .RESET_B(net41),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[22] ));
 sky130_fd_sc_hd__dfrtp_2 _3089_ (.CLK(clknet_4_4_0_clk),
    .D(_0049_),
    .RESET_B(net41),
    .Q(\top8227.internalDataflow.addressHighBusModule.busInputs[23] ));
 sky130_fd_sc_hd__dfrtp_1 _3090_ (.CLK(clknet_4_1_0_clk),
    .D(_0050_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[32] ));
 sky130_fd_sc_hd__dfrtp_1 _3091_ (.CLK(clknet_4_6_0_clk),
    .D(_0051_),
    .RESET_B(net43),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[33] ));
 sky130_fd_sc_hd__dfrtp_1 _3092_ (.CLK(clknet_4_0_0_clk),
    .D(_0052_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[34] ));
 sky130_fd_sc_hd__dfrtp_1 _3093_ (.CLK(clknet_4_3_0_clk),
    .D(_0053_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[35] ));
 sky130_fd_sc_hd__dfrtp_1 _3094_ (.CLK(clknet_4_0_0_clk),
    .D(_0054_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[36] ));
 sky130_fd_sc_hd__dfrtp_1 _3095_ (.CLK(clknet_4_0_0_clk),
    .D(_0055_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[37] ));
 sky130_fd_sc_hd__dfrtp_1 _3096_ (.CLK(clknet_4_1_0_clk),
    .D(_0056_),
    .RESET_B(net40),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[38] ));
 sky130_fd_sc_hd__dfrtp_1 _3097_ (.CLK(clknet_4_0_0_clk),
    .D(_0057_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[39] ));
 sky130_fd_sc_hd__dfrtp_1 _3098_ (.CLK(clknet_4_3_0_clk),
    .D(_0058_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[40] ));
 sky130_fd_sc_hd__dfrtp_1 _3099_ (.CLK(clknet_4_9_0_clk),
    .D(_0059_),
    .RESET_B(net39),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[41] ));
 sky130_fd_sc_hd__dfrtp_1 _3100_ (.CLK(clknet_4_3_0_clk),
    .D(_0060_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[42] ));
 sky130_fd_sc_hd__dfrtp_1 _3101_ (.CLK(clknet_4_3_0_clk),
    .D(_0061_),
    .RESET_B(net36),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[43] ));
 sky130_fd_sc_hd__dfrtp_1 _3102_ (.CLK(clknet_4_0_0_clk),
    .D(_0062_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[44] ));
 sky130_fd_sc_hd__dfrtp_1 _3103_ (.CLK(clknet_4_0_0_clk),
    .D(_0063_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[45] ));
 sky130_fd_sc_hd__dfrtp_1 _3104_ (.CLK(clknet_4_0_0_clk),
    .D(_0064_),
    .RESET_B(net35),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[46] ));
 sky130_fd_sc_hd__dfrtp_1 _3105_ (.CLK(clknet_4_3_0_clk),
    .D(_0065_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[47] ));
 sky130_fd_sc_hd__dfrtp_4 _3106_ (.CLK(clknet_4_8_0_clk),
    .D(_0066_),
    .RESET_B(net45),
    .Q(\top8227.demux.reset ));
 sky130_fd_sc_hd__dfrtp_4 _3107_ (.CLK(clknet_4_1_0_clk),
    .D(_0067_),
    .RESET_B(net40),
    .Q(gpio[8]));
 sky130_fd_sc_hd__dfrtp_4 _3108_ (.CLK(clknet_4_5_0_clk),
    .D(_0068_),
    .RESET_B(net41),
    .Q(gpio[9]));
 sky130_fd_sc_hd__dfrtp_4 _3109_ (.CLK(clknet_4_1_0_clk),
    .D(_0069_),
    .RESET_B(net40),
    .Q(gpio[10]));
 sky130_fd_sc_hd__dfrtp_4 _3110_ (.CLK(clknet_4_7_0_clk),
    .D(_0070_),
    .RESET_B(net42),
    .Q(gpio[11]));
 sky130_fd_sc_hd__dfrtp_4 _3111_ (.CLK(clknet_4_5_0_clk),
    .D(_0071_),
    .RESET_B(net44),
    .Q(gpio[12]));
 sky130_fd_sc_hd__dfrtp_4 _3112_ (.CLK(clknet_4_1_0_clk),
    .D(_0072_),
    .RESET_B(net40),
    .Q(gpio[13]));
 sky130_fd_sc_hd__dfrtp_4 _3113_ (.CLK(clknet_4_5_0_clk),
    .D(_0073_),
    .RESET_B(net44),
    .Q(gpio[14]));
 sky130_fd_sc_hd__dfrtp_4 _3114_ (.CLK(clknet_4_4_0_clk),
    .D(_0074_),
    .RESET_B(net40),
    .Q(gpio[15]));
 sky130_fd_sc_hd__dfrtp_4 _3115_ (.CLK(clknet_4_7_0_clk),
    .D(_0075_),
    .RESET_B(net42),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[16] ));
 sky130_fd_sc_hd__dfrtp_4 _3116_ (.CLK(clknet_4_6_0_clk),
    .D(_0076_),
    .RESET_B(net42),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[17] ));
 sky130_fd_sc_hd__dfrtp_4 _3117_ (.CLK(clknet_4_7_0_clk),
    .D(_0077_),
    .RESET_B(net43),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[18] ));
 sky130_fd_sc_hd__dfrtp_4 _3118_ (.CLK(clknet_4_7_0_clk),
    .D(_0078_),
    .RESET_B(net43),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[19] ));
 sky130_fd_sc_hd__dfrtp_2 _3119_ (.CLK(clknet_4_6_0_clk),
    .D(_0079_),
    .RESET_B(net42),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[20] ));
 sky130_fd_sc_hd__dfrtp_4 _3120_ (.CLK(clknet_4_4_0_clk),
    .D(_0080_),
    .RESET_B(net42),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[21] ));
 sky130_fd_sc_hd__dfrtp_4 _3121_ (.CLK(clknet_4_5_0_clk),
    .D(_0081_),
    .RESET_B(net42),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[22] ));
 sky130_fd_sc_hd__dfrtp_4 _3122_ (.CLK(clknet_4_7_0_clk),
    .D(_0082_),
    .RESET_B(net43),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[23] ));
 sky130_fd_sc_hd__dfrtp_2 _3123_ (.CLK(clknet_4_3_0_clk),
    .D(_0083_),
    .RESET_B(net36),
    .Q(\top8227.internalDataflow.accRegToDB[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3124_ (.CLK(clknet_4_3_0_clk),
    .D(_0084_),
    .RESET_B(net39),
    .Q(\top8227.internalDataflow.accRegToDB[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3125_ (.CLK(clknet_4_1_0_clk),
    .D(_0085_),
    .RESET_B(net40),
    .Q(\top8227.internalDataflow.accRegToDB[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3126_ (.CLK(clknet_4_3_0_clk),
    .D(_0086_),
    .RESET_B(net39),
    .Q(\top8227.internalDataflow.accRegToDB[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3127_ (.CLK(clknet_4_1_0_clk),
    .D(_0087_),
    .RESET_B(net40),
    .Q(\top8227.internalDataflow.accRegToDB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3128_ (.CLK(clknet_4_1_0_clk),
    .D(_0088_),
    .RESET_B(net40),
    .Q(\top8227.internalDataflow.accRegToDB[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3129_ (.CLK(clknet_4_1_0_clk),
    .D(_0089_),
    .RESET_B(net40),
    .Q(\top8227.internalDataflow.accRegToDB[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3130_ (.CLK(clknet_4_1_0_clk),
    .D(_0090_),
    .RESET_B(net40),
    .Q(\top8227.internalDataflow.accRegToDB[7] ));
 sky130_fd_sc_hd__dfrtp_4 _3131_ (.CLK(clknet_4_7_0_clk),
    .D(_0091_),
    .RESET_B(net48),
    .Q(gpio[0]));
 sky130_fd_sc_hd__dfrtp_4 _3132_ (.CLK(clknet_4_11_0_clk),
    .D(_0092_),
    .RESET_B(net45),
    .Q(gpio[1]));
 sky130_fd_sc_hd__dfrtp_4 _3133_ (.CLK(clknet_4_8_0_clk),
    .D(_0093_),
    .RESET_B(net38),
    .Q(gpio[2]));
 sky130_fd_sc_hd__dfrtp_4 _3134_ (.CLK(clknet_4_4_0_clk),
    .D(_0094_),
    .RESET_B(net43),
    .Q(gpio[3]));
 sky130_fd_sc_hd__dfrtp_4 _3135_ (.CLK(clknet_4_7_0_clk),
    .D(_0095_),
    .RESET_B(net48),
    .Q(gpio[4]));
 sky130_fd_sc_hd__dfrtp_4 _3136_ (.CLK(clknet_4_5_0_clk),
    .D(_0096_),
    .RESET_B(net42),
    .Q(gpio[5]));
 sky130_fd_sc_hd__dfrtp_4 _3137_ (.CLK(clknet_4_7_0_clk),
    .D(_0097_),
    .RESET_B(net42),
    .Q(gpio[6]));
 sky130_fd_sc_hd__dfrtp_4 _3138_ (.CLK(clknet_4_11_0_clk),
    .D(_0098_),
    .RESET_B(net45),
    .Q(gpio[7]));
 sky130_fd_sc_hd__dfrtp_1 _3139_ (.CLK(clknet_4_9_0_clk),
    .D(_0099_),
    .RESET_B(net39),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[24] ));
 sky130_fd_sc_hd__dfrtp_2 _3140_ (.CLK(clknet_4_8_0_clk),
    .D(_0100_),
    .RESET_B(net38),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[25] ));
 sky130_fd_sc_hd__dfrtp_1 _3141_ (.CLK(clknet_4_2_0_clk),
    .D(_0101_),
    .RESET_B(net37),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[26] ));
 sky130_fd_sc_hd__dfrtp_1 _3142_ (.CLK(clknet_4_2_0_clk),
    .D(_0102_),
    .RESET_B(net39),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[27] ));
 sky130_fd_sc_hd__dfrtp_4 _3143_ (.CLK(clknet_4_2_0_clk),
    .D(_0103_),
    .RESET_B(net37),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[28] ));
 sky130_fd_sc_hd__dfrtp_2 _3144_ (.CLK(clknet_4_2_0_clk),
    .D(_0104_),
    .RESET_B(net37),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[29] ));
 sky130_fd_sc_hd__dfrtp_2 _3145_ (.CLK(clknet_4_2_0_clk),
    .D(_0105_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[30] ));
 sky130_fd_sc_hd__dfrtp_1 _3146_ (.CLK(clknet_4_2_0_clk),
    .D(_0106_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.addressLowBusModule.busInputs[31] ));
 sky130_fd_sc_hd__dfrtp_1 _3147_ (.CLK(clknet_4_7_0_clk),
    .D(\top8227.pulse_slower.nextEnableState[0] ),
    .RESET_B(net43),
    .Q(\top8227.pulse_slower.currentEnableState[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3148_ (.CLK(clknet_4_7_0_clk),
    .D(\top8227.pulse_slower.nextEnableState[1] ),
    .RESET_B(net48),
    .Q(\top8227.pulse_slower.currentEnableState[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3149_ (.CLK(clknet_4_3_0_clk),
    .D(_0107_),
    .RESET_B(net36),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[32] ));
 sky130_fd_sc_hd__dfrtp_1 _3150_ (.CLK(clknet_4_9_0_clk),
    .D(_0108_),
    .RESET_B(net44),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[33] ));
 sky130_fd_sc_hd__dfrtp_1 _3151_ (.CLK(clknet_4_2_0_clk),
    .D(_0109_),
    .RESET_B(net36),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[34] ));
 sky130_fd_sc_hd__dfrtp_1 _3152_ (.CLK(clknet_4_3_0_clk),
    .D(_0110_),
    .RESET_B(net36),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[35] ));
 sky130_fd_sc_hd__dfrtp_1 _3153_ (.CLK(clknet_4_2_0_clk),
    .D(_0111_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[36] ));
 sky130_fd_sc_hd__dfrtp_1 _3154_ (.CLK(clknet_4_2_0_clk),
    .D(_0112_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[37] ));
 sky130_fd_sc_hd__dfrtp_1 _3155_ (.CLK(clknet_4_2_0_clk),
    .D(_0113_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[38] ));
 sky130_fd_sc_hd__dfrtp_1 _3156_ (.CLK(clknet_4_2_0_clk),
    .D(_0114_),
    .RESET_B(net34),
    .Q(\top8227.internalDataflow.stackBusModule.busInputs[39] ));
 sky130_fd_sc_hd__dfrtp_1 _3157_ (.CLK(clknet_4_6_0_clk),
    .D(_0115_),
    .RESET_B(net43),
    .Q(\top8227.branchBackward ));
 sky130_fd_sc_hd__dfstp_1 _3158_ (.CLK(clknet_4_10_0_clk),
    .D(_0116_),
    .SET_B(net46),
    .Q(\top8227.demux.isAddressing ));
 sky130_fd_sc_hd__dfrtp_4 _3159_ (.CLK(clknet_4_12_0_clk),
    .D(_0117_),
    .RESET_B(net44),
    .Q(\top8227.PSRCurrentValue[7] ));
 sky130_fd_sc_hd__buf_2 _3160_ (.A(clknet_4_2_0_clk),
    .X(gpio[23]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net37),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net44),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net44),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_4 fanout41 (.A(net44),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net50),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net47),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net50),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net9),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\top8227.instructionLoader.interruptInjector.irqSync.nextQ2 ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\top8227.demux.state_machine.currentAddress[4] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\top8227.demux.state_machine.currentAddress[11] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\top8227.instructionLoader.interruptInjector.irqGenerated ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[30] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\top8227.pulse_slower.currentEnableState[0] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\top8227.internalDataflow.stackBusModule.busInputs[44] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\top8227.internalDataflow.stackBusModule.busInputs[46] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\top8227.demux.setInterruptFlag ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\top8227.internalDataflow.stackBusModule.busInputs[42] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[29] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\top8227.internalDataflow.stackBusModule.busInputs[35] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\top8227.internalDataflow.stackBusModule.busInputs[45] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\top8227.internalDataflow.stackBusModule.busInputs[43] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\top8227.demux.state_machine.timeState[3] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[24] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[16] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[22] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\top8227.demux.state_machine.currentAddress[10] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[31] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net12),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\top8227.internalDataflow.stackBusModule.busInputs[32] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\top8227.internalDataflow.stackBusModule.busInputs[47] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\top8227.negEdgeDetector.q1 ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\top8227.internalDataflow.stackBusModule.busInputs[34] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net17),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net11),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net15),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\top8227.internalDataflow.stackBusModule.busInputs[36] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\top8227.internalDataflow.addressLowBusModule.busInputs[20] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\top8227.internalDataflow.stackBusModule.busInputs[39] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\top8227.demux.state_machine.currentAddress[8] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\top8227.internalDataflow.addressHighBusModule.busInputs[17] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\top8227.demux.state_machine.currentAddress[2] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\top8227.internalDataflow.stackBusModule.busInputs[37] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\top8227.instructionLoader.interruptInjector.resetDetected ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\top8227.branchForward ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\top8227.branchBackward ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\top8227.demux.state_machine.currentAddress[3] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\top8227.demux.state_machine.currentAddress[0] ),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(dataBusIn[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(dataBusIn[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(dataBusIn[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(dataBusIn[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(dataBusIn[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(dataBusIn[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(dataBusIn[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(dataBusIn[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(nrst),
    .X(net9));
 sky130_fd_sc_hd__buf_1 max_cap1 (.A(_1395_),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 max_cap19 (.A(_1440_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(_1477_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 max_cap20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 max_cap21 (.A(_1395_),
    .X(net21));
 sky130_fd_sc_hd__buf_2 max_cap22 (.A(_0691_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 max_cap24 (.A(_0119_),
    .X(net24));
 sky130_fd_sc_hd__buf_1 max_cap26 (.A(_1102_),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 max_cap27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 max_cap30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 max_cap32 (.A(_1485_),
    .X(net32));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dataBusOut[0]));
 sky130_fd_sc_hd__clkbuf_4 output11 (.A(net11),
    .X(dataBusOut[1]));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(dataBusOut[2]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dataBusOut[3]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(dataBusOut[4]));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(dataBusOut[5]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(dataBusOut[6]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(dataBusOut[7]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(dataBusSelect));
 sky130_fd_sc_hd__clkbuf_1 wire23 (.A(_0349_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 wire25 (.A(net94),
    .X(net25));
 sky130_fd_sc_hd__buf_1 wire28 (.A(_1418_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 wire29 (.A(_0973_),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 wire31 (.A(_0343_),
    .X(net31));
 sky130_fd_sc_hd__buf_1 wire33 (.A(_0970_),
    .X(net33));
endmodule

